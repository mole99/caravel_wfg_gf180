magic
tech gf180mcuC
magscale 1 10
timestamp 1670096818
<< metal1 >>
rect 1344 76858 78624 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 78624 76858
rect 1344 76772 78624 76806
rect 1344 76074 78624 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 78624 76074
rect 1344 75988 78624 76022
rect 2034 75742 2046 75794
rect 2098 75742 2110 75794
rect 75618 75742 75630 75794
rect 75682 75742 75694 75794
rect 3502 75682 3554 75694
rect 3042 75630 3054 75682
rect 3106 75630 3118 75682
rect 74946 75630 74958 75682
rect 75010 75630 75022 75682
rect 3502 75618 3554 75630
rect 1344 75290 78624 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 78624 75290
rect 1344 75204 78624 75238
rect 3042 74846 3054 74898
rect 3106 74846 3118 74898
rect 74946 74846 74958 74898
rect 75010 74846 75022 74898
rect 3614 74786 3666 74798
rect 1922 74734 1934 74786
rect 1986 74734 1998 74786
rect 75618 74734 75630 74786
rect 75682 74734 75694 74786
rect 3614 74722 3666 74734
rect 1344 74506 78624 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 78624 74506
rect 1344 74420 78624 74454
rect 3266 74174 3278 74226
rect 3330 74174 3342 74226
rect 74946 74174 74958 74226
rect 75010 74174 75022 74226
rect 3838 74002 3890 74014
rect 2258 73950 2270 74002
rect 2322 73950 2334 74002
rect 3838 73938 3890 73950
rect 4174 74002 4226 74014
rect 77310 74002 77362 74014
rect 76290 73950 76302 74002
rect 76354 73950 76366 74002
rect 4174 73938 4226 73950
rect 77310 73938 77362 73950
rect 73614 73890 73666 73902
rect 73614 73826 73666 73838
rect 74062 73890 74114 73902
rect 74062 73826 74114 73838
rect 1344 73722 78624 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 78624 73722
rect 1344 73636 78624 73670
rect 68910 73554 68962 73566
rect 68910 73490 68962 73502
rect 73726 73554 73778 73566
rect 73726 73490 73778 73502
rect 69022 73442 69074 73454
rect 69022 73378 69074 73390
rect 73838 73442 73890 73454
rect 73838 73378 73890 73390
rect 3042 73278 3054 73330
rect 3106 73278 3118 73330
rect 4834 73278 4846 73330
rect 4898 73278 4910 73330
rect 74946 73278 74958 73330
rect 75010 73278 75022 73330
rect 76738 73278 76750 73330
rect 76802 73278 76814 73330
rect 5406 73218 5458 73230
rect 2034 73166 2046 73218
rect 2098 73166 2110 73218
rect 3714 73166 3726 73218
rect 3778 73166 3790 73218
rect 5406 73154 5458 73166
rect 69694 73218 69746 73230
rect 69694 73154 69746 73166
rect 72382 73218 72434 73230
rect 72382 73154 72434 73166
rect 74398 73218 74450 73230
rect 75954 73166 75966 73218
rect 76018 73166 76030 73218
rect 77858 73166 77870 73218
rect 77922 73166 77934 73218
rect 74398 73154 74450 73166
rect 68798 73106 68850 73118
rect 68798 73042 68850 73054
rect 73614 73106 73666 73118
rect 74162 73054 74174 73106
rect 74226 73103 74238 73106
rect 74722 73103 74734 73106
rect 74226 73057 74734 73103
rect 74226 73054 74238 73057
rect 74722 73054 74734 73057
rect 74786 73054 74798 73106
rect 73614 73042 73666 73054
rect 1344 72938 78624 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 78624 72938
rect 1344 72852 78624 72886
rect 74062 72658 74114 72670
rect 74062 72594 74114 72606
rect 74174 72658 74226 72670
rect 74174 72594 74226 72606
rect 72158 72546 72210 72558
rect 3042 72494 3054 72546
rect 3106 72494 3118 72546
rect 73042 72494 73054 72546
rect 73106 72494 73118 72546
rect 75058 72494 75070 72546
rect 75122 72494 75134 72546
rect 72158 72482 72210 72494
rect 69358 72434 69410 72446
rect 1922 72382 1934 72434
rect 1986 72382 1998 72434
rect 69358 72370 69410 72382
rect 70142 72434 70194 72446
rect 70142 72370 70194 72382
rect 71822 72434 71874 72446
rect 71822 72370 71874 72382
rect 73278 72434 73330 72446
rect 76066 72382 76078 72434
rect 76130 72382 76142 72434
rect 73278 72370 73330 72382
rect 3614 72322 3666 72334
rect 3614 72258 3666 72270
rect 3950 72322 4002 72334
rect 3950 72258 4002 72270
rect 69470 72322 69522 72334
rect 69470 72258 69522 72270
rect 69582 72322 69634 72334
rect 69582 72258 69634 72270
rect 73950 72322 74002 72334
rect 73950 72258 74002 72270
rect 1344 72154 78624 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 78624 72154
rect 1344 72068 78624 72102
rect 72494 71986 72546 71998
rect 72494 71922 72546 71934
rect 73390 71986 73442 71998
rect 73390 71922 73442 71934
rect 74062 71986 74114 71998
rect 74062 71922 74114 71934
rect 71262 71874 71314 71886
rect 71262 71810 71314 71822
rect 71598 71874 71650 71886
rect 71598 71810 71650 71822
rect 70814 71762 70866 71774
rect 3042 71710 3054 71762
rect 3106 71710 3118 71762
rect 4834 71710 4846 71762
rect 4898 71710 4910 71762
rect 72258 71710 72270 71762
rect 72322 71710 72334 71762
rect 74946 71710 74958 71762
rect 75010 71710 75022 71762
rect 76738 71710 76750 71762
rect 76802 71710 76814 71762
rect 70814 71698 70866 71710
rect 5406 71650 5458 71662
rect 2034 71598 2046 71650
rect 2098 71598 2110 71650
rect 3714 71598 3726 71650
rect 3778 71598 3790 71650
rect 5406 71586 5458 71598
rect 73502 71650 73554 71662
rect 73502 71586 73554 71598
rect 74174 71650 74226 71662
rect 75618 71598 75630 71650
rect 75682 71598 75694 71650
rect 77858 71598 77870 71650
rect 77922 71598 77934 71650
rect 74174 71586 74226 71598
rect 1344 71370 78624 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 78624 71370
rect 1344 71284 78624 71318
rect 3266 71038 3278 71090
rect 3330 71038 3342 71090
rect 74946 71038 74958 71090
rect 75010 71038 75022 71090
rect 70142 70866 70194 70878
rect 2146 70814 2158 70866
rect 2210 70814 2222 70866
rect 70142 70802 70194 70814
rect 70590 70866 70642 70878
rect 70590 70802 70642 70814
rect 70926 70866 70978 70878
rect 70926 70802 70978 70814
rect 71598 70866 71650 70878
rect 71598 70802 71650 70814
rect 71934 70866 71986 70878
rect 76290 70814 76302 70866
rect 76354 70814 76366 70866
rect 71934 70802 71986 70814
rect 3726 70754 3778 70766
rect 3726 70690 3778 70702
rect 72494 70754 72546 70766
rect 72494 70690 72546 70702
rect 72830 70754 72882 70766
rect 72830 70690 72882 70702
rect 73726 70754 73778 70766
rect 73726 70690 73778 70702
rect 74398 70754 74450 70766
rect 74398 70690 74450 70702
rect 77310 70754 77362 70766
rect 77310 70690 77362 70702
rect 1344 70586 78624 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 78624 70586
rect 1344 70500 78624 70534
rect 71262 70418 71314 70430
rect 71262 70354 71314 70366
rect 3726 70306 3778 70318
rect 1922 70254 1934 70306
rect 1986 70254 1998 70306
rect 3726 70242 3778 70254
rect 69918 70306 69970 70318
rect 76290 70254 76302 70306
rect 76354 70254 76366 70306
rect 69918 70242 69970 70254
rect 69470 70194 69522 70206
rect 69470 70130 69522 70142
rect 70254 70194 70306 70206
rect 70254 70130 70306 70142
rect 70926 70194 70978 70206
rect 70926 70130 70978 70142
rect 71710 70194 71762 70206
rect 71710 70130 71762 70142
rect 76862 70082 76914 70094
rect 3266 70030 3278 70082
rect 3330 70030 3342 70082
rect 75058 70030 75070 70082
rect 75122 70030 75134 70082
rect 76862 70018 76914 70030
rect 1344 69802 78624 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 78624 69802
rect 1344 69716 78624 69750
rect 3266 69470 3278 69522
rect 3330 69470 3342 69522
rect 72930 69470 72942 69522
rect 72994 69470 73006 69522
rect 74946 69470 74958 69522
rect 75010 69470 75022 69522
rect 4174 69298 4226 69310
rect 2258 69246 2270 69298
rect 2322 69246 2334 69298
rect 4174 69234 4226 69246
rect 69694 69298 69746 69310
rect 69694 69234 69746 69246
rect 70254 69298 70306 69310
rect 70254 69234 70306 69246
rect 70590 69298 70642 69310
rect 70590 69234 70642 69246
rect 71150 69298 71202 69310
rect 74274 69246 74286 69298
rect 74338 69246 74350 69298
rect 76290 69246 76302 69298
rect 76354 69246 76366 69298
rect 71150 69234 71202 69246
rect 3726 69186 3778 69198
rect 3726 69122 3778 69134
rect 69358 69186 69410 69198
rect 69358 69122 69410 69134
rect 77310 69186 77362 69198
rect 77310 69122 77362 69134
rect 1344 69018 78624 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 78624 69018
rect 1344 68932 78624 68966
rect 74510 68850 74562 68862
rect 74510 68786 74562 68798
rect 68574 68738 68626 68750
rect 2258 68686 2270 68738
rect 2322 68686 2334 68738
rect 3938 68686 3950 68738
rect 4002 68686 4014 68738
rect 76290 68686 76302 68738
rect 76354 68686 76366 68738
rect 68574 68674 68626 68686
rect 67118 68514 67170 68526
rect 3154 68462 3166 68514
rect 3218 68462 3230 68514
rect 5282 68462 5294 68514
rect 5346 68462 5358 68514
rect 67118 68450 67170 68462
rect 67678 68514 67730 68526
rect 67678 68450 67730 68462
rect 69918 68514 69970 68526
rect 76862 68514 76914 68526
rect 75170 68462 75182 68514
rect 75234 68462 75246 68514
rect 69918 68450 69970 68462
rect 76862 68450 76914 68462
rect 67790 68402 67842 68414
rect 67790 68338 67842 68350
rect 68686 68402 68738 68414
rect 68686 68338 68738 68350
rect 1344 68234 78624 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 78624 68234
rect 1344 68148 78624 68182
rect 3490 68014 3502 68066
rect 3554 68063 3566 68066
rect 4274 68063 4286 68066
rect 3554 68017 4286 68063
rect 3554 68014 3566 68017
rect 4274 68014 4286 68017
rect 4338 68014 4350 68066
rect 3838 67954 3890 67966
rect 3266 67902 3278 67954
rect 3330 67902 3342 67954
rect 3838 67890 3890 67902
rect 66782 67954 66834 67966
rect 66782 67890 66834 67902
rect 67902 67954 67954 67966
rect 67902 67890 67954 67902
rect 68462 67954 68514 67966
rect 68462 67890 68514 67902
rect 69470 67954 69522 67966
rect 74946 67902 74958 67954
rect 75010 67902 75022 67954
rect 69470 67890 69522 67902
rect 4174 67730 4226 67742
rect 2258 67678 2270 67730
rect 2322 67678 2334 67730
rect 4174 67666 4226 67678
rect 67230 67730 67282 67742
rect 77310 67730 77362 67742
rect 76290 67678 76302 67730
rect 76354 67678 76366 67730
rect 67230 67666 67282 67678
rect 77310 67666 77362 67678
rect 66334 67618 66386 67630
rect 66334 67554 66386 67566
rect 67342 67618 67394 67630
rect 67342 67554 67394 67566
rect 68014 67618 68066 67630
rect 68014 67554 68066 67566
rect 69358 67618 69410 67630
rect 69358 67554 69410 67566
rect 1344 67450 78624 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 78624 67450
rect 1344 67364 78624 67398
rect 68350 67282 68402 67294
rect 68350 67218 68402 67230
rect 67006 67170 67058 67182
rect 2146 67118 2158 67170
rect 2210 67118 2222 67170
rect 67006 67106 67058 67118
rect 67454 67170 67506 67182
rect 67454 67106 67506 67118
rect 69470 67170 69522 67182
rect 76290 67118 76302 67170
rect 76354 67118 76366 67170
rect 69470 67106 69522 67118
rect 3726 67058 3778 67070
rect 3726 66994 3778 67006
rect 63534 67058 63586 67070
rect 63534 66994 63586 67006
rect 65662 67058 65714 67070
rect 65662 66994 65714 67006
rect 65886 67058 65938 67070
rect 65886 66994 65938 67006
rect 68126 67058 68178 67070
rect 68798 67058 68850 67070
rect 68450 67006 68462 67058
rect 68514 67006 68526 67058
rect 68126 66994 68178 67006
rect 68798 66994 68850 67006
rect 63422 66946 63474 66958
rect 3266 66894 3278 66946
rect 3330 66894 3342 66946
rect 63422 66882 63474 66894
rect 63982 66946 64034 66958
rect 63982 66882 64034 66894
rect 65774 66946 65826 66958
rect 65774 66882 65826 66894
rect 66110 66946 66162 66958
rect 66110 66882 66162 66894
rect 68238 66946 68290 66958
rect 76862 66946 76914 66958
rect 75170 66894 75182 66946
rect 75234 66894 75246 66946
rect 68238 66882 68290 66894
rect 76862 66882 76914 66894
rect 66334 66834 66386 66846
rect 66334 66770 66386 66782
rect 66894 66834 66946 66846
rect 69358 66834 69410 66846
rect 67330 66782 67342 66834
rect 67394 66831 67406 66834
rect 67890 66831 67902 66834
rect 67394 66785 67902 66831
rect 67394 66782 67406 66785
rect 67890 66782 67902 66785
rect 67954 66782 67966 66834
rect 66894 66770 66946 66782
rect 69358 66770 69410 66782
rect 1344 66666 78624 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 78624 66666
rect 1344 66580 78624 66614
rect 68350 66498 68402 66510
rect 68350 66434 68402 66446
rect 64878 66386 64930 66398
rect 3266 66334 3278 66386
rect 3330 66334 3342 66386
rect 64878 66322 64930 66334
rect 66894 66386 66946 66398
rect 66894 66322 66946 66334
rect 68126 66386 68178 66398
rect 75058 66334 75070 66386
rect 75122 66334 75134 66386
rect 68126 66322 68178 66334
rect 66222 66274 66274 66286
rect 65874 66222 65886 66274
rect 65938 66222 65950 66274
rect 66222 66210 66274 66222
rect 66782 66274 66834 66286
rect 66782 66210 66834 66222
rect 67902 66274 67954 66286
rect 67902 66210 67954 66222
rect 63310 66162 63362 66174
rect 2034 66110 2046 66162
rect 2098 66110 2110 66162
rect 63310 66098 63362 66110
rect 63870 66162 63922 66174
rect 76290 66110 76302 66162
rect 76354 66110 76366 66162
rect 63870 66098 63922 66110
rect 3726 66050 3778 66062
rect 3726 65986 3778 65998
rect 63422 66050 63474 66062
rect 63422 65986 63474 65998
rect 65550 66050 65602 66062
rect 65550 65986 65602 65998
rect 65662 66050 65714 66062
rect 65662 65986 65714 65998
rect 65774 66050 65826 66062
rect 65774 65986 65826 65998
rect 67678 66050 67730 66062
rect 67678 65986 67730 65998
rect 67790 66050 67842 66062
rect 67790 65986 67842 65998
rect 77310 66050 77362 66062
rect 77310 65986 77362 65998
rect 1344 65882 78624 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 78624 65882
rect 1344 65796 78624 65830
rect 68238 65714 68290 65726
rect 68238 65650 68290 65662
rect 64542 65602 64594 65614
rect 1922 65550 1934 65602
rect 1986 65550 1998 65602
rect 64542 65538 64594 65550
rect 65886 65602 65938 65614
rect 76290 65550 76302 65602
rect 76354 65550 76366 65602
rect 65886 65538 65938 65550
rect 62078 65490 62130 65502
rect 66110 65490 66162 65502
rect 65762 65438 65774 65490
rect 65826 65438 65838 65490
rect 62078 65426 62130 65438
rect 66110 65426 66162 65438
rect 68014 65490 68066 65502
rect 68014 65426 68066 65438
rect 68462 65490 68514 65502
rect 68462 65426 68514 65438
rect 68686 65490 68738 65502
rect 68686 65426 68738 65438
rect 3726 65378 3778 65390
rect 3266 65326 3278 65378
rect 3330 65326 3342 65378
rect 3726 65314 3778 65326
rect 61966 65378 62018 65390
rect 61966 65314 62018 65326
rect 62526 65378 62578 65390
rect 62526 65314 62578 65326
rect 65998 65378 66050 65390
rect 65998 65314 66050 65326
rect 66782 65378 66834 65390
rect 66782 65314 66834 65326
rect 67118 65378 67170 65390
rect 67118 65314 67170 65326
rect 68126 65378 68178 65390
rect 76862 65378 76914 65390
rect 74946 65326 74958 65378
rect 75010 65326 75022 65378
rect 68126 65314 68178 65326
rect 76862 65314 76914 65326
rect 64654 65266 64706 65278
rect 64654 65202 64706 65214
rect 65438 65266 65490 65278
rect 65438 65202 65490 65214
rect 1344 65098 78624 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 78624 65098
rect 1344 65012 78624 65046
rect 66446 64818 66498 64830
rect 3266 64766 3278 64818
rect 3330 64766 3342 64818
rect 72930 64766 72942 64818
rect 72994 64766 73006 64818
rect 74946 64766 74958 64818
rect 75010 64766 75022 64818
rect 66446 64754 66498 64766
rect 4174 64706 4226 64718
rect 4174 64642 4226 64654
rect 63758 64706 63810 64718
rect 63758 64642 63810 64654
rect 64318 64706 64370 64718
rect 65774 64706 65826 64718
rect 65426 64654 65438 64706
rect 65490 64654 65502 64706
rect 64318 64642 64370 64654
rect 65774 64642 65826 64654
rect 66334 64706 66386 64718
rect 66334 64642 66386 64654
rect 68238 64706 68290 64718
rect 68238 64642 68290 64654
rect 60734 64594 60786 64606
rect 1922 64542 1934 64594
rect 1986 64542 1998 64594
rect 60734 64530 60786 64542
rect 61742 64594 61794 64606
rect 61742 64530 61794 64542
rect 67006 64594 67058 64606
rect 67006 64530 67058 64542
rect 67342 64594 67394 64606
rect 67342 64530 67394 64542
rect 69358 64594 69410 64606
rect 74274 64542 74286 64594
rect 74338 64542 74350 64594
rect 76290 64542 76302 64594
rect 76354 64542 76366 64594
rect 69358 64530 69410 64542
rect 3726 64482 3778 64494
rect 3726 64418 3778 64430
rect 61854 64482 61906 64494
rect 61854 64418 61906 64430
rect 62302 64482 62354 64494
rect 62302 64418 62354 64430
rect 64206 64482 64258 64494
rect 64206 64418 64258 64430
rect 65102 64482 65154 64494
rect 65102 64418 65154 64430
rect 65214 64482 65266 64494
rect 65214 64418 65266 64430
rect 65326 64482 65378 64494
rect 65326 64418 65378 64430
rect 68574 64482 68626 64494
rect 68574 64418 68626 64430
rect 69694 64482 69746 64494
rect 69694 64418 69746 64430
rect 77310 64482 77362 64494
rect 77310 64418 77362 64430
rect 1344 64314 78624 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 78624 64314
rect 1344 64228 78624 64262
rect 65774 64146 65826 64158
rect 65774 64082 65826 64094
rect 66334 64146 66386 64158
rect 66334 64082 66386 64094
rect 67678 64146 67730 64158
rect 67678 64082 67730 64094
rect 74510 64146 74562 64158
rect 74510 64082 74562 64094
rect 61182 64034 61234 64046
rect 2034 63982 2046 64034
rect 2098 63982 2110 64034
rect 3938 63982 3950 64034
rect 4002 63982 4014 64034
rect 61182 63970 61234 63982
rect 62526 64034 62578 64046
rect 62526 63970 62578 63982
rect 63534 64034 63586 64046
rect 63534 63970 63586 63982
rect 64654 64034 64706 64046
rect 76290 63982 76302 64034
rect 76354 63982 76366 64034
rect 64654 63970 64706 63982
rect 61070 63922 61122 63934
rect 61070 63858 61122 63870
rect 61630 63922 61682 63934
rect 63310 63922 63362 63934
rect 66670 63922 66722 63934
rect 62290 63870 62302 63922
rect 62354 63870 62366 63922
rect 65538 63870 65550 63922
rect 65602 63870 65614 63922
rect 61630 63858 61682 63870
rect 63310 63858 63362 63870
rect 66670 63858 66722 63870
rect 67342 63922 67394 63934
rect 67342 63858 67394 63870
rect 76862 63922 76914 63934
rect 76862 63858 76914 63870
rect 63422 63810 63474 63822
rect 3266 63758 3278 63810
rect 3330 63758 3342 63810
rect 5282 63758 5294 63810
rect 5346 63758 5358 63810
rect 63422 63746 63474 63758
rect 63758 63810 63810 63822
rect 75170 63758 75182 63810
rect 75234 63758 75246 63810
rect 63758 63746 63810 63758
rect 63982 63698 64034 63710
rect 63982 63634 64034 63646
rect 64542 63698 64594 63710
rect 64542 63634 64594 63646
rect 1344 63530 78624 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 78624 63530
rect 1344 63444 78624 63478
rect 63870 63362 63922 63374
rect 63870 63298 63922 63310
rect 3838 63250 3890 63262
rect 3266 63198 3278 63250
rect 3330 63198 3342 63250
rect 3838 63186 3890 63198
rect 59278 63250 59330 63262
rect 59278 63186 59330 63198
rect 59838 63250 59890 63262
rect 59838 63186 59890 63198
rect 63646 63250 63698 63262
rect 63646 63186 63698 63198
rect 64990 63250 65042 63262
rect 64990 63186 65042 63198
rect 65326 63250 65378 63262
rect 74946 63198 74958 63250
rect 75010 63198 75022 63250
rect 65326 63186 65378 63198
rect 63198 63138 63250 63150
rect 63198 63074 63250 63086
rect 61406 63026 61458 63038
rect 2146 62974 2158 63026
rect 2210 62974 2222 63026
rect 61406 62962 61458 62974
rect 61966 63026 62018 63038
rect 76290 62974 76302 63026
rect 76354 62974 76366 63026
rect 61966 62962 62018 62974
rect 4174 62914 4226 62926
rect 4174 62850 4226 62862
rect 59390 62914 59442 62926
rect 59390 62850 59442 62862
rect 61518 62914 61570 62926
rect 61518 62850 61570 62862
rect 63310 62914 63362 62926
rect 63310 62850 63362 62862
rect 63422 62914 63474 62926
rect 63422 62850 63474 62862
rect 65998 62914 66050 62926
rect 65998 62850 66050 62862
rect 67006 62914 67058 62926
rect 67006 62850 67058 62862
rect 77310 62914 77362 62926
rect 77310 62850 77362 62862
rect 1344 62746 78624 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 78624 62746
rect 1344 62660 78624 62694
rect 62750 62578 62802 62590
rect 62750 62514 62802 62526
rect 62974 62578 63026 62590
rect 62974 62514 63026 62526
rect 63758 62578 63810 62590
rect 63758 62514 63810 62526
rect 3726 62466 3778 62478
rect 1922 62414 1934 62466
rect 1986 62414 1998 62466
rect 3726 62402 3778 62414
rect 61630 62466 61682 62478
rect 61630 62402 61682 62414
rect 68238 62466 68290 62478
rect 68238 62402 68290 62414
rect 68686 62466 68738 62478
rect 76290 62414 76302 62466
rect 76354 62414 76366 62466
rect 68686 62402 68738 62414
rect 59726 62354 59778 62366
rect 59726 62290 59778 62302
rect 61182 62354 61234 62366
rect 61182 62290 61234 62302
rect 62526 62354 62578 62366
rect 62526 62290 62578 62302
rect 63982 62354 64034 62366
rect 64082 62302 64094 62354
rect 64146 62302 64158 62354
rect 63982 62290 64034 62302
rect 59614 62242 59666 62254
rect 3266 62190 3278 62242
rect 3330 62190 3342 62242
rect 59614 62178 59666 62190
rect 60174 62242 60226 62254
rect 60174 62178 60226 62190
rect 61742 62242 61794 62254
rect 61742 62178 61794 62190
rect 62302 62242 62354 62254
rect 62302 62178 62354 62190
rect 62862 62242 62914 62254
rect 62862 62178 62914 62190
rect 63870 62242 63922 62254
rect 63870 62178 63922 62190
rect 64430 62242 64482 62254
rect 64430 62178 64482 62190
rect 68126 62242 68178 62254
rect 76862 62242 76914 62254
rect 75058 62190 75070 62242
rect 75122 62190 75134 62242
rect 68126 62178 68178 62190
rect 76862 62178 76914 62190
rect 1344 61962 78624 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 78624 61962
rect 1344 61876 78624 61910
rect 3266 61630 3278 61682
rect 3330 61630 3342 61682
rect 74946 61630 74958 61682
rect 75010 61630 75022 61682
rect 60286 61458 60338 61470
rect 2034 61406 2046 61458
rect 2098 61406 2110 61458
rect 60286 61394 60338 61406
rect 61518 61458 61570 61470
rect 61518 61394 61570 61406
rect 63646 61458 63698 61470
rect 76290 61406 76302 61458
rect 76354 61406 76366 61458
rect 63646 61394 63698 61406
rect 3726 61346 3778 61358
rect 3726 61282 3778 61294
rect 59054 61346 59106 61358
rect 59054 61282 59106 61294
rect 59838 61346 59890 61358
rect 59838 61282 59890 61294
rect 60398 61346 60450 61358
rect 60398 61282 60450 61294
rect 61630 61346 61682 61358
rect 61630 61282 61682 61294
rect 62190 61346 62242 61358
rect 62190 61282 62242 61294
rect 62750 61346 62802 61358
rect 62750 61282 62802 61294
rect 63310 61346 63362 61358
rect 63310 61282 63362 61294
rect 77310 61346 77362 61358
rect 77310 61282 77362 61294
rect 1344 61178 78624 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 78624 61178
rect 1344 61092 78624 61126
rect 58494 61010 58546 61022
rect 58494 60946 58546 60958
rect 62414 61010 62466 61022
rect 62414 60946 62466 60958
rect 59726 60898 59778 60910
rect 2146 60846 2158 60898
rect 2210 60846 2222 60898
rect 59726 60834 59778 60846
rect 60734 60898 60786 60910
rect 60734 60834 60786 60846
rect 62638 60898 62690 60910
rect 76290 60846 76302 60898
rect 76354 60846 76366 60898
rect 62638 60834 62690 60846
rect 57598 60786 57650 60798
rect 57598 60722 57650 60734
rect 59390 60786 59442 60798
rect 59390 60722 59442 60734
rect 60958 60786 61010 60798
rect 60958 60722 61010 60734
rect 61966 60786 62018 60798
rect 61966 60722 62018 60734
rect 3726 60674 3778 60686
rect 3266 60622 3278 60674
rect 3330 60622 3342 60674
rect 3726 60610 3778 60622
rect 57486 60674 57538 60686
rect 57486 60610 57538 60622
rect 58046 60674 58098 60686
rect 58046 60610 58098 60622
rect 60846 60674 60898 60686
rect 60846 60610 60898 60622
rect 61182 60674 61234 60686
rect 61182 60610 61234 60622
rect 62190 60674 62242 60686
rect 62190 60610 62242 60622
rect 62526 60674 62578 60686
rect 62526 60610 62578 60622
rect 64542 60674 64594 60686
rect 64542 60610 64594 60622
rect 65326 60674 65378 60686
rect 76862 60674 76914 60686
rect 74946 60622 74958 60674
rect 75010 60622 75022 60674
rect 65326 60610 65378 60622
rect 76862 60610 76914 60622
rect 61406 60562 61458 60574
rect 61406 60498 61458 60510
rect 64430 60562 64482 60574
rect 64430 60498 64482 60510
rect 1344 60394 78624 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 78624 60394
rect 1344 60308 78624 60342
rect 58830 60114 58882 60126
rect 3266 60062 3278 60114
rect 3330 60062 3342 60114
rect 58830 60050 58882 60062
rect 60398 60114 60450 60126
rect 60398 60050 60450 60062
rect 66558 60114 66610 60126
rect 66558 60050 66610 60062
rect 67118 60114 67170 60126
rect 72930 60062 72942 60114
rect 72994 60062 73006 60114
rect 74946 60062 74958 60114
rect 75010 60062 75022 60114
rect 67118 60050 67170 60062
rect 58046 60002 58098 60014
rect 58046 59938 58098 59950
rect 59950 60002 60002 60014
rect 59950 59938 60002 59950
rect 60622 60002 60674 60014
rect 60622 59938 60674 59950
rect 66446 60002 66498 60014
rect 66446 59938 66498 59950
rect 56814 59890 56866 59902
rect 2258 59838 2270 59890
rect 2322 59838 2334 59890
rect 56814 59826 56866 59838
rect 57150 59890 57202 59902
rect 57150 59826 57202 59838
rect 58158 59890 58210 59902
rect 58158 59826 58210 59838
rect 60174 59890 60226 59902
rect 60174 59826 60226 59838
rect 61518 59890 61570 59902
rect 61518 59826 61570 59838
rect 62078 59890 62130 59902
rect 74274 59838 74286 59890
rect 74338 59838 74350 59890
rect 76290 59838 76302 59890
rect 76354 59838 76366 59890
rect 62078 59826 62130 59838
rect 3726 59778 3778 59790
rect 3726 59714 3778 59726
rect 4174 59778 4226 59790
rect 4174 59714 4226 59726
rect 56366 59778 56418 59790
rect 56366 59714 56418 59726
rect 58942 59778 58994 59790
rect 58942 59714 58994 59726
rect 60062 59778 60114 59790
rect 60062 59714 60114 59726
rect 61406 59778 61458 59790
rect 61406 59714 61458 59726
rect 77310 59778 77362 59790
rect 77310 59714 77362 59726
rect 1344 59610 78624 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 78624 59610
rect 1344 59524 78624 59558
rect 57822 59442 57874 59454
rect 57822 59378 57874 59390
rect 59614 59442 59666 59454
rect 59614 59378 59666 59390
rect 59838 59442 59890 59454
rect 59838 59378 59890 59390
rect 61070 59442 61122 59454
rect 61070 59378 61122 59390
rect 74510 59442 74562 59454
rect 74510 59378 74562 59390
rect 1922 59278 1934 59330
rect 1986 59278 1998 59330
rect 3938 59278 3950 59330
rect 4002 59278 4014 59330
rect 76290 59278 76302 59330
rect 76354 59278 76366 59330
rect 58382 59218 58434 59230
rect 58382 59154 58434 59166
rect 58942 59218 58994 59230
rect 58942 59154 58994 59166
rect 60286 59218 60338 59230
rect 61282 59166 61294 59218
rect 61346 59166 61358 59218
rect 60286 59154 60338 59166
rect 59726 59106 59778 59118
rect 3266 59054 3278 59106
rect 3330 59054 3342 59106
rect 5282 59054 5294 59106
rect 5346 59054 5358 59106
rect 59726 59042 59778 59054
rect 60062 59106 60114 59118
rect 60062 59042 60114 59054
rect 61854 59106 61906 59118
rect 76862 59106 76914 59118
rect 75170 59054 75182 59106
rect 75234 59054 75246 59106
rect 61854 59042 61906 59054
rect 76862 59042 76914 59054
rect 58494 58994 58546 59006
rect 58494 58930 58546 58942
rect 1344 58826 78624 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 78624 58826
rect 1344 58740 78624 58774
rect 58606 58658 58658 58670
rect 58606 58594 58658 58606
rect 3838 58546 3890 58558
rect 3266 58494 3278 58546
rect 3330 58494 3342 58546
rect 75058 58494 75070 58546
rect 75122 58494 75134 58546
rect 3838 58482 3890 58494
rect 57262 58434 57314 58446
rect 57262 58370 57314 58382
rect 58158 58434 58210 58446
rect 58258 58382 58270 58434
rect 58322 58382 58334 58434
rect 58158 58370 58210 58382
rect 57150 58322 57202 58334
rect 2034 58270 2046 58322
rect 2098 58270 2110 58322
rect 57150 58258 57202 58270
rect 59278 58322 59330 58334
rect 76290 58270 76302 58322
rect 76354 58270 76366 58322
rect 59278 58258 59330 58270
rect 4174 58210 4226 58222
rect 4174 58146 4226 58158
rect 56702 58210 56754 58222
rect 56702 58146 56754 58158
rect 57934 58210 57986 58222
rect 57934 58146 57986 58158
rect 58046 58210 58098 58222
rect 58046 58146 58098 58158
rect 59166 58210 59218 58222
rect 59166 58146 59218 58158
rect 59838 58210 59890 58222
rect 59838 58146 59890 58158
rect 77310 58210 77362 58222
rect 77310 58146 77362 58158
rect 1344 58042 78624 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 78624 58042
rect 1344 57956 78624 57990
rect 57822 57874 57874 57886
rect 57822 57810 57874 57822
rect 63310 57874 63362 57886
rect 63310 57810 63362 57822
rect 62862 57762 62914 57774
rect 1922 57710 1934 57762
rect 1986 57710 1998 57762
rect 76290 57710 76302 57762
rect 76354 57710 76366 57762
rect 62862 57698 62914 57710
rect 54574 57650 54626 57662
rect 54574 57586 54626 57598
rect 55134 57650 55186 57662
rect 55134 57586 55186 57598
rect 56142 57650 56194 57662
rect 56142 57586 56194 57598
rect 58046 57650 58098 57662
rect 58046 57586 58098 57598
rect 58270 57650 58322 57662
rect 58270 57586 58322 57598
rect 58494 57650 58546 57662
rect 58494 57586 58546 57598
rect 3726 57538 3778 57550
rect 3154 57486 3166 57538
rect 3218 57486 3230 57538
rect 3726 57474 3778 57486
rect 56030 57538 56082 57550
rect 56030 57474 56082 57486
rect 56590 57538 56642 57550
rect 56590 57474 56642 57486
rect 57934 57538 57986 57550
rect 76862 57538 76914 57550
rect 74946 57486 74958 57538
rect 75010 57486 75022 57538
rect 57934 57474 57986 57486
rect 76862 57474 76914 57486
rect 55246 57426 55298 57438
rect 55246 57362 55298 57374
rect 62750 57426 62802 57438
rect 62750 57362 62802 57374
rect 1344 57258 78624 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 78624 57258
rect 1344 57172 78624 57206
rect 58046 57090 58098 57102
rect 58046 57026 58098 57038
rect 57822 56978 57874 56990
rect 3266 56926 3278 56978
rect 3330 56926 3342 56978
rect 74946 56926 74958 56978
rect 75010 56926 75022 56978
rect 57822 56914 57874 56926
rect 57598 56866 57650 56878
rect 57598 56802 57650 56814
rect 3726 56754 3778 56766
rect 2258 56702 2270 56754
rect 2322 56702 2334 56754
rect 3726 56690 3778 56702
rect 56142 56754 56194 56766
rect 56142 56690 56194 56702
rect 56590 56754 56642 56766
rect 56590 56690 56642 56702
rect 58942 56754 58994 56766
rect 58942 56690 58994 56702
rect 59502 56754 59554 56766
rect 76290 56702 76302 56754
rect 76354 56702 76366 56754
rect 59502 56690 59554 56702
rect 56702 56642 56754 56654
rect 56702 56578 56754 56590
rect 57374 56642 57426 56654
rect 57374 56578 57426 56590
rect 57486 56642 57538 56654
rect 57486 56578 57538 56590
rect 58830 56642 58882 56654
rect 58830 56578 58882 56590
rect 77310 56642 77362 56654
rect 77310 56578 77362 56590
rect 1344 56474 78624 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 78624 56474
rect 1344 56388 78624 56422
rect 57598 56306 57650 56318
rect 57598 56242 57650 56254
rect 57822 56306 57874 56318
rect 57822 56242 57874 56254
rect 3726 56194 3778 56206
rect 76862 56194 76914 56206
rect 2258 56142 2270 56194
rect 2322 56142 2334 56194
rect 76290 56142 76302 56194
rect 76354 56142 76366 56194
rect 3726 56130 3778 56142
rect 76862 56130 76914 56142
rect 53230 56082 53282 56094
rect 53230 56018 53282 56030
rect 55358 56082 55410 56094
rect 55358 56018 55410 56030
rect 55582 56082 55634 56094
rect 56702 56082 56754 56094
rect 55682 56030 55694 56082
rect 55746 56030 55758 56082
rect 55582 56018 55634 56030
rect 56702 56018 56754 56030
rect 58046 56082 58098 56094
rect 58046 56018 58098 56030
rect 58270 56082 58322 56094
rect 58270 56018 58322 56030
rect 53118 55970 53170 55982
rect 3266 55918 3278 55970
rect 3330 55918 3342 55970
rect 53118 55906 53170 55918
rect 53678 55970 53730 55982
rect 53678 55906 53730 55918
rect 54798 55970 54850 55982
rect 54798 55906 54850 55918
rect 55470 55970 55522 55982
rect 55470 55906 55522 55918
rect 57710 55970 57762 55982
rect 75058 55918 75070 55970
rect 75122 55918 75134 55970
rect 57710 55906 57762 55918
rect 56030 55858 56082 55870
rect 56030 55794 56082 55806
rect 56590 55858 56642 55870
rect 56590 55794 56642 55806
rect 1344 55690 78624 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 78624 55690
rect 1344 55604 78624 55638
rect 57474 55470 57486 55522
rect 57538 55519 57550 55522
rect 57698 55519 57710 55522
rect 57538 55473 57710 55519
rect 57538 55470 57550 55473
rect 57698 55470 57710 55473
rect 57762 55470 57774 55522
rect 55694 55410 55746 55422
rect 3266 55358 3278 55410
rect 3330 55358 3342 55410
rect 55694 55346 55746 55358
rect 57822 55410 57874 55422
rect 75170 55358 75182 55410
rect 75234 55358 75246 55410
rect 57822 55346 57874 55358
rect 55246 55298 55298 55310
rect 54226 55246 54238 55298
rect 54290 55246 54302 55298
rect 55246 55234 55298 55246
rect 55918 55298 55970 55310
rect 55918 55234 55970 55246
rect 50654 55186 50706 55198
rect 2034 55134 2046 55186
rect 2098 55134 2110 55186
rect 50654 55122 50706 55134
rect 50766 55186 50818 55198
rect 50766 55122 50818 55134
rect 54462 55186 54514 55198
rect 54462 55122 54514 55134
rect 55470 55186 55522 55198
rect 55470 55122 55522 55134
rect 56926 55186 56978 55198
rect 56926 55122 56978 55134
rect 57262 55186 57314 55198
rect 76290 55134 76302 55186
rect 76354 55134 76366 55186
rect 57262 55122 57314 55134
rect 3726 55074 3778 55086
rect 3726 55010 3778 55022
rect 51214 55074 51266 55086
rect 51214 55010 51266 55022
rect 53678 55074 53730 55086
rect 53678 55010 53730 55022
rect 55358 55074 55410 55086
rect 55358 55010 55410 55022
rect 56366 55074 56418 55086
rect 56366 55010 56418 55022
rect 77310 55074 77362 55086
rect 77310 55010 77362 55022
rect 1344 54906 78624 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 78624 54906
rect 1344 54820 78624 54854
rect 3726 54738 3778 54750
rect 3726 54674 3778 54686
rect 56590 54738 56642 54750
rect 56590 54674 56642 54686
rect 52222 54626 52274 54638
rect 2146 54574 2158 54626
rect 2210 54574 2222 54626
rect 52222 54562 52274 54574
rect 53902 54626 53954 54638
rect 53902 54562 53954 54574
rect 54910 54626 54962 54638
rect 54910 54562 54962 54574
rect 56030 54626 56082 54638
rect 56030 54562 56082 54574
rect 56702 54626 56754 54638
rect 56702 54562 56754 54574
rect 57374 54626 57426 54638
rect 76290 54574 76302 54626
rect 76354 54574 76366 54626
rect 57374 54562 57426 54574
rect 51550 54514 51602 54526
rect 51550 54450 51602 54462
rect 52110 54514 52162 54526
rect 52110 54450 52162 54462
rect 54686 54514 54738 54526
rect 55010 54462 55022 54514
rect 55074 54462 55086 54514
rect 54686 54450 54738 54462
rect 52782 54402 52834 54414
rect 3266 54350 3278 54402
rect 3330 54350 3342 54402
rect 52782 54338 52834 54350
rect 53342 54402 53394 54414
rect 53342 54338 53394 54350
rect 54798 54402 54850 54414
rect 76862 54402 76914 54414
rect 75058 54350 75070 54402
rect 75122 54350 75134 54402
rect 54798 54338 54850 54350
rect 76862 54338 76914 54350
rect 52894 54290 52946 54302
rect 52894 54226 52946 54238
rect 54014 54290 54066 54302
rect 54014 54226 54066 54238
rect 55358 54290 55410 54302
rect 55358 54226 55410 54238
rect 55918 54290 55970 54302
rect 55918 54226 55970 54238
rect 1344 54122 78624 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 78624 54122
rect 1344 54036 78624 54070
rect 54238 53954 54290 53966
rect 56130 53902 56142 53954
rect 56194 53951 56206 53954
rect 56466 53951 56478 53954
rect 56194 53905 56478 53951
rect 56194 53902 56206 53905
rect 56466 53902 56478 53905
rect 56530 53902 56542 53954
rect 54238 53890 54290 53902
rect 54462 53842 54514 53854
rect 3266 53790 3278 53842
rect 3330 53790 3342 53842
rect 54462 53778 54514 53790
rect 56478 53842 56530 53854
rect 74946 53790 74958 53842
rect 75010 53790 75022 53842
rect 56478 53778 56530 53790
rect 52222 53730 52274 53742
rect 52222 53666 52274 53678
rect 54686 53730 54738 53742
rect 54686 53666 54738 53678
rect 53566 53618 53618 53630
rect 2034 53566 2046 53618
rect 2098 53566 2110 53618
rect 53566 53554 53618 53566
rect 55918 53618 55970 53630
rect 55918 53554 55970 53566
rect 57038 53618 57090 53630
rect 57038 53554 57090 53566
rect 57374 53618 57426 53630
rect 76290 53566 76302 53618
rect 76354 53566 76366 53618
rect 57374 53554 57426 53566
rect 3726 53506 3778 53518
rect 3726 53442 3778 53454
rect 53454 53506 53506 53518
rect 53454 53442 53506 53454
rect 54798 53506 54850 53518
rect 54798 53442 54850 53454
rect 54910 53506 54962 53518
rect 54910 53442 54962 53454
rect 55582 53506 55634 53518
rect 55582 53442 55634 53454
rect 77310 53506 77362 53518
rect 77310 53442 77362 53454
rect 1344 53338 78624 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 78624 53338
rect 1344 53252 78624 53286
rect 58046 53170 58098 53182
rect 58046 53106 58098 53118
rect 51998 53058 52050 53070
rect 1922 53006 1934 53058
rect 1986 53006 1998 53058
rect 51998 52994 52050 53006
rect 57598 53058 57650 53070
rect 76290 53006 76302 53058
rect 76354 53006 76366 53058
rect 57598 52994 57650 53006
rect 47742 52946 47794 52958
rect 47742 52882 47794 52894
rect 48302 52946 48354 52958
rect 48302 52882 48354 52894
rect 50542 52946 50594 52958
rect 52894 52946 52946 52958
rect 51762 52894 51774 52946
rect 51826 52894 51838 52946
rect 50542 52882 50594 52894
rect 52894 52882 52946 52894
rect 53118 52946 53170 52958
rect 53118 52882 53170 52894
rect 53566 52946 53618 52958
rect 53566 52882 53618 52894
rect 3726 52834 3778 52846
rect 3266 52782 3278 52834
rect 3330 52782 3342 52834
rect 3726 52770 3778 52782
rect 50430 52834 50482 52846
rect 50430 52770 50482 52782
rect 50990 52834 51042 52846
rect 50990 52770 51042 52782
rect 53006 52834 53058 52846
rect 53006 52770 53058 52782
rect 53342 52834 53394 52846
rect 53342 52770 53394 52782
rect 54126 52834 54178 52846
rect 54126 52770 54178 52782
rect 56702 52834 56754 52846
rect 76862 52834 76914 52846
rect 75058 52782 75070 52834
rect 75122 52782 75134 52834
rect 56702 52770 56754 52782
rect 76862 52770 76914 52782
rect 48414 52722 48466 52734
rect 48414 52658 48466 52670
rect 57486 52722 57538 52734
rect 57486 52658 57538 52670
rect 1344 52554 78624 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 78624 52554
rect 1344 52468 78624 52502
rect 54238 52386 54290 52398
rect 54238 52322 54290 52334
rect 60510 52386 60562 52398
rect 60510 52322 60562 52334
rect 48302 52274 48354 52286
rect 3266 52222 3278 52274
rect 3330 52222 3342 52274
rect 48302 52210 48354 52222
rect 48862 52274 48914 52286
rect 48862 52210 48914 52222
rect 49534 52274 49586 52286
rect 49534 52210 49586 52222
rect 51326 52274 51378 52286
rect 51326 52210 51378 52222
rect 52670 52274 52722 52286
rect 52670 52210 52722 52222
rect 54014 52274 54066 52286
rect 54014 52210 54066 52222
rect 59278 52274 59330 52286
rect 59278 52210 59330 52222
rect 60622 52274 60674 52286
rect 60622 52210 60674 52222
rect 61406 52274 61458 52286
rect 75170 52222 75182 52274
rect 75234 52222 75246 52274
rect 61406 52210 61458 52222
rect 3726 52162 3778 52174
rect 3726 52098 3778 52110
rect 50878 52162 50930 52174
rect 59390 52162 59442 52174
rect 52322 52110 52334 52162
rect 52386 52110 52398 52162
rect 56130 52110 56142 52162
rect 56194 52110 56206 52162
rect 50878 52098 50930 52110
rect 59390 52098 59442 52110
rect 59950 52162 60002 52174
rect 59950 52098 60002 52110
rect 77310 52162 77362 52174
rect 77310 52098 77362 52110
rect 56366 52050 56418 52062
rect 2034 51998 2046 52050
rect 2098 51998 2110 52050
rect 56366 51986 56418 51998
rect 56926 52050 56978 52062
rect 56926 51986 56978 51998
rect 57262 52050 57314 52062
rect 76290 51998 76302 52050
rect 76354 51998 76366 52050
rect 57262 51986 57314 51998
rect 48414 51938 48466 51950
rect 48414 51874 48466 51886
rect 49646 51938 49698 51950
rect 49646 51874 49698 51886
rect 50542 51938 50594 51950
rect 50542 51874 50594 51886
rect 51998 51938 52050 51950
rect 51998 51874 52050 51886
rect 52110 51938 52162 51950
rect 52110 51874 52162 51886
rect 52222 51938 52274 51950
rect 52222 51874 52274 51886
rect 53566 51938 53618 51950
rect 53566 51874 53618 51886
rect 53678 51938 53730 51950
rect 53678 51874 53730 51886
rect 53790 51938 53842 51950
rect 53790 51874 53842 51886
rect 55582 51938 55634 51950
rect 55582 51874 55634 51886
rect 1344 51770 78624 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 78624 51770
rect 1344 51684 78624 51718
rect 49534 51602 49586 51614
rect 49534 51538 49586 51550
rect 51886 51602 51938 51614
rect 51886 51538 51938 51550
rect 53342 51602 53394 51614
rect 53342 51538 53394 51550
rect 52110 51490 52162 51502
rect 2146 51438 2158 51490
rect 2210 51438 2222 51490
rect 52110 51426 52162 51438
rect 53678 51490 53730 51502
rect 53678 51426 53730 51438
rect 56590 51490 56642 51502
rect 76290 51438 76302 51490
rect 76354 51438 76366 51490
rect 56590 51426 56642 51438
rect 52334 51378 52386 51390
rect 52334 51314 52386 51326
rect 52558 51378 52610 51390
rect 52558 51314 52610 51326
rect 56254 51378 56306 51390
rect 56254 51314 56306 51326
rect 3726 51266 3778 51278
rect 3266 51214 3278 51266
rect 3330 51214 3342 51266
rect 3726 51202 3778 51214
rect 51998 51266 52050 51278
rect 51998 51202 52050 51214
rect 55694 51266 55746 51278
rect 76862 51266 76914 51278
rect 75058 51214 75070 51266
rect 75122 51214 75134 51266
rect 55694 51202 55746 51214
rect 76862 51202 76914 51214
rect 1344 50986 78624 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 78624 50986
rect 1344 50900 78624 50934
rect 48974 50706 49026 50718
rect 3266 50654 3278 50706
rect 3330 50654 3342 50706
rect 48974 50642 49026 50654
rect 49422 50706 49474 50718
rect 49422 50642 49474 50654
rect 50542 50706 50594 50718
rect 50542 50642 50594 50654
rect 50878 50706 50930 50718
rect 50878 50642 50930 50654
rect 72158 50706 72210 50718
rect 72158 50642 72210 50654
rect 72606 50706 72658 50718
rect 72606 50642 72658 50654
rect 73502 50706 73554 50718
rect 73502 50642 73554 50654
rect 74062 50706 74114 50718
rect 74946 50654 74958 50706
rect 75010 50654 75022 50706
rect 74062 50642 74114 50654
rect 3726 50594 3778 50606
rect 3726 50530 3778 50542
rect 51102 50594 51154 50606
rect 51102 50530 51154 50542
rect 51662 50594 51714 50606
rect 51662 50530 51714 50542
rect 51774 50594 51826 50606
rect 51774 50530 51826 50542
rect 52334 50594 52386 50606
rect 53666 50542 53678 50594
rect 53730 50542 53742 50594
rect 52334 50530 52386 50542
rect 49534 50482 49586 50494
rect 1922 50430 1934 50482
rect 1986 50430 1998 50482
rect 49534 50418 49586 50430
rect 50430 50482 50482 50494
rect 50430 50418 50482 50430
rect 50654 50482 50706 50494
rect 77310 50482 77362 50494
rect 76290 50430 76302 50482
rect 76354 50430 76366 50482
rect 50654 50418 50706 50430
rect 77310 50418 77362 50430
rect 53454 50370 53506 50382
rect 53454 50306 53506 50318
rect 72718 50370 72770 50382
rect 72718 50306 72770 50318
rect 73390 50370 73442 50382
rect 73390 50306 73442 50318
rect 1344 50202 78624 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 78624 50202
rect 1344 50116 78624 50150
rect 50206 50034 50258 50046
rect 50206 49970 50258 49982
rect 73838 50034 73890 50046
rect 73838 49970 73890 49982
rect 46734 49922 46786 49934
rect 2034 49870 2046 49922
rect 2098 49870 2110 49922
rect 46734 49858 46786 49870
rect 50430 49922 50482 49934
rect 76290 49870 76302 49922
rect 76354 49870 76366 49922
rect 50430 49858 50482 49870
rect 46622 49810 46674 49822
rect 46622 49746 46674 49758
rect 47182 49810 47234 49822
rect 47182 49746 47234 49758
rect 50654 49810 50706 49822
rect 50654 49746 50706 49758
rect 73390 49810 73442 49822
rect 73390 49746 73442 49758
rect 73614 49810 73666 49822
rect 73614 49746 73666 49758
rect 74062 49810 74114 49822
rect 74062 49746 74114 49758
rect 3726 49698 3778 49710
rect 3266 49646 3278 49698
rect 3330 49646 3342 49698
rect 3726 49634 3778 49646
rect 48190 49698 48242 49710
rect 48190 49634 48242 49646
rect 48750 49698 48802 49710
rect 48750 49634 48802 49646
rect 50318 49698 50370 49710
rect 50318 49634 50370 49646
rect 51550 49698 51602 49710
rect 51550 49634 51602 49646
rect 51998 49698 52050 49710
rect 51998 49634 52050 49646
rect 72606 49698 72658 49710
rect 72606 49634 72658 49646
rect 73950 49698 74002 49710
rect 76862 49698 76914 49710
rect 75170 49646 75182 49698
rect 75234 49646 75246 49698
rect 73950 49634 74002 49646
rect 76862 49634 76914 49646
rect 48302 49586 48354 49598
rect 48302 49522 48354 49534
rect 50878 49586 50930 49598
rect 50878 49522 50930 49534
rect 51438 49586 51490 49598
rect 51438 49522 51490 49534
rect 1344 49418 78624 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 78624 49418
rect 1344 49332 78624 49366
rect 48078 49138 48130 49150
rect 3266 49086 3278 49138
rect 3330 49086 3342 49138
rect 48078 49074 48130 49086
rect 49422 49138 49474 49150
rect 49422 49074 49474 49086
rect 50654 49138 50706 49150
rect 50654 49074 50706 49086
rect 51214 49138 51266 49150
rect 51214 49074 51266 49086
rect 66670 49138 66722 49150
rect 66670 49074 66722 49086
rect 67118 49138 67170 49150
rect 67118 49074 67170 49086
rect 68350 49138 68402 49150
rect 68350 49074 68402 49086
rect 69470 49138 69522 49150
rect 74946 49086 74958 49138
rect 75010 49086 75022 49138
rect 69470 49074 69522 49086
rect 49198 49026 49250 49038
rect 49198 48962 49250 48974
rect 49870 49026 49922 49038
rect 49870 48962 49922 48974
rect 68574 49026 68626 49038
rect 68574 48962 68626 48974
rect 69358 49026 69410 49038
rect 69358 48962 69410 48974
rect 70030 48914 70082 48926
rect 1922 48862 1934 48914
rect 1986 48862 1998 48914
rect 76290 48862 76302 48914
rect 76354 48862 76366 48914
rect 70030 48850 70082 48862
rect 3838 48802 3890 48814
rect 3838 48738 3890 48750
rect 4174 48802 4226 48814
rect 4174 48738 4226 48750
rect 49646 48802 49698 48814
rect 49646 48738 49698 48750
rect 49758 48802 49810 48814
rect 49758 48738 49810 48750
rect 50542 48802 50594 48814
rect 50542 48738 50594 48750
rect 67230 48802 67282 48814
rect 67230 48738 67282 48750
rect 67902 48802 67954 48814
rect 67902 48738 67954 48750
rect 68014 48802 68066 48814
rect 68014 48738 68066 48750
rect 68126 48802 68178 48814
rect 68126 48738 68178 48750
rect 73054 48802 73106 48814
rect 73054 48738 73106 48750
rect 77310 48802 77362 48814
rect 77310 48738 77362 48750
rect 1344 48634 78624 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 78624 48634
rect 1344 48548 78624 48582
rect 48526 48466 48578 48478
rect 48526 48402 48578 48414
rect 49646 48466 49698 48478
rect 49646 48402 49698 48414
rect 68910 48466 68962 48478
rect 68910 48402 68962 48414
rect 48414 48354 48466 48366
rect 48414 48290 48466 48302
rect 49870 48242 49922 48254
rect 3042 48190 3054 48242
rect 3106 48190 3118 48242
rect 4834 48190 4846 48242
rect 4898 48190 4910 48242
rect 49870 48178 49922 48190
rect 50094 48242 50146 48254
rect 50094 48178 50146 48190
rect 50318 48242 50370 48254
rect 74946 48190 74958 48242
rect 75010 48190 75022 48242
rect 76738 48190 76750 48242
rect 76802 48190 76814 48242
rect 50318 48178 50370 48190
rect 5406 48130 5458 48142
rect 2034 48078 2046 48130
rect 2098 48078 2110 48130
rect 3714 48078 3726 48130
rect 3778 48078 3790 48130
rect 5406 48066 5458 48078
rect 47742 48130 47794 48142
rect 47742 48066 47794 48078
rect 49758 48130 49810 48142
rect 49758 48066 49810 48078
rect 74510 48130 74562 48142
rect 75954 48078 75966 48130
rect 76018 48078 76030 48130
rect 77858 48078 77870 48130
rect 77922 48078 77934 48130
rect 74510 48066 74562 48078
rect 1344 47850 78624 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 78624 47850
rect 1344 47764 78624 47798
rect 49534 47682 49586 47694
rect 49534 47618 49586 47630
rect 3042 47406 3054 47458
rect 3106 47406 3118 47458
rect 74946 47406 74958 47458
rect 75010 47406 75022 47458
rect 47070 47346 47122 47358
rect 1922 47294 1934 47346
rect 1986 47294 1998 47346
rect 47070 47282 47122 47294
rect 47406 47346 47458 47358
rect 47406 47282 47458 47294
rect 48078 47346 48130 47358
rect 48078 47282 48130 47294
rect 49646 47346 49698 47358
rect 49646 47282 49698 47294
rect 50206 47346 50258 47358
rect 76066 47294 76078 47346
rect 76130 47294 76142 47346
rect 50206 47282 50258 47294
rect 3502 47234 3554 47246
rect 3502 47170 3554 47182
rect 48414 47234 48466 47246
rect 48414 47170 48466 47182
rect 48862 47234 48914 47246
rect 48862 47170 48914 47182
rect 74398 47234 74450 47246
rect 74398 47170 74450 47182
rect 77198 47234 77250 47246
rect 77198 47170 77250 47182
rect 1344 47066 78624 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 78624 47066
rect 1344 46980 78624 47014
rect 46398 46786 46450 46798
rect 46398 46722 46450 46734
rect 47742 46786 47794 46798
rect 47742 46722 47794 46734
rect 45950 46674 46002 46686
rect 3042 46622 3054 46674
rect 3106 46622 3118 46674
rect 45950 46610 46002 46622
rect 46734 46674 46786 46686
rect 47506 46622 47518 46674
rect 47570 46622 47582 46674
rect 74946 46622 74958 46674
rect 75010 46622 75022 46674
rect 46734 46610 46786 46622
rect 3614 46562 3666 46574
rect 2034 46510 2046 46562
rect 2098 46510 2110 46562
rect 3614 46498 3666 46510
rect 48190 46562 48242 46574
rect 48190 46498 48242 46510
rect 74510 46562 74562 46574
rect 75954 46510 75966 46562
rect 76018 46510 76030 46562
rect 74510 46498 74562 46510
rect 1344 46282 78624 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 78624 46282
rect 1344 46196 78624 46230
rect 46062 45890 46114 45902
rect 3042 45838 3054 45890
rect 3106 45838 3118 45890
rect 46946 45838 46958 45890
rect 47010 45838 47022 45890
rect 74946 45838 74958 45890
rect 75010 45838 75022 45890
rect 46062 45826 46114 45838
rect 47182 45778 47234 45790
rect 1922 45726 1934 45778
rect 1986 45726 1998 45778
rect 76066 45726 76078 45778
rect 76130 45726 76142 45778
rect 47182 45714 47234 45726
rect 3502 45666 3554 45678
rect 3502 45602 3554 45614
rect 45726 45666 45778 45678
rect 45726 45602 45778 45614
rect 47742 45666 47794 45678
rect 47742 45602 47794 45614
rect 48190 45666 48242 45678
rect 48190 45602 48242 45614
rect 74398 45666 74450 45678
rect 74398 45602 74450 45614
rect 1344 45498 78624 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 78624 45498
rect 1344 45412 78624 45446
rect 44382 45330 44434 45342
rect 44382 45266 44434 45278
rect 45614 45330 45666 45342
rect 45614 45266 45666 45278
rect 46174 45218 46226 45230
rect 46174 45154 46226 45166
rect 47406 45218 47458 45230
rect 47406 45154 47458 45166
rect 43934 45106 43986 45118
rect 3042 45054 3054 45106
rect 3106 45054 3118 45106
rect 43934 45042 43986 45054
rect 44718 45106 44770 45118
rect 46510 45106 46562 45118
rect 45378 45054 45390 45106
rect 45442 45054 45454 45106
rect 47170 45054 47182 45106
rect 47234 45054 47246 45106
rect 74946 45054 74958 45106
rect 75010 45054 75022 45106
rect 44718 45042 44770 45054
rect 46510 45042 46562 45054
rect 3614 44994 3666 45006
rect 2034 44942 2046 44994
rect 2098 44942 2110 44994
rect 3614 44930 3666 44942
rect 47854 44994 47906 45006
rect 47854 44930 47906 44942
rect 48302 44994 48354 45006
rect 48302 44930 48354 44942
rect 74510 44994 74562 45006
rect 75954 44942 75966 44994
rect 76018 44942 76030 44994
rect 74510 44930 74562 44942
rect 1344 44714 78624 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 78624 44714
rect 1344 44628 78624 44662
rect 3042 44270 3054 44322
rect 3106 44270 3118 44322
rect 74946 44270 74958 44322
rect 75010 44270 75022 44322
rect 43710 44210 43762 44222
rect 1922 44158 1934 44210
rect 1986 44158 1998 44210
rect 43710 44146 43762 44158
rect 44046 44210 44098 44222
rect 44046 44146 44098 44158
rect 44606 44210 44658 44222
rect 44606 44146 44658 44158
rect 45502 44210 45554 44222
rect 45502 44146 45554 44158
rect 46398 44210 46450 44222
rect 76066 44158 76078 44210
rect 76130 44158 76142 44210
rect 46398 44146 46450 44158
rect 3502 44098 3554 44110
rect 3502 44034 3554 44046
rect 45838 44098 45890 44110
rect 45838 44034 45890 44046
rect 46734 44098 46786 44110
rect 46734 44034 46786 44046
rect 74398 44098 74450 44110
rect 74398 44034 74450 44046
rect 1344 43930 78624 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 78624 43930
rect 1344 43844 78624 43878
rect 43038 43762 43090 43774
rect 43038 43698 43090 43710
rect 44494 43762 44546 43774
rect 44494 43698 44546 43710
rect 42590 43538 42642 43550
rect 3042 43486 3054 43538
rect 3106 43486 3118 43538
rect 42590 43474 42642 43486
rect 43374 43538 43426 43550
rect 44258 43486 44270 43538
rect 44322 43486 44334 43538
rect 74946 43486 74958 43538
rect 75010 43486 75022 43538
rect 43374 43474 43426 43486
rect 3614 43426 3666 43438
rect 1922 43374 1934 43426
rect 1986 43374 1998 43426
rect 3614 43362 3666 43374
rect 44942 43426 44994 43438
rect 44942 43362 44994 43374
rect 74510 43426 74562 43438
rect 76066 43374 76078 43426
rect 76130 43374 76142 43426
rect 74510 43362 74562 43374
rect 1344 43146 78624 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 78624 43146
rect 1344 43060 78624 43094
rect 3042 42702 3054 42754
rect 3106 42702 3118 42754
rect 43474 42702 43486 42754
rect 43538 42702 43550 42754
rect 74946 42702 74958 42754
rect 75010 42702 75022 42754
rect 3502 42642 3554 42654
rect 1922 42590 1934 42642
rect 1986 42590 1998 42642
rect 3502 42578 3554 42590
rect 42366 42642 42418 42654
rect 42366 42578 42418 42590
rect 42702 42642 42754 42654
rect 42702 42578 42754 42590
rect 44270 42642 44322 42654
rect 76066 42590 76078 42642
rect 76130 42590 76142 42642
rect 44270 42578 44322 42590
rect 41918 42530 41970 42542
rect 41918 42466 41970 42478
rect 43710 42530 43762 42542
rect 43710 42466 43762 42478
rect 74398 42530 74450 42542
rect 74398 42466 74450 42478
rect 1344 42362 78624 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 78624 42362
rect 1344 42276 78624 42310
rect 41806 42194 41858 42206
rect 41806 42130 41858 42142
rect 43150 42082 43202 42094
rect 43150 42018 43202 42030
rect 42142 41970 42194 41982
rect 3042 41918 3054 41970
rect 3106 41918 3118 41970
rect 42914 41918 42926 41970
rect 42978 41918 42990 41970
rect 74946 41918 74958 41970
rect 75010 41918 75022 41970
rect 42142 41906 42194 41918
rect 3614 41858 3666 41870
rect 1922 41806 1934 41858
rect 1986 41806 1998 41858
rect 3614 41794 3666 41806
rect 43598 41858 43650 41870
rect 43598 41794 43650 41806
rect 74510 41858 74562 41870
rect 76066 41806 76078 41858
rect 76130 41806 76142 41858
rect 74510 41794 74562 41806
rect 1344 41578 78624 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 78624 41578
rect 1344 41492 78624 41526
rect 3042 41134 3054 41186
rect 3106 41134 3118 41186
rect 74946 41134 74958 41186
rect 75010 41134 75022 41186
rect 41022 41074 41074 41086
rect 1922 41022 1934 41074
rect 1986 41022 1998 41074
rect 41022 41010 41074 41022
rect 41358 41074 41410 41086
rect 41358 41010 41410 41022
rect 42142 41074 42194 41086
rect 76066 41022 76078 41074
rect 76130 41022 76142 41074
rect 42142 41010 42194 41022
rect 3502 40962 3554 40974
rect 3502 40898 3554 40910
rect 40126 40962 40178 40974
rect 40126 40898 40178 40910
rect 40574 40962 40626 40974
rect 40574 40898 40626 40910
rect 42478 40962 42530 40974
rect 42478 40898 42530 40910
rect 42926 40962 42978 40974
rect 42926 40898 42978 40910
rect 74398 40962 74450 40974
rect 74398 40898 74450 40910
rect 1344 40794 78624 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 78624 40794
rect 1344 40708 78624 40742
rect 40350 40626 40402 40638
rect 40350 40562 40402 40574
rect 42366 40626 42418 40638
rect 42366 40562 42418 40574
rect 39454 40514 39506 40526
rect 39454 40450 39506 40462
rect 41918 40514 41970 40526
rect 41918 40450 41970 40462
rect 3614 40402 3666 40414
rect 3042 40350 3054 40402
rect 3106 40350 3118 40402
rect 3614 40338 3666 40350
rect 39790 40402 39842 40414
rect 39790 40338 39842 40350
rect 40686 40402 40738 40414
rect 40686 40338 40738 40350
rect 41582 40402 41634 40414
rect 41582 40338 41634 40350
rect 42814 40402 42866 40414
rect 42814 40338 42866 40350
rect 74510 40402 74562 40414
rect 76078 40402 76130 40414
rect 74946 40350 74958 40402
rect 75010 40350 75022 40402
rect 74510 40338 74562 40350
rect 76078 40338 76130 40350
rect 39006 40290 39058 40302
rect 1922 40238 1934 40290
rect 1986 40238 1998 40290
rect 39006 40226 39058 40238
rect 1344 40010 78624 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 78624 40010
rect 1344 39924 78624 39958
rect 1934 39618 1986 39630
rect 76078 39618 76130 39630
rect 3042 39566 3054 39618
rect 3106 39566 3118 39618
rect 74946 39566 74958 39618
rect 75010 39566 75022 39618
rect 1934 39554 1986 39566
rect 76078 39554 76130 39566
rect 3614 39506 3666 39518
rect 3614 39442 3666 39454
rect 38894 39506 38946 39518
rect 38894 39442 38946 39454
rect 39230 39506 39282 39518
rect 39230 39442 39282 39454
rect 39790 39506 39842 39518
rect 39790 39442 39842 39454
rect 40686 39506 40738 39518
rect 40686 39442 40738 39454
rect 41022 39506 41074 39518
rect 41022 39442 41074 39454
rect 38446 39394 38498 39406
rect 38446 39330 38498 39342
rect 40126 39394 40178 39406
rect 40126 39330 40178 39342
rect 41470 39394 41522 39406
rect 41470 39330 41522 39342
rect 74510 39394 74562 39406
rect 74510 39330 74562 39342
rect 1344 39226 78624 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 78624 39226
rect 1344 39140 78624 39174
rect 38334 38946 38386 38958
rect 1922 38894 1934 38946
rect 1986 38894 1998 38946
rect 38334 38882 38386 38894
rect 39678 38946 39730 38958
rect 39678 38882 39730 38894
rect 74510 38946 74562 38958
rect 76066 38894 76078 38946
rect 76130 38894 76142 38946
rect 74510 38882 74562 38894
rect 3614 38834 3666 38846
rect 3042 38782 3054 38834
rect 3106 38782 3118 38834
rect 3614 38770 3666 38782
rect 38670 38834 38722 38846
rect 39442 38782 39454 38834
rect 39506 38782 39518 38834
rect 74946 38782 74958 38834
rect 75010 38782 75022 38834
rect 38670 38770 38722 38782
rect 37886 38722 37938 38734
rect 37886 38658 37938 38670
rect 40350 38722 40402 38734
rect 40350 38658 40402 38670
rect 1344 38442 78624 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 78624 38442
rect 1344 38356 78624 38390
rect 1922 38110 1934 38162
rect 1986 38110 1998 38162
rect 76066 38110 76078 38162
rect 76130 38110 76142 38162
rect 3042 37998 3054 38050
rect 3106 37998 3118 38050
rect 38882 37998 38894 38050
rect 38946 37998 38958 38050
rect 74946 37998 74958 38050
rect 75010 37998 75022 38050
rect 37998 37938 38050 37950
rect 37998 37874 38050 37886
rect 40014 37938 40066 37950
rect 40014 37874 40066 37886
rect 3614 37826 3666 37838
rect 3614 37762 3666 37774
rect 37662 37826 37714 37838
rect 37662 37762 37714 37774
rect 39118 37826 39170 37838
rect 39118 37762 39170 37774
rect 39566 37826 39618 37838
rect 39566 37762 39618 37774
rect 74510 37826 74562 37838
rect 74510 37762 74562 37774
rect 1344 37658 78624 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 78624 37658
rect 1344 37572 78624 37606
rect 36990 37378 37042 37390
rect 1922 37326 1934 37378
rect 1986 37326 1998 37378
rect 36990 37314 37042 37326
rect 38446 37378 38498 37390
rect 38446 37314 38498 37326
rect 74510 37378 74562 37390
rect 76066 37326 76078 37378
rect 76130 37326 76142 37378
rect 74510 37314 74562 37326
rect 36542 37266 36594 37278
rect 3042 37214 3054 37266
rect 3106 37214 3118 37266
rect 36542 37202 36594 37214
rect 37326 37266 37378 37278
rect 37326 37202 37378 37214
rect 38110 37266 38162 37278
rect 38110 37202 38162 37214
rect 39342 37266 39394 37278
rect 74946 37214 74958 37266
rect 75010 37214 75022 37266
rect 39342 37202 39394 37214
rect 3614 37154 3666 37166
rect 3614 37090 3666 37102
rect 38894 37154 38946 37166
rect 38894 37090 38946 37102
rect 39106 36990 39118 37042
rect 39170 37039 39182 37042
rect 39442 37039 39454 37042
rect 39170 36993 39454 37039
rect 39170 36990 39182 36993
rect 39442 36990 39454 36993
rect 39506 36990 39518 37042
rect 1344 36874 78624 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 78624 36874
rect 1344 36788 78624 36822
rect 1922 36542 1934 36594
rect 1986 36542 1998 36594
rect 76066 36542 76078 36594
rect 76130 36542 76142 36594
rect 3042 36430 3054 36482
rect 3106 36430 3118 36482
rect 36530 36430 36542 36482
rect 36594 36430 36606 36482
rect 74946 36430 74958 36482
rect 75010 36430 75022 36482
rect 35870 36370 35922 36382
rect 35870 36306 35922 36318
rect 37550 36370 37602 36382
rect 37550 36306 37602 36318
rect 3614 36258 3666 36270
rect 3614 36194 3666 36206
rect 35422 36258 35474 36270
rect 35422 36194 35474 36206
rect 36318 36258 36370 36270
rect 36318 36194 36370 36206
rect 37886 36258 37938 36270
rect 37886 36194 37938 36206
rect 74510 36258 74562 36270
rect 74510 36194 74562 36206
rect 1344 36090 78624 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 78624 36090
rect 1344 36004 78624 36038
rect 34750 35810 34802 35822
rect 1922 35758 1934 35810
rect 1986 35758 1998 35810
rect 34750 35746 34802 35758
rect 35646 35810 35698 35822
rect 35646 35746 35698 35758
rect 36990 35810 37042 35822
rect 36990 35746 37042 35758
rect 74510 35810 74562 35822
rect 76066 35758 76078 35810
rect 76130 35758 76142 35810
rect 74510 35746 74562 35758
rect 35982 35698 36034 35710
rect 3042 35646 3054 35698
rect 3106 35646 3118 35698
rect 4834 35646 4846 35698
rect 4898 35646 4910 35698
rect 34962 35646 34974 35698
rect 35026 35646 35038 35698
rect 35982 35634 36034 35646
rect 36654 35698 36706 35710
rect 36654 35634 36706 35646
rect 37886 35698 37938 35710
rect 37886 35634 37938 35646
rect 38334 35698 38386 35710
rect 74946 35646 74958 35698
rect 75010 35646 75022 35698
rect 76738 35646 76750 35698
rect 76802 35646 76814 35698
rect 38334 35634 38386 35646
rect 5406 35586 5458 35598
rect 3714 35534 3726 35586
rect 3778 35534 3790 35586
rect 5406 35522 5458 35534
rect 37438 35586 37490 35598
rect 77858 35534 77870 35586
rect 77922 35534 77934 35586
rect 37438 35522 37490 35534
rect 1344 35306 78624 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 78624 35306
rect 1344 35220 78624 35254
rect 3614 35026 3666 35038
rect 1922 34974 1934 35026
rect 1986 34974 1998 35026
rect 3614 34962 3666 34974
rect 37438 35026 37490 35038
rect 76066 34974 76078 35026
rect 76130 34974 76142 35026
rect 37438 34962 37490 34974
rect 36094 34914 36146 34926
rect 3042 34862 3054 34914
rect 3106 34862 3118 34914
rect 35298 34862 35310 34914
rect 35362 34862 35374 34914
rect 74946 34862 74958 34914
rect 75010 34862 75022 34914
rect 36094 34850 36146 34862
rect 33854 34802 33906 34814
rect 33854 34738 33906 34750
rect 34302 34802 34354 34814
rect 34302 34738 34354 34750
rect 34638 34802 34690 34814
rect 34638 34738 34690 34750
rect 36430 34802 36482 34814
rect 36430 34738 36482 34750
rect 74510 34802 74562 34814
rect 74510 34738 74562 34750
rect 4062 34690 4114 34702
rect 4062 34626 4114 34638
rect 35534 34690 35586 34702
rect 35534 34626 35586 34638
rect 77198 34690 77250 34702
rect 77198 34626 77250 34638
rect 1344 34522 78624 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 78624 34522
rect 1344 34436 78624 34470
rect 33742 34242 33794 34254
rect 1922 34190 1934 34242
rect 1986 34190 1998 34242
rect 33742 34178 33794 34190
rect 35086 34242 35138 34254
rect 35086 34178 35138 34190
rect 74510 34242 74562 34254
rect 76066 34190 76078 34242
rect 76130 34190 76142 34242
rect 74510 34178 74562 34190
rect 34078 34130 34130 34142
rect 36206 34130 36258 34142
rect 3042 34078 3054 34130
rect 3106 34078 3118 34130
rect 34850 34078 34862 34130
rect 34914 34078 34926 34130
rect 74946 34078 74958 34130
rect 75010 34078 75022 34130
rect 34078 34066 34130 34078
rect 36206 34066 36258 34078
rect 3614 34018 3666 34030
rect 3614 33954 3666 33966
rect 35758 34018 35810 34030
rect 35758 33954 35810 33966
rect 1344 33738 78624 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 78624 33738
rect 1344 33652 78624 33686
rect 34862 33458 34914 33470
rect 1922 33406 1934 33458
rect 1986 33406 1998 33458
rect 76066 33406 76078 33458
rect 76130 33406 76142 33458
rect 34862 33394 34914 33406
rect 34078 33346 34130 33358
rect 3042 33294 3054 33346
rect 3106 33294 3118 33346
rect 33170 33294 33182 33346
rect 33234 33294 33246 33346
rect 74946 33294 74958 33346
rect 75010 33294 75022 33346
rect 34078 33282 34130 33294
rect 3614 33234 3666 33246
rect 3614 33170 3666 33182
rect 32958 33234 33010 33246
rect 32958 33170 33010 33182
rect 32510 33122 32562 33134
rect 32510 33058 32562 33070
rect 34414 33122 34466 33134
rect 34414 33058 34466 33070
rect 74510 33122 74562 33134
rect 74510 33058 74562 33070
rect 1344 32954 78624 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 78624 32954
rect 1344 32868 78624 32902
rect 34414 32786 34466 32798
rect 34414 32722 34466 32734
rect 32286 32674 32338 32686
rect 1922 32622 1934 32674
rect 1986 32622 1998 32674
rect 32286 32610 32338 32622
rect 33966 32674 34018 32686
rect 33966 32610 34018 32622
rect 74510 32674 74562 32686
rect 76066 32622 76078 32674
rect 76130 32622 76142 32674
rect 74510 32610 74562 32622
rect 33630 32562 33682 32574
rect 3042 32510 3054 32562
rect 3106 32510 3118 32562
rect 32498 32510 32510 32562
rect 32562 32510 32574 32562
rect 74946 32510 74958 32562
rect 75010 32510 75022 32562
rect 33630 32498 33682 32510
rect 3614 32450 3666 32462
rect 3614 32386 3666 32398
rect 31838 32450 31890 32462
rect 31838 32386 31890 32398
rect 1344 32170 78624 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 78624 32170
rect 1344 32084 78624 32118
rect 33518 31890 33570 31902
rect 1922 31838 1934 31890
rect 1986 31838 1998 31890
rect 76066 31838 76078 31890
rect 76130 31838 76142 31890
rect 33518 31826 33570 31838
rect 31950 31778 32002 31790
rect 33966 31778 34018 31790
rect 3042 31726 3054 31778
rect 3106 31726 3118 31778
rect 32834 31726 32846 31778
rect 32898 31726 32910 31778
rect 74946 31726 74958 31778
rect 75010 31726 75022 31778
rect 31950 31714 32002 31726
rect 33966 31714 34018 31726
rect 3614 31554 3666 31566
rect 3614 31490 3666 31502
rect 30718 31554 30770 31566
rect 30718 31490 30770 31502
rect 31166 31554 31218 31566
rect 31166 31490 31218 31502
rect 31614 31554 31666 31566
rect 31614 31490 31666 31502
rect 33070 31554 33122 31566
rect 33070 31490 33122 31502
rect 74510 31554 74562 31566
rect 74510 31490 74562 31502
rect 1344 31386 78624 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 78624 31386
rect 1344 31300 78624 31334
rect 30046 31106 30098 31118
rect 1922 31054 1934 31106
rect 1986 31054 1998 31106
rect 30046 31042 30098 31054
rect 30942 31106 30994 31118
rect 30942 31042 30994 31054
rect 32286 31106 32338 31118
rect 32286 31042 32338 31054
rect 74510 31106 74562 31118
rect 76066 31054 76078 31106
rect 76130 31054 76142 31106
rect 74510 31042 74562 31054
rect 30382 30994 30434 31006
rect 3042 30942 3054 30994
rect 3106 30942 3118 30994
rect 4834 30942 4846 30994
rect 4898 30942 4910 30994
rect 30382 30930 30434 30942
rect 31278 30994 31330 31006
rect 32734 30994 32786 31006
rect 32050 30942 32062 30994
rect 32114 30942 32126 30994
rect 74946 30942 74958 30994
rect 75010 30942 75022 30994
rect 76738 30942 76750 30994
rect 76802 30942 76814 30994
rect 31278 30930 31330 30942
rect 32734 30930 32786 30942
rect 5406 30882 5458 30894
rect 3714 30830 3726 30882
rect 3778 30830 3790 30882
rect 5406 30818 5458 30830
rect 29374 30882 29426 30894
rect 77858 30830 77870 30882
rect 77922 30830 77934 30882
rect 29374 30818 29426 30830
rect 1344 30602 78624 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 78624 30602
rect 1344 30516 78624 30550
rect 32174 30322 32226 30334
rect 1922 30270 1934 30322
rect 1986 30270 1998 30322
rect 32174 30258 32226 30270
rect 3614 30210 3666 30222
rect 76078 30210 76130 30222
rect 3042 30158 3054 30210
rect 3106 30158 3118 30210
rect 74946 30158 74958 30210
rect 75010 30158 75022 30210
rect 3614 30146 3666 30158
rect 76078 30146 76130 30158
rect 29598 30098 29650 30110
rect 29598 30034 29650 30046
rect 29934 30098 29986 30110
rect 29934 30034 29986 30046
rect 30494 30098 30546 30110
rect 30494 30034 30546 30046
rect 31390 30098 31442 30110
rect 31390 30034 31442 30046
rect 31726 30098 31778 30110
rect 31726 30034 31778 30046
rect 74510 30098 74562 30110
rect 74510 30034 74562 30046
rect 4062 29986 4114 29998
rect 4062 29922 4114 29934
rect 28814 29986 28866 29998
rect 28814 29922 28866 29934
rect 30830 29986 30882 29998
rect 30830 29922 30882 29934
rect 77198 29986 77250 29998
rect 77198 29922 77250 29934
rect 1344 29818 78624 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 78624 29818
rect 1344 29732 78624 29766
rect 28926 29538 28978 29550
rect 1922 29486 1934 29538
rect 1986 29486 1998 29538
rect 28926 29474 28978 29486
rect 30382 29538 30434 29550
rect 30382 29474 30434 29486
rect 74510 29538 74562 29550
rect 76066 29486 76078 29538
rect 76130 29486 76142 29538
rect 74510 29474 74562 29486
rect 28478 29426 28530 29438
rect 3042 29374 3054 29426
rect 3106 29374 3118 29426
rect 28478 29362 28530 29374
rect 29262 29426 29314 29438
rect 29262 29362 29314 29374
rect 30046 29426 30098 29438
rect 30046 29362 30098 29374
rect 31054 29426 31106 29438
rect 74946 29374 74958 29426
rect 75010 29374 75022 29426
rect 31054 29362 31106 29374
rect 3614 29314 3666 29326
rect 3614 29250 3666 29262
rect 31502 29314 31554 29326
rect 31502 29250 31554 29262
rect 1344 29034 78624 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 78624 29034
rect 1344 28948 78624 28982
rect 1922 28702 1934 28754
rect 1986 28702 1998 28754
rect 76066 28702 76078 28754
rect 76130 28702 76142 28754
rect 3614 28642 3666 28654
rect 3042 28590 3054 28642
rect 3106 28590 3118 28642
rect 3614 28578 3666 28590
rect 27806 28642 27858 28654
rect 27806 28578 27858 28590
rect 74510 28642 74562 28654
rect 74946 28590 74958 28642
rect 75010 28590 75022 28642
rect 74510 28578 74562 28590
rect 28254 28530 28306 28542
rect 28254 28466 28306 28478
rect 28590 28530 28642 28542
rect 28590 28466 28642 28478
rect 29598 28530 29650 28542
rect 29598 28466 29650 28478
rect 29934 28418 29986 28430
rect 29934 28354 29986 28366
rect 1344 28250 78624 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 78624 28250
rect 1344 28164 78624 28198
rect 29374 28082 29426 28094
rect 29374 28018 29426 28030
rect 27582 27970 27634 27982
rect 1922 27918 1934 27970
rect 1986 27918 1998 27970
rect 27582 27906 27634 27918
rect 28926 27970 28978 27982
rect 28926 27906 28978 27918
rect 74510 27970 74562 27982
rect 76066 27918 76078 27970
rect 76130 27918 76142 27970
rect 74510 27906 74562 27918
rect 28590 27858 28642 27870
rect 3042 27806 3054 27858
rect 3106 27806 3118 27858
rect 27794 27806 27806 27858
rect 27858 27806 27870 27858
rect 28590 27794 28642 27806
rect 29822 27858 29874 27870
rect 74946 27806 74958 27858
rect 75010 27806 75022 27858
rect 29822 27794 29874 27806
rect 3614 27746 3666 27758
rect 3614 27682 3666 27694
rect 27134 27746 27186 27758
rect 27134 27682 27186 27694
rect 1344 27466 78624 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 78624 27466
rect 1344 27380 78624 27414
rect 1922 27134 1934 27186
rect 1986 27134 1998 27186
rect 76066 27134 76078 27186
rect 76130 27134 76142 27186
rect 3614 27074 3666 27086
rect 3042 27022 3054 27074
rect 3106 27022 3118 27074
rect 74946 27022 74958 27074
rect 75010 27022 75022 27074
rect 3614 27010 3666 27022
rect 26462 26962 26514 26974
rect 26462 26898 26514 26910
rect 27246 26962 27298 26974
rect 27246 26898 27298 26910
rect 27918 26962 27970 26974
rect 27918 26898 27970 26910
rect 28814 26962 28866 26974
rect 28814 26898 28866 26910
rect 74510 26962 74562 26974
rect 74510 26898 74562 26910
rect 26910 26850 26962 26862
rect 26910 26786 26962 26798
rect 28254 26850 28306 26862
rect 28254 26786 28306 26798
rect 1344 26682 78624 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 78624 26682
rect 1344 26596 78624 26630
rect 26238 26402 26290 26414
rect 1922 26350 1934 26402
rect 1986 26350 1998 26402
rect 26238 26338 26290 26350
rect 27694 26402 27746 26414
rect 27694 26338 27746 26350
rect 74510 26402 74562 26414
rect 76066 26350 76078 26402
rect 76130 26350 76142 26402
rect 74510 26338 74562 26350
rect 25790 26290 25842 26302
rect 2930 26238 2942 26290
rect 2994 26238 3006 26290
rect 4834 26238 4846 26290
rect 4898 26238 4910 26290
rect 25790 26226 25842 26238
rect 26574 26290 26626 26302
rect 26574 26226 26626 26238
rect 27358 26290 27410 26302
rect 74946 26238 74958 26290
rect 75010 26238 75022 26290
rect 76962 26238 76974 26290
rect 77026 26238 77038 26290
rect 27358 26226 27410 26238
rect 5406 26178 5458 26190
rect 3714 26126 3726 26178
rect 3778 26126 3790 26178
rect 5406 26114 5458 26126
rect 25006 26178 25058 26190
rect 77858 26126 77870 26178
rect 77922 26126 77934 26178
rect 25006 26114 25058 26126
rect 1344 25898 78624 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 78624 25898
rect 1344 25812 78624 25846
rect 1922 25566 1934 25618
rect 1986 25566 1998 25618
rect 76066 25566 76078 25618
rect 76130 25566 76142 25618
rect 25566 25506 25618 25518
rect 27582 25506 27634 25518
rect 3042 25454 3054 25506
rect 3106 25454 3118 25506
rect 26450 25454 26462 25506
rect 26514 25454 26526 25506
rect 74946 25454 74958 25506
rect 75010 25454 75022 25506
rect 25566 25442 25618 25454
rect 27582 25442 27634 25454
rect 4062 25394 4114 25406
rect 4062 25330 4114 25342
rect 24334 25394 24386 25406
rect 24334 25330 24386 25342
rect 24670 25394 24722 25406
rect 24670 25330 24722 25342
rect 25230 25394 25282 25406
rect 25230 25330 25282 25342
rect 27134 25394 27186 25406
rect 27134 25330 27186 25342
rect 3614 25282 3666 25294
rect 3614 25218 3666 25230
rect 26686 25282 26738 25294
rect 26686 25218 26738 25230
rect 74510 25282 74562 25294
rect 74510 25218 74562 25230
rect 77198 25282 77250 25294
rect 77198 25218 77250 25230
rect 1344 25114 78624 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 78624 25114
rect 1344 25028 78624 25062
rect 23662 24834 23714 24846
rect 1922 24782 1934 24834
rect 1986 24782 1998 24834
rect 23662 24770 23714 24782
rect 24894 24834 24946 24846
rect 24894 24770 24946 24782
rect 26126 24834 26178 24846
rect 76066 24782 76078 24834
rect 76130 24782 76142 24834
rect 26126 24770 26178 24782
rect 22766 24722 22818 24734
rect 3042 24670 3054 24722
rect 3106 24670 3118 24722
rect 22766 24658 22818 24670
rect 23102 24722 23154 24734
rect 23102 24658 23154 24670
rect 23998 24722 24050 24734
rect 23998 24658 24050 24670
rect 24558 24722 24610 24734
rect 74510 24722 74562 24734
rect 25890 24670 25902 24722
rect 25954 24670 25966 24722
rect 74946 24670 74958 24722
rect 75010 24670 75022 24722
rect 24558 24658 24610 24670
rect 74510 24658 74562 24670
rect 3614 24610 3666 24622
rect 3614 24546 3666 24558
rect 26574 24610 26626 24622
rect 26574 24546 26626 24558
rect 1344 24330 78624 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 78624 24330
rect 1344 24244 78624 24278
rect 1922 23998 1934 24050
rect 1986 23998 1998 24050
rect 76066 23998 76078 24050
rect 76130 23998 76142 24050
rect 3042 23886 3054 23938
rect 3106 23886 3118 23938
rect 74946 23886 74958 23938
rect 75010 23886 75022 23938
rect 23998 23826 24050 23838
rect 23998 23762 24050 23774
rect 25342 23826 25394 23838
rect 25342 23762 25394 23774
rect 3614 23714 3666 23726
rect 3614 23650 3666 23662
rect 23102 23714 23154 23726
rect 23102 23650 23154 23662
rect 23662 23714 23714 23726
rect 23662 23650 23714 23662
rect 24894 23714 24946 23726
rect 24894 23650 24946 23662
rect 25678 23714 25730 23726
rect 25678 23650 25730 23662
rect 26126 23714 26178 23726
rect 26126 23650 26178 23662
rect 74510 23714 74562 23726
rect 74510 23650 74562 23662
rect 1344 23546 78624 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 78624 23546
rect 1344 23460 78624 23494
rect 22430 23266 22482 23278
rect 1922 23214 1934 23266
rect 1986 23214 1998 23266
rect 22430 23202 22482 23214
rect 23886 23266 23938 23278
rect 23886 23202 23938 23214
rect 74510 23266 74562 23278
rect 76066 23214 76078 23266
rect 76130 23214 76142 23266
rect 74510 23202 74562 23214
rect 22766 23154 22818 23166
rect 3042 23102 3054 23154
rect 3106 23102 3118 23154
rect 23650 23102 23662 23154
rect 23714 23102 23726 23154
rect 74946 23102 74958 23154
rect 75010 23102 75022 23154
rect 22766 23090 22818 23102
rect 3614 23042 3666 23054
rect 3614 22978 3666 22990
rect 24334 23042 24386 23054
rect 24334 22978 24386 22990
rect 1344 22762 78624 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 78624 22762
rect 1344 22676 78624 22710
rect 1922 22430 1934 22482
rect 1986 22430 1998 22482
rect 76066 22430 76078 22482
rect 76130 22430 76142 22482
rect 3042 22318 3054 22370
rect 3106 22318 3118 22370
rect 23090 22318 23102 22370
rect 23154 22318 23166 22370
rect 74946 22318 74958 22370
rect 75010 22318 75022 22370
rect 22430 22258 22482 22270
rect 22430 22194 22482 22206
rect 3614 22146 3666 22158
rect 3614 22082 3666 22094
rect 22094 22146 22146 22158
rect 22094 22082 22146 22094
rect 23326 22146 23378 22158
rect 23326 22082 23378 22094
rect 23774 22146 23826 22158
rect 23774 22082 23826 22094
rect 24334 22146 24386 22158
rect 24334 22082 24386 22094
rect 74510 22146 74562 22158
rect 74510 22082 74562 22094
rect 1344 21978 78624 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 78624 21978
rect 1344 21892 78624 21926
rect 22654 21810 22706 21822
rect 22654 21746 22706 21758
rect 21758 21698 21810 21710
rect 1922 21646 1934 21698
rect 1986 21646 1998 21698
rect 21758 21634 21810 21646
rect 23998 21698 24050 21710
rect 23998 21634 24050 21646
rect 74510 21698 74562 21710
rect 76066 21646 76078 21698
rect 76130 21646 76142 21698
rect 74510 21634 74562 21646
rect 22094 21586 22146 21598
rect 2930 21534 2942 21586
rect 2994 21534 3006 21586
rect 4834 21534 4846 21586
rect 4898 21534 4910 21586
rect 22094 21522 22146 21534
rect 23102 21586 23154 21598
rect 23102 21522 23154 21534
rect 23662 21586 23714 21598
rect 23662 21522 23714 21534
rect 24446 21586 24498 21598
rect 74946 21534 74958 21586
rect 75010 21534 75022 21586
rect 76962 21534 76974 21586
rect 77026 21534 77038 21586
rect 24446 21522 24498 21534
rect 5406 21474 5458 21486
rect 3714 21422 3726 21474
rect 3778 21422 3790 21474
rect 77858 21422 77870 21474
rect 77922 21422 77934 21474
rect 5406 21410 5458 21422
rect 1344 21194 78624 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 78624 21194
rect 1344 21108 78624 21142
rect 3614 20914 3666 20926
rect 1922 20862 1934 20914
rect 1986 20862 1998 20914
rect 76066 20862 76078 20914
rect 76130 20862 76142 20914
rect 3614 20850 3666 20862
rect 22766 20802 22818 20814
rect 3042 20750 3054 20802
rect 3106 20750 3118 20802
rect 21858 20750 21870 20802
rect 21922 20750 21934 20802
rect 22766 20738 22818 20750
rect 23214 20802 23266 20814
rect 74946 20750 74958 20802
rect 75010 20750 75022 20802
rect 23214 20738 23266 20750
rect 4062 20690 4114 20702
rect 4062 20626 4114 20638
rect 21646 20690 21698 20702
rect 21646 20626 21698 20638
rect 20974 20578 21026 20590
rect 20974 20514 21026 20526
rect 23550 20578 23602 20590
rect 23550 20514 23602 20526
rect 74510 20578 74562 20590
rect 74510 20514 74562 20526
rect 77198 20578 77250 20590
rect 77198 20514 77250 20526
rect 1344 20410 78624 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 78624 20410
rect 1344 20324 78624 20358
rect 19966 20242 20018 20254
rect 19966 20178 20018 20190
rect 21198 20242 21250 20254
rect 21198 20178 21250 20190
rect 1922 20078 1934 20130
rect 1986 20078 1998 20130
rect 76066 20078 76078 20130
rect 76130 20078 76142 20130
rect 19518 20018 19570 20030
rect 3042 19966 3054 20018
rect 3106 19966 3118 20018
rect 19518 19954 19570 19966
rect 20302 20018 20354 20030
rect 20302 19954 20354 19966
rect 20862 20018 20914 20030
rect 20862 19954 20914 19966
rect 21646 20018 21698 20030
rect 74946 19966 74958 20018
rect 75010 19966 75022 20018
rect 21646 19954 21698 19966
rect 3614 19906 3666 19918
rect 3614 19842 3666 19854
rect 74510 19906 74562 19918
rect 74510 19842 74562 19854
rect 1344 19626 78624 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 78624 19626
rect 1344 19540 78624 19574
rect 1922 19294 1934 19346
rect 1986 19294 1998 19346
rect 76066 19294 76078 19346
rect 76130 19294 76142 19346
rect 3042 19182 3054 19234
rect 3106 19182 3118 19234
rect 18946 19182 18958 19234
rect 19010 19182 19022 19234
rect 74946 19182 74958 19234
rect 75010 19182 75022 19234
rect 19630 19122 19682 19134
rect 19630 19058 19682 19070
rect 19966 19122 20018 19134
rect 19966 19058 20018 19070
rect 20526 19122 20578 19134
rect 20526 19058 20578 19070
rect 21646 19122 21698 19134
rect 21646 19058 21698 19070
rect 21982 19122 22034 19134
rect 21982 19058 22034 19070
rect 74510 19122 74562 19134
rect 74510 19058 74562 19070
rect 3614 19010 3666 19022
rect 3614 18946 3666 18958
rect 18286 19010 18338 19022
rect 18286 18946 18338 18958
rect 18734 19010 18786 19022
rect 18734 18946 18786 18958
rect 20862 19010 20914 19022
rect 20862 18946 20914 18958
rect 22430 19010 22482 19022
rect 22430 18946 22482 18958
rect 1344 18842 78624 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 78624 18842
rect 1344 18756 78624 18790
rect 21534 18674 21586 18686
rect 56242 18622 56254 18674
rect 56306 18622 56318 18674
rect 21534 18610 21586 18622
rect 18622 18562 18674 18574
rect 1922 18510 1934 18562
rect 1986 18510 1998 18562
rect 18622 18498 18674 18510
rect 21086 18562 21138 18574
rect 21086 18498 21138 18510
rect 55582 18562 55634 18574
rect 55582 18498 55634 18510
rect 18958 18450 19010 18462
rect 3042 18398 3054 18450
rect 3106 18398 3118 18450
rect 18958 18386 19010 18398
rect 20750 18450 20802 18462
rect 20750 18386 20802 18398
rect 55806 18450 55858 18462
rect 55806 18386 55858 18398
rect 56030 18450 56082 18462
rect 56030 18386 56082 18398
rect 56254 18450 56306 18462
rect 56254 18386 56306 18398
rect 74510 18450 74562 18462
rect 76078 18450 76130 18462
rect 74946 18398 74958 18450
rect 75010 18398 75022 18450
rect 74510 18386 74562 18398
rect 76078 18386 76130 18398
rect 3614 18338 3666 18350
rect 3614 18274 3666 18286
rect 18174 18338 18226 18350
rect 18174 18274 18226 18286
rect 19742 18338 19794 18350
rect 19742 18274 19794 18286
rect 20190 18338 20242 18350
rect 20190 18274 20242 18286
rect 54574 18338 54626 18350
rect 54574 18274 54626 18286
rect 55022 18338 55074 18350
rect 55022 18274 55074 18286
rect 1344 18058 78624 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 78624 18058
rect 1344 17972 78624 18006
rect 20750 17890 20802 17902
rect 20750 17826 20802 17838
rect 56254 17890 56306 17902
rect 56254 17826 56306 17838
rect 55694 17778 55746 17790
rect 1922 17726 1934 17778
rect 1986 17726 1998 17778
rect 26226 17726 26238 17778
rect 26290 17726 26302 17778
rect 76066 17726 76078 17778
rect 76130 17726 76142 17778
rect 55694 17714 55746 17726
rect 17166 17666 17218 17678
rect 3042 17614 3054 17666
rect 3106 17614 3118 17666
rect 17166 17602 17218 17614
rect 20190 17666 20242 17678
rect 20190 17602 20242 17614
rect 20302 17666 20354 17678
rect 20302 17602 20354 17614
rect 20526 17666 20578 17678
rect 20526 17602 20578 17614
rect 54126 17666 54178 17678
rect 54126 17602 54178 17614
rect 55022 17666 55074 17678
rect 55022 17602 55074 17614
rect 55582 17666 55634 17678
rect 55582 17602 55634 17614
rect 56142 17666 56194 17678
rect 74946 17614 74958 17666
rect 75010 17614 75022 17666
rect 56142 17602 56194 17614
rect 17950 17554 18002 17566
rect 17950 17490 18002 17502
rect 18510 17554 18562 17566
rect 18510 17490 18562 17502
rect 18846 17554 18898 17566
rect 18846 17490 18898 17502
rect 20862 17554 20914 17566
rect 20862 17490 20914 17502
rect 25902 17554 25954 17566
rect 25902 17490 25954 17502
rect 74510 17554 74562 17566
rect 74510 17490 74562 17502
rect 3614 17442 3666 17454
rect 3614 17378 3666 17390
rect 16382 17442 16434 17454
rect 16382 17378 16434 17390
rect 17614 17442 17666 17454
rect 17614 17378 17666 17390
rect 19294 17442 19346 17454
rect 19294 17378 19346 17390
rect 21534 17442 21586 17454
rect 21534 17378 21586 17390
rect 21982 17442 22034 17454
rect 21982 17378 22034 17390
rect 24110 17442 24162 17454
rect 24110 17378 24162 17390
rect 25006 17442 25058 17454
rect 25006 17378 25058 17390
rect 25342 17442 25394 17454
rect 25342 17378 25394 17390
rect 26126 17442 26178 17454
rect 26126 17378 26178 17390
rect 53678 17442 53730 17454
rect 53678 17378 53730 17390
rect 55134 17442 55186 17454
rect 55134 17378 55186 17390
rect 55358 17442 55410 17454
rect 55358 17378 55410 17390
rect 56702 17442 56754 17454
rect 56702 17378 56754 17390
rect 1344 17274 78624 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 78624 17274
rect 1344 17188 78624 17222
rect 19966 17106 20018 17118
rect 19966 17042 20018 17054
rect 21086 17106 21138 17118
rect 21086 17042 21138 17054
rect 24446 17106 24498 17118
rect 24446 17042 24498 17054
rect 15710 16994 15762 17006
rect 1922 16942 1934 16994
rect 1986 16942 1998 16994
rect 15710 16930 15762 16942
rect 16606 16994 16658 17006
rect 16606 16930 16658 16942
rect 18510 16994 18562 17006
rect 18510 16930 18562 16942
rect 19518 16994 19570 17006
rect 19518 16930 19570 16942
rect 26014 16994 26066 17006
rect 26014 16930 26066 16942
rect 74510 16994 74562 17006
rect 76066 16942 76078 16994
rect 76130 16942 76142 16994
rect 74510 16930 74562 16942
rect 5406 16882 5458 16894
rect 3042 16830 3054 16882
rect 3106 16830 3118 16882
rect 4834 16830 4846 16882
rect 4898 16830 4910 16882
rect 5406 16818 5458 16830
rect 16046 16882 16098 16894
rect 16046 16818 16098 16830
rect 16942 16882 16994 16894
rect 16942 16818 16994 16830
rect 18174 16882 18226 16894
rect 18174 16818 18226 16830
rect 19182 16882 19234 16894
rect 19182 16818 19234 16830
rect 20414 16882 20466 16894
rect 24894 16882 24946 16894
rect 23650 16830 23662 16882
rect 23714 16830 23726 16882
rect 20414 16818 20466 16830
rect 24894 16818 24946 16830
rect 25678 16882 25730 16894
rect 25678 16818 25730 16830
rect 25902 16882 25954 16894
rect 26686 16882 26738 16894
rect 26226 16830 26238 16882
rect 26290 16830 26302 16882
rect 25902 16818 25954 16830
rect 26686 16818 26738 16830
rect 54574 16882 54626 16894
rect 77870 16882 77922 16894
rect 74946 16830 74958 16882
rect 75010 16830 75022 16882
rect 76738 16830 76750 16882
rect 76802 16830 76814 16882
rect 54574 16818 54626 16830
rect 77870 16818 77922 16830
rect 17614 16770 17666 16782
rect 3714 16718 3726 16770
rect 3778 16718 3790 16770
rect 17614 16706 17666 16718
rect 22318 16770 22370 16782
rect 22318 16706 22370 16718
rect 22990 16770 23042 16782
rect 22990 16706 23042 16718
rect 23214 16770 23266 16782
rect 23214 16706 23266 16718
rect 22878 16658 22930 16670
rect 22878 16594 22930 16606
rect 23438 16658 23490 16670
rect 23438 16594 23490 16606
rect 1344 16490 78624 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 78624 16490
rect 1344 16404 78624 16438
rect 18734 16322 18786 16334
rect 18734 16258 18786 16270
rect 22878 16322 22930 16334
rect 23202 16270 23214 16322
rect 23266 16270 23278 16322
rect 22878 16258 22930 16270
rect 3614 16210 3666 16222
rect 1922 16158 1934 16210
rect 1986 16158 1998 16210
rect 76066 16158 76078 16210
rect 76130 16158 76142 16210
rect 3614 16146 3666 16158
rect 18286 16098 18338 16110
rect 3042 16046 3054 16098
rect 3106 16046 3118 16098
rect 18050 16046 18062 16098
rect 18114 16046 18126 16098
rect 18286 16034 18338 16046
rect 18510 16098 18562 16110
rect 18510 16034 18562 16046
rect 18846 16098 18898 16110
rect 18846 16034 18898 16046
rect 22654 16098 22706 16110
rect 22654 16034 22706 16046
rect 74510 16098 74562 16110
rect 74946 16046 74958 16098
rect 75010 16046 75022 16098
rect 74510 16034 74562 16046
rect 15822 15986 15874 15998
rect 15822 15922 15874 15934
rect 16158 15986 16210 15998
rect 16158 15922 16210 15934
rect 19406 15986 19458 15998
rect 19406 15922 19458 15934
rect 20190 15986 20242 15998
rect 20190 15922 20242 15934
rect 4062 15874 4114 15886
rect 4062 15810 4114 15822
rect 16718 15874 16770 15886
rect 16718 15810 16770 15822
rect 17166 15874 17218 15886
rect 17166 15810 17218 15822
rect 19742 15874 19794 15886
rect 19742 15810 19794 15822
rect 23886 15874 23938 15886
rect 23886 15810 23938 15822
rect 24334 15874 24386 15886
rect 24334 15810 24386 15822
rect 77198 15874 77250 15886
rect 77198 15810 77250 15822
rect 1344 15706 78624 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 78624 15706
rect 1344 15620 78624 15654
rect 14702 15426 14754 15438
rect 1922 15374 1934 15426
rect 1986 15374 1998 15426
rect 14702 15362 14754 15374
rect 18174 15426 18226 15438
rect 18174 15362 18226 15374
rect 56366 15426 56418 15438
rect 56366 15362 56418 15374
rect 74510 15426 74562 15438
rect 76066 15374 76078 15426
rect 76130 15374 76142 15426
rect 74510 15362 74562 15374
rect 15038 15314 15090 15326
rect 3042 15262 3054 15314
rect 3106 15262 3118 15314
rect 15038 15250 15090 15262
rect 16382 15314 16434 15326
rect 16382 15250 16434 15262
rect 56030 15314 56082 15326
rect 74946 15262 74958 15314
rect 75010 15262 75022 15314
rect 56030 15250 56082 15262
rect 3614 15202 3666 15214
rect 3614 15138 3666 15150
rect 15486 15202 15538 15214
rect 15486 15138 15538 15150
rect 17726 15202 17778 15214
rect 17726 15138 17778 15150
rect 19070 15202 19122 15214
rect 19070 15138 19122 15150
rect 55470 15202 55522 15214
rect 55470 15138 55522 15150
rect 1344 14922 78624 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 78624 14922
rect 1344 14836 78624 14870
rect 55358 14754 55410 14766
rect 55358 14690 55410 14702
rect 54126 14642 54178 14654
rect 1922 14590 1934 14642
rect 1986 14590 1998 14642
rect 76066 14590 76078 14642
rect 76130 14590 76142 14642
rect 54126 14578 54178 14590
rect 55134 14530 55186 14542
rect 56814 14530 56866 14542
rect 3042 14478 3054 14530
rect 3106 14478 3118 14530
rect 54898 14478 54910 14530
rect 54962 14478 54974 14530
rect 56130 14478 56142 14530
rect 56194 14478 56206 14530
rect 74946 14478 74958 14530
rect 75010 14478 75022 14530
rect 55134 14466 55186 14478
rect 56814 14466 56866 14478
rect 14366 14418 14418 14430
rect 14366 14354 14418 14366
rect 3614 14306 3666 14318
rect 3614 14242 3666 14254
rect 14030 14306 14082 14318
rect 14030 14242 14082 14254
rect 14814 14306 14866 14318
rect 14814 14242 14866 14254
rect 53678 14306 53730 14318
rect 53678 14242 53730 14254
rect 55022 14306 55074 14318
rect 55022 14242 55074 14254
rect 56366 14306 56418 14318
rect 56366 14242 56418 14254
rect 74510 14306 74562 14318
rect 74510 14242 74562 14254
rect 1344 14138 78624 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 78624 14138
rect 1344 14052 78624 14086
rect 12462 13858 12514 13870
rect 1922 13806 1934 13858
rect 1986 13806 1998 13858
rect 12462 13794 12514 13806
rect 13358 13858 13410 13870
rect 13358 13794 13410 13806
rect 55694 13858 55746 13870
rect 55694 13794 55746 13806
rect 57822 13858 57874 13870
rect 57822 13794 57874 13806
rect 74510 13858 74562 13870
rect 76066 13806 76078 13858
rect 76130 13806 76142 13858
rect 74510 13794 74562 13806
rect 12798 13746 12850 13758
rect 3042 13694 3054 13746
rect 3106 13694 3118 13746
rect 12798 13682 12850 13694
rect 13694 13746 13746 13758
rect 13694 13682 13746 13694
rect 14142 13746 14194 13758
rect 14142 13682 14194 13694
rect 54574 13746 54626 13758
rect 54574 13682 54626 13694
rect 55358 13746 55410 13758
rect 55358 13682 55410 13694
rect 57486 13746 57538 13758
rect 74946 13694 74958 13746
rect 75010 13694 75022 13746
rect 57486 13682 57538 13694
rect 3614 13634 3666 13646
rect 3614 13570 3666 13582
rect 12014 13634 12066 13646
rect 12014 13570 12066 13582
rect 56702 13634 56754 13646
rect 56702 13570 56754 13582
rect 1344 13354 78624 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 78624 13354
rect 1344 13268 78624 13302
rect 55022 13074 55074 13086
rect 1922 13022 1934 13074
rect 1986 13022 1998 13074
rect 55022 13010 55074 13022
rect 74510 13074 74562 13086
rect 76066 13022 76078 13074
rect 76130 13022 76142 13074
rect 74510 13010 74562 13022
rect 3042 12910 3054 12962
rect 3106 12910 3118 12962
rect 74946 12910 74958 12962
rect 75010 12910 75022 12962
rect 3614 12738 3666 12750
rect 3614 12674 3666 12686
rect 12014 12738 12066 12750
rect 12014 12674 12066 12686
rect 12910 12738 12962 12750
rect 12910 12674 12962 12686
rect 1344 12570 78624 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 78624 12570
rect 1344 12484 78624 12518
rect 11342 12290 11394 12302
rect 1922 12238 1934 12290
rect 1986 12238 1998 12290
rect 11342 12226 11394 12238
rect 12238 12290 12290 12302
rect 12238 12226 12290 12238
rect 13470 12290 13522 12302
rect 13470 12226 13522 12238
rect 74510 12290 74562 12302
rect 76066 12238 76078 12290
rect 76130 12238 76142 12290
rect 74510 12226 74562 12238
rect 11678 12178 11730 12190
rect 3042 12126 3054 12178
rect 3106 12126 3118 12178
rect 4834 12126 4846 12178
rect 4898 12126 4910 12178
rect 11678 12114 11730 12126
rect 12574 12178 12626 12190
rect 13234 12126 13246 12178
rect 13298 12126 13310 12178
rect 74946 12126 74958 12178
rect 75010 12126 75022 12178
rect 76738 12126 76750 12178
rect 76802 12126 76814 12178
rect 12574 12114 12626 12126
rect 13918 12066 13970 12078
rect 3714 12014 3726 12066
rect 3778 12014 3790 12066
rect 77858 12014 77870 12066
rect 77922 12014 77934 12066
rect 13918 12002 13970 12014
rect 1344 11786 78624 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 78624 11786
rect 1344 11700 78624 11734
rect 3614 11506 3666 11518
rect 1922 11454 1934 11506
rect 1986 11454 1998 11506
rect 3614 11442 3666 11454
rect 4062 11506 4114 11518
rect 76066 11454 76078 11506
rect 76130 11454 76142 11506
rect 4062 11442 4114 11454
rect 13582 11394 13634 11406
rect 3042 11342 3054 11394
rect 3106 11342 3118 11394
rect 12562 11342 12574 11394
rect 12626 11342 12638 11394
rect 74946 11342 74958 11394
rect 75010 11342 75022 11394
rect 13582 11330 13634 11342
rect 10670 11282 10722 11294
rect 10670 11218 10722 11230
rect 11006 11282 11058 11294
rect 11006 11218 11058 11230
rect 11566 11282 11618 11294
rect 11566 11218 11618 11230
rect 12798 11282 12850 11294
rect 12798 11218 12850 11230
rect 74510 11282 74562 11294
rect 74510 11218 74562 11230
rect 11902 11170 11954 11182
rect 11902 11106 11954 11118
rect 77198 11170 77250 11182
rect 77198 11106 77250 11118
rect 1344 11002 78624 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 78624 11002
rect 1344 10916 78624 10950
rect 10110 10722 10162 10734
rect 1922 10670 1934 10722
rect 1986 10670 1998 10722
rect 10110 10658 10162 10670
rect 11454 10722 11506 10734
rect 11454 10658 11506 10670
rect 74510 10722 74562 10734
rect 76066 10670 76078 10722
rect 76130 10670 76142 10722
rect 74510 10658 74562 10670
rect 10446 10610 10498 10622
rect 3042 10558 3054 10610
rect 3106 10558 3118 10610
rect 10446 10546 10498 10558
rect 11118 10610 11170 10622
rect 74946 10558 74958 10610
rect 75010 10558 75022 10610
rect 11118 10546 11170 10558
rect 1344 10218 78624 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 78624 10218
rect 1344 10132 78624 10166
rect 1922 9886 1934 9938
rect 1986 9886 1998 9938
rect 76066 9886 76078 9938
rect 76130 9886 76142 9938
rect 3042 9774 3054 9826
rect 3106 9774 3118 9826
rect 9650 9774 9662 9826
rect 9714 9774 9726 9826
rect 74946 9774 74958 9826
rect 75010 9774 75022 9826
rect 9438 9714 9490 9726
rect 9438 9650 9490 9662
rect 10558 9714 10610 9726
rect 10558 9650 10610 9662
rect 10894 9602 10946 9614
rect 10894 9538 10946 9550
rect 74510 9602 74562 9614
rect 74510 9538 74562 9550
rect 1344 9434 78624 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 78624 9434
rect 1344 9348 78624 9382
rect 8654 9154 8706 9166
rect 1922 9102 1934 9154
rect 1986 9102 1998 9154
rect 8654 9090 8706 9102
rect 10222 9154 10274 9166
rect 10222 9090 10274 9102
rect 74510 9154 74562 9166
rect 76066 9102 76078 9154
rect 76130 9102 76142 9154
rect 74510 9090 74562 9102
rect 8990 9042 9042 9054
rect 3042 8990 3054 9042
rect 3106 8990 3118 9042
rect 8990 8978 9042 8990
rect 9886 9042 9938 9054
rect 74946 8990 74958 9042
rect 75010 8990 75022 9042
rect 9886 8978 9938 8990
rect 1344 8650 78624 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 78624 8650
rect 1344 8564 78624 8598
rect 1922 8318 1934 8370
rect 1986 8318 1998 8370
rect 76066 8318 76078 8370
rect 76130 8318 76142 8370
rect 3042 8206 3054 8258
rect 3106 8206 3118 8258
rect 74946 8206 74958 8258
rect 75010 8206 75022 8258
rect 8094 8146 8146 8158
rect 8094 8082 8146 8094
rect 8430 8146 8482 8158
rect 8430 8082 8482 8094
rect 9102 8146 9154 8158
rect 9102 8082 9154 8094
rect 9438 8034 9490 8046
rect 9438 7970 9490 7982
rect 74510 8034 74562 8046
rect 74510 7970 74562 7982
rect 1344 7866 78624 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 78624 7866
rect 1344 7780 78624 7814
rect 6526 7586 6578 7598
rect 1922 7534 1934 7586
rect 1986 7534 1998 7586
rect 6526 7522 6578 7534
rect 7422 7586 7474 7598
rect 7422 7522 7474 7534
rect 8766 7586 8818 7598
rect 8766 7522 8818 7534
rect 74510 7586 74562 7598
rect 76066 7534 76078 7586
rect 76130 7534 76142 7586
rect 74510 7522 74562 7534
rect 6862 7474 6914 7486
rect 8430 7474 8482 7486
rect 3042 7422 3054 7474
rect 3106 7422 3118 7474
rect 4834 7422 4846 7474
rect 4898 7422 4910 7474
rect 7634 7422 7646 7474
rect 7698 7422 7710 7474
rect 74946 7422 74958 7474
rect 75010 7422 75022 7474
rect 76738 7422 76750 7474
rect 76802 7422 76814 7474
rect 6862 7410 6914 7422
rect 8430 7410 8482 7422
rect 18062 7362 18114 7374
rect 3714 7310 3726 7362
rect 3778 7310 3790 7362
rect 77858 7310 77870 7362
rect 77922 7310 77934 7362
rect 18062 7298 18114 7310
rect 1344 7082 78624 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 78624 7082
rect 1344 6996 78624 7030
rect 1922 6750 1934 6802
rect 1986 6750 1998 6802
rect 16258 6750 16270 6802
rect 16322 6750 16334 6802
rect 19506 6750 19518 6802
rect 19570 6750 19582 6802
rect 23650 6750 23662 6802
rect 23714 6750 23726 6802
rect 27010 6750 27022 6802
rect 27074 6750 27086 6802
rect 70018 6750 70030 6802
rect 70082 6750 70094 6802
rect 6974 6690 7026 6702
rect 3042 6638 3054 6690
rect 3106 6638 3118 6690
rect 6290 6638 6302 6690
rect 6354 6638 6366 6690
rect 6974 6626 7026 6638
rect 7870 6690 7922 6702
rect 7870 6626 7922 6638
rect 68686 6690 68738 6702
rect 76078 6690 76130 6702
rect 69346 6638 69358 6690
rect 69410 6638 69422 6690
rect 74946 6638 74958 6690
rect 75010 6638 75022 6690
rect 68686 6626 68738 6638
rect 76078 6626 76130 6638
rect 6078 6578 6130 6590
rect 6078 6514 6130 6526
rect 7310 6578 7362 6590
rect 66782 6578 66834 6590
rect 17266 6526 17278 6578
rect 17330 6526 17342 6578
rect 18498 6526 18510 6578
rect 18562 6526 18574 6578
rect 22418 6526 22430 6578
rect 22482 6526 22494 6578
rect 28018 6526 28030 6578
rect 28082 6526 28094 6578
rect 7310 6514 7362 6526
rect 66782 6514 66834 6526
rect 77198 6578 77250 6590
rect 77198 6514 77250 6526
rect 8206 6466 8258 6478
rect 8206 6402 8258 6414
rect 8654 6466 8706 6478
rect 8654 6402 8706 6414
rect 20638 6466 20690 6478
rect 20638 6402 20690 6414
rect 21870 6466 21922 6478
rect 21870 6402 21922 6414
rect 26574 6466 26626 6478
rect 26574 6402 26626 6414
rect 31054 6466 31106 6478
rect 31054 6402 31106 6414
rect 74510 6466 74562 6478
rect 74510 6402 74562 6414
rect 1344 6298 78624 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 78624 6298
rect 1344 6212 78624 6246
rect 53006 6130 53058 6142
rect 53006 6066 53058 6078
rect 54238 6130 54290 6142
rect 54238 6066 54290 6078
rect 55022 6130 55074 6142
rect 55022 6066 55074 6078
rect 55358 6130 55410 6142
rect 55358 6066 55410 6078
rect 57374 6130 57426 6142
rect 57374 6066 57426 6078
rect 58158 6130 58210 6142
rect 58158 6066 58210 6078
rect 58718 6130 58770 6142
rect 58718 6066 58770 6078
rect 59166 6130 59218 6142
rect 59166 6066 59218 6078
rect 59614 6130 59666 6142
rect 59614 6066 59666 6078
rect 60286 6130 60338 6142
rect 60286 6066 60338 6078
rect 61182 6130 61234 6142
rect 61182 6066 61234 6078
rect 61518 6130 61570 6142
rect 61518 6066 61570 6078
rect 62078 6130 62130 6142
rect 62078 6066 62130 6078
rect 64206 6130 64258 6142
rect 64206 6066 64258 6078
rect 65326 6130 65378 6142
rect 65326 6066 65378 6078
rect 65774 6130 65826 6142
rect 65774 6066 65826 6078
rect 66334 6130 66386 6142
rect 66334 6066 66386 6078
rect 66782 6130 66834 6142
rect 66782 6066 66834 6078
rect 4622 6018 4674 6030
rect 1922 5966 1934 6018
rect 1986 5966 1998 6018
rect 6850 5966 6862 6018
rect 6914 5966 6926 6018
rect 8642 5966 8654 6018
rect 8706 5966 8718 6018
rect 15922 5966 15934 6018
rect 15986 5966 15998 6018
rect 20290 5966 20302 6018
rect 20354 5966 20366 6018
rect 21970 5966 21982 6018
rect 22034 5966 22046 6018
rect 23090 5966 23102 6018
rect 23154 5966 23166 6018
rect 28690 5966 28702 6018
rect 28754 5966 28766 6018
rect 30370 5966 30382 6018
rect 30434 5966 30446 6018
rect 32386 5966 32398 6018
rect 32450 5966 32462 6018
rect 35186 5966 35198 6018
rect 35250 5966 35262 6018
rect 47282 5966 47294 6018
rect 47346 5966 47358 6018
rect 76066 5966 76078 6018
rect 76130 5966 76142 6018
rect 4622 5954 4674 5966
rect 4958 5906 5010 5918
rect 3042 5854 3054 5906
rect 3106 5854 3118 5906
rect 4958 5842 5010 5854
rect 18398 5906 18450 5918
rect 51214 5906 51266 5918
rect 70814 5906 70866 5918
rect 50530 5854 50542 5906
rect 50594 5854 50606 5906
rect 67330 5854 67342 5906
rect 67394 5854 67406 5906
rect 70130 5854 70142 5906
rect 70194 5854 70206 5906
rect 74946 5854 74958 5906
rect 75010 5854 75022 5906
rect 76738 5854 76750 5906
rect 76802 5854 76814 5906
rect 18398 5842 18450 5854
rect 51214 5842 51266 5854
rect 70814 5842 70866 5854
rect 4174 5794 4226 5806
rect 11118 5794 11170 5806
rect 5506 5742 5518 5794
rect 5570 5742 5582 5794
rect 7746 5742 7758 5794
rect 7810 5742 7822 5794
rect 4174 5730 4226 5742
rect 11118 5730 11170 5742
rect 11902 5794 11954 5806
rect 11902 5730 11954 5742
rect 13470 5794 13522 5806
rect 13470 5730 13522 5742
rect 13918 5794 13970 5806
rect 13918 5730 13970 5742
rect 14478 5794 14530 5806
rect 17950 5794 18002 5806
rect 33518 5794 33570 5806
rect 16706 5742 16718 5794
rect 16770 5742 16782 5794
rect 18946 5742 18958 5794
rect 19010 5742 19022 5794
rect 20962 5742 20974 5794
rect 21026 5742 21038 5794
rect 24210 5742 24222 5794
rect 24274 5742 24286 5794
rect 27346 5742 27358 5794
rect 27410 5742 27422 5794
rect 29362 5742 29374 5794
rect 29426 5742 29438 5794
rect 31602 5742 31614 5794
rect 31666 5742 31678 5794
rect 14478 5730 14530 5742
rect 17950 5730 18002 5742
rect 33518 5730 33570 5742
rect 34638 5794 34690 5806
rect 38782 5794 38834 5806
rect 36306 5742 36318 5794
rect 36370 5742 36382 5794
rect 34638 5730 34690 5742
rect 38782 5730 38834 5742
rect 40238 5794 40290 5806
rect 40238 5730 40290 5742
rect 42254 5794 42306 5806
rect 42254 5730 42306 5742
rect 45390 5794 45442 5806
rect 45390 5730 45442 5742
rect 46734 5794 46786 5806
rect 51662 5794 51714 5806
rect 48402 5742 48414 5794
rect 48466 5742 48478 5794
rect 49634 5742 49646 5794
rect 49698 5742 49710 5794
rect 46734 5730 46786 5742
rect 51662 5730 51714 5742
rect 55806 5794 55858 5806
rect 55806 5730 55858 5742
rect 56366 5794 56418 5806
rect 73390 5794 73442 5806
rect 68002 5742 68014 5794
rect 68066 5742 68078 5794
rect 69234 5742 69246 5794
rect 69298 5742 69310 5794
rect 56366 5730 56418 5742
rect 73390 5730 73442 5742
rect 73838 5794 73890 5806
rect 73838 5730 73890 5742
rect 74510 5794 74562 5806
rect 77858 5742 77870 5794
rect 77922 5742 77934 5794
rect 74510 5730 74562 5742
rect 73490 5630 73502 5682
rect 73554 5679 73566 5682
rect 73826 5679 73838 5682
rect 73554 5633 73838 5679
rect 73554 5630 73566 5633
rect 73826 5630 73838 5633
rect 73890 5630 73902 5682
rect 1344 5514 78624 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 78624 5514
rect 1344 5428 78624 5462
rect 21982 5234 22034 5246
rect 29486 5234 29538 5246
rect 1922 5182 1934 5234
rect 1986 5182 1998 5234
rect 7634 5182 7646 5234
rect 7698 5182 7710 5234
rect 9650 5182 9662 5234
rect 9714 5182 9726 5234
rect 11554 5182 11566 5234
rect 11618 5182 11630 5234
rect 16706 5182 16718 5234
rect 16770 5182 16782 5234
rect 18610 5182 18622 5234
rect 18674 5182 18686 5234
rect 20850 5182 20862 5234
rect 20914 5182 20926 5234
rect 24658 5182 24670 5234
rect 24722 5182 24734 5234
rect 25442 5182 25454 5234
rect 25506 5182 25518 5234
rect 27570 5182 27582 5234
rect 27634 5182 27646 5234
rect 31266 5182 31278 5234
rect 31330 5182 31342 5234
rect 34514 5182 34526 5234
rect 34578 5182 34590 5234
rect 35298 5182 35310 5234
rect 35362 5182 35374 5234
rect 39666 5182 39678 5234
rect 39730 5182 39742 5234
rect 40450 5182 40462 5234
rect 40514 5182 40526 5234
rect 43698 5182 43710 5234
rect 43762 5182 43774 5234
rect 46946 5182 46958 5234
rect 47010 5182 47022 5234
rect 48738 5182 48750 5234
rect 48802 5182 48814 5234
rect 51986 5182 51998 5234
rect 52050 5182 52062 5234
rect 55906 5182 55918 5234
rect 55970 5182 55982 5234
rect 59938 5182 59950 5234
rect 60002 5182 60014 5234
rect 62066 5182 62078 5234
rect 62130 5182 62142 5234
rect 67778 5182 67790 5234
rect 67842 5182 67854 5234
rect 70130 5182 70142 5234
rect 70194 5182 70206 5234
rect 73266 5182 73278 5234
rect 73330 5182 73342 5234
rect 74050 5182 74062 5234
rect 74114 5182 74126 5234
rect 21982 5170 22034 5182
rect 29486 5170 29538 5182
rect 14478 5122 14530 5134
rect 3042 5070 3054 5122
rect 3106 5070 3118 5122
rect 14478 5058 14530 5070
rect 21646 5122 21698 5134
rect 21646 5058 21698 5070
rect 22766 5122 22818 5134
rect 22766 5058 22818 5070
rect 30830 5122 30882 5134
rect 30830 5058 30882 5070
rect 37438 5122 37490 5134
rect 37438 5058 37490 5070
rect 44830 5122 44882 5134
rect 44830 5058 44882 5070
rect 49646 5122 49698 5134
rect 57374 5122 57426 5134
rect 71598 5122 71650 5134
rect 50754 5070 50766 5122
rect 50818 5070 50830 5122
rect 51314 5070 51326 5122
rect 51378 5070 51390 5122
rect 54450 5070 54462 5122
rect 54514 5070 54526 5122
rect 55234 5070 55246 5122
rect 55298 5070 55310 5122
rect 58482 5070 58494 5122
rect 58546 5070 58558 5122
rect 59266 5070 59278 5122
rect 59330 5070 59342 5122
rect 61394 5070 61406 5122
rect 61458 5070 61470 5122
rect 64530 5070 64542 5122
rect 64594 5070 64606 5122
rect 66322 5070 66334 5122
rect 66386 5070 66398 5122
rect 67106 5070 67118 5122
rect 67170 5070 67182 5122
rect 69346 5070 69358 5122
rect 69410 5070 69422 5122
rect 49646 5058 49698 5070
rect 57374 5058 57426 5070
rect 71598 5058 71650 5070
rect 76526 5122 76578 5134
rect 76526 5058 76578 5070
rect 4622 5010 4674 5022
rect 4622 4946 4674 4958
rect 6414 5010 6466 5022
rect 13694 5010 13746 5022
rect 8418 4958 8430 5010
rect 8482 4958 8494 5010
rect 10434 4958 10446 5010
rect 10498 4958 10510 5010
rect 12450 4958 12462 5010
rect 12514 4958 12526 5010
rect 6414 4946 6466 4958
rect 13694 4946 13746 4958
rect 14030 5010 14082 5022
rect 29934 5010 29986 5022
rect 15810 4958 15822 5010
rect 15874 4958 15886 5010
rect 17826 4958 17838 5010
rect 17890 4958 17902 5010
rect 19506 4958 19518 5010
rect 19570 4958 19582 5010
rect 23762 4958 23774 5010
rect 23826 4958 23838 5010
rect 26674 4958 26686 5010
rect 26738 4958 26750 5010
rect 28354 4958 28366 5010
rect 28418 4958 28430 5010
rect 32274 4958 32286 5010
rect 32338 4958 32350 5010
rect 33730 4958 33742 5010
rect 33794 4958 33806 5010
rect 36306 4958 36318 5010
rect 36370 4958 36382 5010
rect 38658 4958 38670 5010
rect 38722 4958 38734 5010
rect 41458 4958 41470 5010
rect 41522 4958 41534 5010
rect 42578 4958 42590 5010
rect 42642 4958 42654 5010
rect 45602 4958 45614 5010
rect 45666 4958 45678 5010
rect 47618 4958 47630 5010
rect 47682 4958 47694 5010
rect 53554 4958 53566 5010
rect 53618 4958 53630 5010
rect 63410 4958 63422 5010
rect 63474 4958 63486 5010
rect 65426 4958 65438 5010
rect 65490 4958 65502 5010
rect 72258 4958 72270 5010
rect 72322 4958 72334 5010
rect 75058 4958 75070 5010
rect 75122 4958 75134 5010
rect 14030 4946 14082 4958
rect 29934 4946 29986 4958
rect 4958 4898 5010 4910
rect 4958 4834 5010 4846
rect 6750 4898 6802 4910
rect 6750 4834 6802 4846
rect 37998 4898 38050 4910
rect 37998 4834 38050 4846
rect 1344 4730 78624 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 78624 4730
rect 1344 4644 78624 4678
rect 4622 4562 4674 4574
rect 4622 4498 4674 4510
rect 16830 4562 16882 4574
rect 16830 4498 16882 4510
rect 69470 4562 69522 4574
rect 69470 4498 69522 4510
rect 6738 4398 6750 4450
rect 6802 4398 6814 4450
rect 7970 4398 7982 4450
rect 8034 4398 8046 4450
rect 11218 4398 11230 4450
rect 11282 4398 11294 4450
rect 12674 4398 12686 4450
rect 12738 4398 12750 4450
rect 14354 4398 14366 4450
rect 14418 4398 14430 4450
rect 19842 4398 19854 4450
rect 19906 4398 19918 4450
rect 21858 4398 21870 4450
rect 21922 4398 21934 4450
rect 24770 4398 24782 4450
rect 24834 4398 24846 4450
rect 28690 4398 28702 4450
rect 28754 4398 28766 4450
rect 29810 4398 29822 4450
rect 29874 4398 29886 4450
rect 32722 4398 32734 4450
rect 32786 4398 32798 4450
rect 35522 4398 35534 4450
rect 35586 4398 35598 4450
rect 38098 4398 38110 4450
rect 38162 4398 38174 4450
rect 40114 4398 40126 4450
rect 40178 4398 40190 4450
rect 41682 4398 41694 4450
rect 41746 4398 41758 4450
rect 44594 4398 44606 4450
rect 44658 4398 44670 4450
rect 45714 4398 45726 4450
rect 45778 4398 45790 4450
rect 50530 4398 50542 4450
rect 50594 4398 50606 4450
rect 70802 4398 70814 4450
rect 70866 4398 70878 4450
rect 74386 4398 74398 4450
rect 74450 4398 74462 4450
rect 76402 4398 76414 4450
rect 76466 4398 76478 4450
rect 9662 4338 9714 4350
rect 4834 4286 4846 4338
rect 4898 4286 4910 4338
rect 9662 4274 9714 4286
rect 26014 4338 26066 4350
rect 26014 4274 26066 4286
rect 33518 4338 33570 4350
rect 64542 4338 64594 4350
rect 68910 4338 68962 4350
rect 51538 4286 51550 4338
rect 51602 4286 51614 4338
rect 53330 4286 53342 4338
rect 53394 4286 53406 4338
rect 56130 4286 56142 4338
rect 56194 4286 56206 4338
rect 57474 4286 57486 4338
rect 57538 4286 57550 4338
rect 59378 4286 59390 4338
rect 59442 4286 59454 4338
rect 61058 4286 61070 4338
rect 61122 4286 61134 4338
rect 63858 4286 63870 4338
rect 63922 4286 63934 4338
rect 65650 4286 65662 4338
rect 65714 4286 65726 4338
rect 68226 4286 68238 4338
rect 68290 4286 68302 4338
rect 33518 4274 33570 4286
rect 64542 4274 64594 4286
rect 68910 4274 68962 4286
rect 17614 4226 17666 4238
rect 5730 4174 5742 4226
rect 5794 4174 5806 4226
rect 8978 4174 8990 4226
rect 9042 4174 9054 4226
rect 10434 4174 10446 4226
rect 10498 4174 10510 4226
rect 13570 4174 13582 4226
rect 13634 4174 13646 4226
rect 17614 4162 17666 4174
rect 18062 4226 18114 4238
rect 18062 4162 18114 4174
rect 18846 4226 18898 4238
rect 25566 4226 25618 4238
rect 20738 4174 20750 4226
rect 20802 4174 20814 4226
rect 22642 4174 22654 4226
rect 22706 4174 22718 4226
rect 23426 4174 23438 4226
rect 23490 4174 23502 4226
rect 18846 4162 18898 4174
rect 25566 4162 25618 4174
rect 26798 4226 26850 4238
rect 33966 4226 34018 4238
rect 27458 4174 27470 4226
rect 27522 4174 27534 4226
rect 30594 4174 30606 4226
rect 30658 4174 30670 4226
rect 31490 4174 31502 4226
rect 31554 4174 31566 4226
rect 26798 4162 26850 4174
rect 33966 4162 34018 4174
rect 34526 4226 34578 4238
rect 47518 4226 47570 4238
rect 36530 4174 36542 4226
rect 36594 4174 36606 4226
rect 37314 4174 37326 4226
rect 37378 4174 37390 4226
rect 39106 4174 39118 4226
rect 39170 4174 39182 4226
rect 42802 4174 42814 4226
rect 42866 4174 42878 4226
rect 43586 4174 43598 4226
rect 43650 4174 43662 4226
rect 46834 4174 46846 4226
rect 46898 4174 46910 4226
rect 34526 4162 34578 4174
rect 47518 4162 47570 4174
rect 48750 4226 48802 4238
rect 70254 4226 70306 4238
rect 72718 4226 72770 4238
rect 49522 4174 49534 4226
rect 49586 4174 49598 4226
rect 52210 4174 52222 4226
rect 52274 4174 52286 4226
rect 54002 4174 54014 4226
rect 54066 4174 54078 4226
rect 55458 4174 55470 4226
rect 55522 4174 55534 4226
rect 58146 4174 58158 4226
rect 58210 4174 58222 4226
rect 59938 4174 59950 4226
rect 60002 4174 60014 4226
rect 61730 4174 61742 4226
rect 61794 4174 61806 4226
rect 62962 4174 62974 4226
rect 63026 4174 63038 4226
rect 66098 4174 66110 4226
rect 66162 4174 66174 4226
rect 67330 4174 67342 4226
rect 67394 4174 67406 4226
rect 71922 4174 71934 4226
rect 71986 4174 71998 4226
rect 73378 4174 73390 4226
rect 73442 4174 73454 4226
rect 75394 4174 75406 4226
rect 75458 4174 75470 4226
rect 48750 4162 48802 4174
rect 70254 4162 70306 4174
rect 72718 4162 72770 4174
rect 1344 3946 78624 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 78624 3946
rect 1344 3860 78624 3894
rect 16830 3778 16882 3790
rect 16830 3714 16882 3726
rect 9550 3666 9602 3678
rect 19742 3666 19794 3678
rect 4946 3614 4958 3666
rect 5010 3614 5022 3666
rect 8866 3614 8878 3666
rect 8930 3614 8942 3666
rect 12562 3614 12574 3666
rect 12626 3614 12638 3666
rect 9550 3602 9602 3614
rect 19742 3602 19794 3614
rect 21310 3666 21362 3678
rect 37886 3666 37938 3678
rect 44270 3666 44322 3678
rect 46846 3666 46898 3678
rect 51102 3666 51154 3678
rect 24322 3614 24334 3666
rect 24386 3614 24398 3666
rect 28466 3614 28478 3666
rect 28530 3614 28542 3666
rect 32162 3614 32174 3666
rect 32226 3614 32238 3666
rect 36306 3614 36318 3666
rect 36370 3614 36382 3666
rect 38994 3614 39006 3666
rect 39058 3614 39070 3666
rect 41794 3614 41806 3666
rect 41858 3614 41870 3666
rect 44930 3614 44942 3666
rect 44994 3614 45006 3666
rect 48850 3614 48862 3666
rect 48914 3614 48926 3666
rect 21310 3602 21362 3614
rect 37886 3602 37938 3614
rect 44270 3602 44322 3614
rect 46846 3602 46898 3614
rect 51102 3602 51154 3614
rect 51550 3666 51602 3678
rect 51550 3602 51602 3614
rect 52110 3666 52162 3678
rect 68350 3666 68402 3678
rect 75630 3666 75682 3678
rect 53554 3614 53566 3666
rect 53618 3614 53630 3666
rect 57362 3614 57374 3666
rect 57426 3614 57438 3666
rect 59154 3614 59166 3666
rect 59218 3614 59230 3666
rect 61282 3614 61294 3666
rect 61346 3614 61358 3666
rect 63074 3614 63086 3666
rect 63138 3614 63150 3666
rect 65202 3614 65214 3666
rect 65266 3614 65278 3666
rect 71250 3614 71262 3666
rect 71314 3614 71326 3666
rect 72370 3614 72382 3666
rect 72434 3614 72446 3666
rect 76962 3614 76974 3666
rect 77026 3614 77038 3666
rect 52110 3602 52162 3614
rect 68350 3602 68402 3614
rect 75630 3602 75682 3614
rect 22542 3554 22594 3566
rect 22542 3490 22594 3502
rect 36990 3554 37042 3566
rect 52770 3502 52782 3554
rect 52834 3502 52846 3554
rect 54562 3502 54574 3554
rect 54626 3502 54638 3554
rect 56690 3502 56702 3554
rect 56754 3502 56766 3554
rect 58482 3502 58494 3554
rect 58546 3502 58558 3554
rect 60610 3502 60622 3554
rect 60674 3502 60686 3554
rect 62402 3502 62414 3554
rect 62466 3502 62478 3554
rect 64530 3502 64542 3554
rect 64594 3502 64606 3554
rect 67442 3502 67454 3554
rect 67506 3502 67518 3554
rect 76290 3502 76302 3554
rect 76354 3502 76366 3554
rect 36990 3490 37042 3502
rect 5742 3442 5794 3454
rect 3938 3390 3950 3442
rect 4002 3390 4014 3442
rect 5742 3378 5794 3390
rect 6862 3442 6914 3454
rect 9998 3442 10050 3454
rect 7858 3390 7870 3442
rect 7922 3390 7934 3442
rect 6862 3378 6914 3390
rect 9998 3378 10050 3390
rect 10894 3442 10946 3454
rect 13806 3442 13858 3454
rect 25342 3442 25394 3454
rect 29150 3442 29202 3454
rect 11666 3390 11678 3442
rect 11730 3390 11742 3442
rect 14690 3390 14702 3442
rect 14754 3390 14766 3442
rect 17602 3390 17614 3442
rect 17666 3390 17678 3442
rect 23426 3390 23438 3442
rect 23490 3390 23502 3442
rect 27458 3390 27470 3442
rect 27522 3390 27534 3442
rect 10894 3378 10946 3390
rect 13806 3378 13858 3390
rect 25342 3378 25394 3390
rect 29150 3378 29202 3390
rect 29710 3442 29762 3454
rect 33182 3442 33234 3454
rect 31378 3390 31390 3442
rect 31442 3390 31454 3442
rect 29710 3378 29762 3390
rect 33182 3378 33234 3390
rect 34414 3442 34466 3454
rect 38334 3442 38386 3454
rect 41246 3442 41298 3454
rect 43710 3442 43762 3454
rect 48190 3442 48242 3454
rect 69582 3442 69634 3454
rect 75070 3442 75122 3454
rect 35186 3390 35198 3442
rect 35250 3390 35262 3442
rect 39778 3390 39790 3442
rect 39842 3390 39854 3442
rect 42802 3390 42814 3442
rect 42866 3390 42878 3442
rect 45938 3390 45950 3442
rect 46002 3390 46014 3442
rect 49858 3390 49870 3442
rect 49922 3390 49934 3442
rect 55682 3390 55694 3442
rect 55746 3390 55758 3442
rect 66434 3390 66446 3442
rect 66498 3390 66510 3442
rect 70130 3390 70142 3442
rect 70194 3390 70206 3442
rect 73378 3390 73390 3442
rect 73442 3390 73454 3442
rect 34414 3378 34466 3390
rect 38334 3378 38386 3390
rect 41246 3378 41298 3390
rect 43710 3378 43762 3390
rect 48190 3378 48242 3390
rect 69582 3378 69634 3390
rect 75070 3378 75122 3390
rect 1344 3162 78624 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 78624 3162
rect 1344 3076 78624 3110
<< via1 >>
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 2046 75742 2098 75794
rect 75630 75742 75682 75794
rect 3054 75630 3106 75682
rect 3502 75630 3554 75682
rect 74958 75630 75010 75682
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 3054 74846 3106 74898
rect 74958 74846 75010 74898
rect 1934 74734 1986 74786
rect 3614 74734 3666 74786
rect 75630 74734 75682 74786
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 3278 74174 3330 74226
rect 74958 74174 75010 74226
rect 2270 73950 2322 74002
rect 3838 73950 3890 74002
rect 4174 73950 4226 74002
rect 76302 73950 76354 74002
rect 77310 73950 77362 74002
rect 73614 73838 73666 73890
rect 74062 73838 74114 73890
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 68910 73502 68962 73554
rect 73726 73502 73778 73554
rect 69022 73390 69074 73442
rect 73838 73390 73890 73442
rect 3054 73278 3106 73330
rect 4846 73278 4898 73330
rect 74958 73278 75010 73330
rect 76750 73278 76802 73330
rect 2046 73166 2098 73218
rect 3726 73166 3778 73218
rect 5406 73166 5458 73218
rect 69694 73166 69746 73218
rect 72382 73166 72434 73218
rect 74398 73166 74450 73218
rect 75966 73166 76018 73218
rect 77870 73166 77922 73218
rect 68798 73054 68850 73106
rect 73614 73054 73666 73106
rect 74174 73054 74226 73106
rect 74734 73054 74786 73106
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 74062 72606 74114 72658
rect 74174 72606 74226 72658
rect 3054 72494 3106 72546
rect 72158 72494 72210 72546
rect 73054 72494 73106 72546
rect 75070 72494 75122 72546
rect 1934 72382 1986 72434
rect 69358 72382 69410 72434
rect 70142 72382 70194 72434
rect 71822 72382 71874 72434
rect 73278 72382 73330 72434
rect 76078 72382 76130 72434
rect 3614 72270 3666 72322
rect 3950 72270 4002 72322
rect 69470 72270 69522 72322
rect 69582 72270 69634 72322
rect 73950 72270 74002 72322
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 72494 71934 72546 71986
rect 73390 71934 73442 71986
rect 74062 71934 74114 71986
rect 71262 71822 71314 71874
rect 71598 71822 71650 71874
rect 3054 71710 3106 71762
rect 4846 71710 4898 71762
rect 70814 71710 70866 71762
rect 72270 71710 72322 71762
rect 74958 71710 75010 71762
rect 76750 71710 76802 71762
rect 2046 71598 2098 71650
rect 3726 71598 3778 71650
rect 5406 71598 5458 71650
rect 73502 71598 73554 71650
rect 74174 71598 74226 71650
rect 75630 71598 75682 71650
rect 77870 71598 77922 71650
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 3278 71038 3330 71090
rect 74958 71038 75010 71090
rect 2158 70814 2210 70866
rect 70142 70814 70194 70866
rect 70590 70814 70642 70866
rect 70926 70814 70978 70866
rect 71598 70814 71650 70866
rect 71934 70814 71986 70866
rect 76302 70814 76354 70866
rect 3726 70702 3778 70754
rect 72494 70702 72546 70754
rect 72830 70702 72882 70754
rect 73726 70702 73778 70754
rect 74398 70702 74450 70754
rect 77310 70702 77362 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 71262 70366 71314 70418
rect 1934 70254 1986 70306
rect 3726 70254 3778 70306
rect 69918 70254 69970 70306
rect 76302 70254 76354 70306
rect 69470 70142 69522 70194
rect 70254 70142 70306 70194
rect 70926 70142 70978 70194
rect 71710 70142 71762 70194
rect 3278 70030 3330 70082
rect 75070 70030 75122 70082
rect 76862 70030 76914 70082
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 3278 69470 3330 69522
rect 72942 69470 72994 69522
rect 74958 69470 75010 69522
rect 2270 69246 2322 69298
rect 4174 69246 4226 69298
rect 69694 69246 69746 69298
rect 70254 69246 70306 69298
rect 70590 69246 70642 69298
rect 71150 69246 71202 69298
rect 74286 69246 74338 69298
rect 76302 69246 76354 69298
rect 3726 69134 3778 69186
rect 69358 69134 69410 69186
rect 77310 69134 77362 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 74510 68798 74562 68850
rect 2270 68686 2322 68738
rect 3950 68686 4002 68738
rect 68574 68686 68626 68738
rect 76302 68686 76354 68738
rect 3166 68462 3218 68514
rect 5294 68462 5346 68514
rect 67118 68462 67170 68514
rect 67678 68462 67730 68514
rect 69918 68462 69970 68514
rect 75182 68462 75234 68514
rect 76862 68462 76914 68514
rect 67790 68350 67842 68402
rect 68686 68350 68738 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 3502 68014 3554 68066
rect 4286 68014 4338 68066
rect 3278 67902 3330 67954
rect 3838 67902 3890 67954
rect 66782 67902 66834 67954
rect 67902 67902 67954 67954
rect 68462 67902 68514 67954
rect 69470 67902 69522 67954
rect 74958 67902 75010 67954
rect 2270 67678 2322 67730
rect 4174 67678 4226 67730
rect 67230 67678 67282 67730
rect 76302 67678 76354 67730
rect 77310 67678 77362 67730
rect 66334 67566 66386 67618
rect 67342 67566 67394 67618
rect 68014 67566 68066 67618
rect 69358 67566 69410 67618
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 68350 67230 68402 67282
rect 2158 67118 2210 67170
rect 67006 67118 67058 67170
rect 67454 67118 67506 67170
rect 69470 67118 69522 67170
rect 76302 67118 76354 67170
rect 3726 67006 3778 67058
rect 63534 67006 63586 67058
rect 65662 67006 65714 67058
rect 65886 67006 65938 67058
rect 68126 67006 68178 67058
rect 68462 67006 68514 67058
rect 68798 67006 68850 67058
rect 3278 66894 3330 66946
rect 63422 66894 63474 66946
rect 63982 66894 64034 66946
rect 65774 66894 65826 66946
rect 66110 66894 66162 66946
rect 68238 66894 68290 66946
rect 75182 66894 75234 66946
rect 76862 66894 76914 66946
rect 66334 66782 66386 66834
rect 66894 66782 66946 66834
rect 67342 66782 67394 66834
rect 67902 66782 67954 66834
rect 69358 66782 69410 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 68350 66446 68402 66498
rect 3278 66334 3330 66386
rect 64878 66334 64930 66386
rect 66894 66334 66946 66386
rect 68126 66334 68178 66386
rect 75070 66334 75122 66386
rect 65886 66222 65938 66274
rect 66222 66222 66274 66274
rect 66782 66222 66834 66274
rect 67902 66222 67954 66274
rect 2046 66110 2098 66162
rect 63310 66110 63362 66162
rect 63870 66110 63922 66162
rect 76302 66110 76354 66162
rect 3726 65998 3778 66050
rect 63422 65998 63474 66050
rect 65550 65998 65602 66050
rect 65662 65998 65714 66050
rect 65774 65998 65826 66050
rect 67678 65998 67730 66050
rect 67790 65998 67842 66050
rect 77310 65998 77362 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 68238 65662 68290 65714
rect 1934 65550 1986 65602
rect 64542 65550 64594 65602
rect 65886 65550 65938 65602
rect 76302 65550 76354 65602
rect 62078 65438 62130 65490
rect 65774 65438 65826 65490
rect 66110 65438 66162 65490
rect 68014 65438 68066 65490
rect 68462 65438 68514 65490
rect 68686 65438 68738 65490
rect 3278 65326 3330 65378
rect 3726 65326 3778 65378
rect 61966 65326 62018 65378
rect 62526 65326 62578 65378
rect 65998 65326 66050 65378
rect 66782 65326 66834 65378
rect 67118 65326 67170 65378
rect 68126 65326 68178 65378
rect 74958 65326 75010 65378
rect 76862 65326 76914 65378
rect 64654 65214 64706 65266
rect 65438 65214 65490 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 3278 64766 3330 64818
rect 66446 64766 66498 64818
rect 72942 64766 72994 64818
rect 74958 64766 75010 64818
rect 4174 64654 4226 64706
rect 63758 64654 63810 64706
rect 64318 64654 64370 64706
rect 65438 64654 65490 64706
rect 65774 64654 65826 64706
rect 66334 64654 66386 64706
rect 68238 64654 68290 64706
rect 1934 64542 1986 64594
rect 60734 64542 60786 64594
rect 61742 64542 61794 64594
rect 67006 64542 67058 64594
rect 67342 64542 67394 64594
rect 69358 64542 69410 64594
rect 74286 64542 74338 64594
rect 76302 64542 76354 64594
rect 3726 64430 3778 64482
rect 61854 64430 61906 64482
rect 62302 64430 62354 64482
rect 64206 64430 64258 64482
rect 65102 64430 65154 64482
rect 65214 64430 65266 64482
rect 65326 64430 65378 64482
rect 68574 64430 68626 64482
rect 69694 64430 69746 64482
rect 77310 64430 77362 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 65774 64094 65826 64146
rect 66334 64094 66386 64146
rect 67678 64094 67730 64146
rect 74510 64094 74562 64146
rect 2046 63982 2098 64034
rect 3950 63982 4002 64034
rect 61182 63982 61234 64034
rect 62526 63982 62578 64034
rect 63534 63982 63586 64034
rect 64654 63982 64706 64034
rect 76302 63982 76354 64034
rect 61070 63870 61122 63922
rect 61630 63870 61682 63922
rect 62302 63870 62354 63922
rect 63310 63870 63362 63922
rect 65550 63870 65602 63922
rect 66670 63870 66722 63922
rect 67342 63870 67394 63922
rect 76862 63870 76914 63922
rect 3278 63758 3330 63810
rect 5294 63758 5346 63810
rect 63422 63758 63474 63810
rect 63758 63758 63810 63810
rect 75182 63758 75234 63810
rect 63982 63646 64034 63698
rect 64542 63646 64594 63698
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 63870 63310 63922 63362
rect 3278 63198 3330 63250
rect 3838 63198 3890 63250
rect 59278 63198 59330 63250
rect 59838 63198 59890 63250
rect 63646 63198 63698 63250
rect 64990 63198 65042 63250
rect 65326 63198 65378 63250
rect 74958 63198 75010 63250
rect 63198 63086 63250 63138
rect 2158 62974 2210 63026
rect 61406 62974 61458 63026
rect 61966 62974 62018 63026
rect 76302 62974 76354 63026
rect 4174 62862 4226 62914
rect 59390 62862 59442 62914
rect 61518 62862 61570 62914
rect 63310 62862 63362 62914
rect 63422 62862 63474 62914
rect 65998 62862 66050 62914
rect 67006 62862 67058 62914
rect 77310 62862 77362 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 62750 62526 62802 62578
rect 62974 62526 63026 62578
rect 63758 62526 63810 62578
rect 1934 62414 1986 62466
rect 3726 62414 3778 62466
rect 61630 62414 61682 62466
rect 68238 62414 68290 62466
rect 68686 62414 68738 62466
rect 76302 62414 76354 62466
rect 59726 62302 59778 62354
rect 61182 62302 61234 62354
rect 62526 62302 62578 62354
rect 63982 62302 64034 62354
rect 64094 62302 64146 62354
rect 3278 62190 3330 62242
rect 59614 62190 59666 62242
rect 60174 62190 60226 62242
rect 61742 62190 61794 62242
rect 62302 62190 62354 62242
rect 62862 62190 62914 62242
rect 63870 62190 63922 62242
rect 64430 62190 64482 62242
rect 68126 62190 68178 62242
rect 75070 62190 75122 62242
rect 76862 62190 76914 62242
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 3278 61630 3330 61682
rect 74958 61630 75010 61682
rect 2046 61406 2098 61458
rect 60286 61406 60338 61458
rect 61518 61406 61570 61458
rect 63646 61406 63698 61458
rect 76302 61406 76354 61458
rect 3726 61294 3778 61346
rect 59054 61294 59106 61346
rect 59838 61294 59890 61346
rect 60398 61294 60450 61346
rect 61630 61294 61682 61346
rect 62190 61294 62242 61346
rect 62750 61294 62802 61346
rect 63310 61294 63362 61346
rect 77310 61294 77362 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 58494 60958 58546 61010
rect 62414 60958 62466 61010
rect 2158 60846 2210 60898
rect 59726 60846 59778 60898
rect 60734 60846 60786 60898
rect 62638 60846 62690 60898
rect 76302 60846 76354 60898
rect 57598 60734 57650 60786
rect 59390 60734 59442 60786
rect 60958 60734 61010 60786
rect 61966 60734 62018 60786
rect 3278 60622 3330 60674
rect 3726 60622 3778 60674
rect 57486 60622 57538 60674
rect 58046 60622 58098 60674
rect 60846 60622 60898 60674
rect 61182 60622 61234 60674
rect 62190 60622 62242 60674
rect 62526 60622 62578 60674
rect 64542 60622 64594 60674
rect 65326 60622 65378 60674
rect 74958 60622 75010 60674
rect 76862 60622 76914 60674
rect 61406 60510 61458 60562
rect 64430 60510 64482 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 3278 60062 3330 60114
rect 58830 60062 58882 60114
rect 60398 60062 60450 60114
rect 66558 60062 66610 60114
rect 67118 60062 67170 60114
rect 72942 60062 72994 60114
rect 74958 60062 75010 60114
rect 58046 59950 58098 60002
rect 59950 59950 60002 60002
rect 60622 59950 60674 60002
rect 66446 59950 66498 60002
rect 2270 59838 2322 59890
rect 56814 59838 56866 59890
rect 57150 59838 57202 59890
rect 58158 59838 58210 59890
rect 60174 59838 60226 59890
rect 61518 59838 61570 59890
rect 62078 59838 62130 59890
rect 74286 59838 74338 59890
rect 76302 59838 76354 59890
rect 3726 59726 3778 59778
rect 4174 59726 4226 59778
rect 56366 59726 56418 59778
rect 58942 59726 58994 59778
rect 60062 59726 60114 59778
rect 61406 59726 61458 59778
rect 77310 59726 77362 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 57822 59390 57874 59442
rect 59614 59390 59666 59442
rect 59838 59390 59890 59442
rect 61070 59390 61122 59442
rect 74510 59390 74562 59442
rect 1934 59278 1986 59330
rect 3950 59278 4002 59330
rect 76302 59278 76354 59330
rect 58382 59166 58434 59218
rect 58942 59166 58994 59218
rect 60286 59166 60338 59218
rect 61294 59166 61346 59218
rect 3278 59054 3330 59106
rect 5294 59054 5346 59106
rect 59726 59054 59778 59106
rect 60062 59054 60114 59106
rect 61854 59054 61906 59106
rect 75182 59054 75234 59106
rect 76862 59054 76914 59106
rect 58494 58942 58546 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 58606 58606 58658 58658
rect 3278 58494 3330 58546
rect 3838 58494 3890 58546
rect 75070 58494 75122 58546
rect 57262 58382 57314 58434
rect 58158 58382 58210 58434
rect 58270 58382 58322 58434
rect 2046 58270 2098 58322
rect 57150 58270 57202 58322
rect 59278 58270 59330 58322
rect 76302 58270 76354 58322
rect 4174 58158 4226 58210
rect 56702 58158 56754 58210
rect 57934 58158 57986 58210
rect 58046 58158 58098 58210
rect 59166 58158 59218 58210
rect 59838 58158 59890 58210
rect 77310 58158 77362 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 57822 57822 57874 57874
rect 63310 57822 63362 57874
rect 1934 57710 1986 57762
rect 62862 57710 62914 57762
rect 76302 57710 76354 57762
rect 54574 57598 54626 57650
rect 55134 57598 55186 57650
rect 56142 57598 56194 57650
rect 58046 57598 58098 57650
rect 58270 57598 58322 57650
rect 58494 57598 58546 57650
rect 3166 57486 3218 57538
rect 3726 57486 3778 57538
rect 56030 57486 56082 57538
rect 56590 57486 56642 57538
rect 57934 57486 57986 57538
rect 74958 57486 75010 57538
rect 76862 57486 76914 57538
rect 55246 57374 55298 57426
rect 62750 57374 62802 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 58046 57038 58098 57090
rect 3278 56926 3330 56978
rect 57822 56926 57874 56978
rect 74958 56926 75010 56978
rect 57598 56814 57650 56866
rect 2270 56702 2322 56754
rect 3726 56702 3778 56754
rect 56142 56702 56194 56754
rect 56590 56702 56642 56754
rect 58942 56702 58994 56754
rect 59502 56702 59554 56754
rect 76302 56702 76354 56754
rect 56702 56590 56754 56642
rect 57374 56590 57426 56642
rect 57486 56590 57538 56642
rect 58830 56590 58882 56642
rect 77310 56590 77362 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 57598 56254 57650 56306
rect 57822 56254 57874 56306
rect 2270 56142 2322 56194
rect 3726 56142 3778 56194
rect 76302 56142 76354 56194
rect 76862 56142 76914 56194
rect 53230 56030 53282 56082
rect 55358 56030 55410 56082
rect 55582 56030 55634 56082
rect 55694 56030 55746 56082
rect 56702 56030 56754 56082
rect 58046 56030 58098 56082
rect 58270 56030 58322 56082
rect 3278 55918 3330 55970
rect 53118 55918 53170 55970
rect 53678 55918 53730 55970
rect 54798 55918 54850 55970
rect 55470 55918 55522 55970
rect 57710 55918 57762 55970
rect 75070 55918 75122 55970
rect 56030 55806 56082 55858
rect 56590 55806 56642 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 57486 55470 57538 55522
rect 57710 55470 57762 55522
rect 3278 55358 3330 55410
rect 55694 55358 55746 55410
rect 57822 55358 57874 55410
rect 75182 55358 75234 55410
rect 54238 55246 54290 55298
rect 55246 55246 55298 55298
rect 55918 55246 55970 55298
rect 2046 55134 2098 55186
rect 50654 55134 50706 55186
rect 50766 55134 50818 55186
rect 54462 55134 54514 55186
rect 55470 55134 55522 55186
rect 56926 55134 56978 55186
rect 57262 55134 57314 55186
rect 76302 55134 76354 55186
rect 3726 55022 3778 55074
rect 51214 55022 51266 55074
rect 53678 55022 53730 55074
rect 55358 55022 55410 55074
rect 56366 55022 56418 55074
rect 77310 55022 77362 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 3726 54686 3778 54738
rect 56590 54686 56642 54738
rect 2158 54574 2210 54626
rect 52222 54574 52274 54626
rect 53902 54574 53954 54626
rect 54910 54574 54962 54626
rect 56030 54574 56082 54626
rect 56702 54574 56754 54626
rect 57374 54574 57426 54626
rect 76302 54574 76354 54626
rect 51550 54462 51602 54514
rect 52110 54462 52162 54514
rect 54686 54462 54738 54514
rect 55022 54462 55074 54514
rect 3278 54350 3330 54402
rect 52782 54350 52834 54402
rect 53342 54350 53394 54402
rect 54798 54350 54850 54402
rect 75070 54350 75122 54402
rect 76862 54350 76914 54402
rect 52894 54238 52946 54290
rect 54014 54238 54066 54290
rect 55358 54238 55410 54290
rect 55918 54238 55970 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 54238 53902 54290 53954
rect 56142 53902 56194 53954
rect 56478 53902 56530 53954
rect 3278 53790 3330 53842
rect 54462 53790 54514 53842
rect 56478 53790 56530 53842
rect 74958 53790 75010 53842
rect 52222 53678 52274 53730
rect 54686 53678 54738 53730
rect 2046 53566 2098 53618
rect 53566 53566 53618 53618
rect 55918 53566 55970 53618
rect 57038 53566 57090 53618
rect 57374 53566 57426 53618
rect 76302 53566 76354 53618
rect 3726 53454 3778 53506
rect 53454 53454 53506 53506
rect 54798 53454 54850 53506
rect 54910 53454 54962 53506
rect 55582 53454 55634 53506
rect 77310 53454 77362 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 58046 53118 58098 53170
rect 1934 53006 1986 53058
rect 51998 53006 52050 53058
rect 57598 53006 57650 53058
rect 76302 53006 76354 53058
rect 47742 52894 47794 52946
rect 48302 52894 48354 52946
rect 50542 52894 50594 52946
rect 51774 52894 51826 52946
rect 52894 52894 52946 52946
rect 53118 52894 53170 52946
rect 53566 52894 53618 52946
rect 3278 52782 3330 52834
rect 3726 52782 3778 52834
rect 50430 52782 50482 52834
rect 50990 52782 51042 52834
rect 53006 52782 53058 52834
rect 53342 52782 53394 52834
rect 54126 52782 54178 52834
rect 56702 52782 56754 52834
rect 75070 52782 75122 52834
rect 76862 52782 76914 52834
rect 48414 52670 48466 52722
rect 57486 52670 57538 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 54238 52334 54290 52386
rect 60510 52334 60562 52386
rect 3278 52222 3330 52274
rect 48302 52222 48354 52274
rect 48862 52222 48914 52274
rect 49534 52222 49586 52274
rect 51326 52222 51378 52274
rect 52670 52222 52722 52274
rect 54014 52222 54066 52274
rect 59278 52222 59330 52274
rect 60622 52222 60674 52274
rect 61406 52222 61458 52274
rect 75182 52222 75234 52274
rect 3726 52110 3778 52162
rect 50878 52110 50930 52162
rect 52334 52110 52386 52162
rect 56142 52110 56194 52162
rect 59390 52110 59442 52162
rect 59950 52110 60002 52162
rect 77310 52110 77362 52162
rect 2046 51998 2098 52050
rect 56366 51998 56418 52050
rect 56926 51998 56978 52050
rect 57262 51998 57314 52050
rect 76302 51998 76354 52050
rect 48414 51886 48466 51938
rect 49646 51886 49698 51938
rect 50542 51886 50594 51938
rect 51998 51886 52050 51938
rect 52110 51886 52162 51938
rect 52222 51886 52274 51938
rect 53566 51886 53618 51938
rect 53678 51886 53730 51938
rect 53790 51886 53842 51938
rect 55582 51886 55634 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 49534 51550 49586 51602
rect 51886 51550 51938 51602
rect 53342 51550 53394 51602
rect 2158 51438 2210 51490
rect 52110 51438 52162 51490
rect 53678 51438 53730 51490
rect 56590 51438 56642 51490
rect 76302 51438 76354 51490
rect 52334 51326 52386 51378
rect 52558 51326 52610 51378
rect 56254 51326 56306 51378
rect 3278 51214 3330 51266
rect 3726 51214 3778 51266
rect 51998 51214 52050 51266
rect 55694 51214 55746 51266
rect 75070 51214 75122 51266
rect 76862 51214 76914 51266
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 3278 50654 3330 50706
rect 48974 50654 49026 50706
rect 49422 50654 49474 50706
rect 50542 50654 50594 50706
rect 50878 50654 50930 50706
rect 72158 50654 72210 50706
rect 72606 50654 72658 50706
rect 73502 50654 73554 50706
rect 74062 50654 74114 50706
rect 74958 50654 75010 50706
rect 3726 50542 3778 50594
rect 51102 50542 51154 50594
rect 51662 50542 51714 50594
rect 51774 50542 51826 50594
rect 52334 50542 52386 50594
rect 53678 50542 53730 50594
rect 1934 50430 1986 50482
rect 49534 50430 49586 50482
rect 50430 50430 50482 50482
rect 50654 50430 50706 50482
rect 76302 50430 76354 50482
rect 77310 50430 77362 50482
rect 53454 50318 53506 50370
rect 72718 50318 72770 50370
rect 73390 50318 73442 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 50206 49982 50258 50034
rect 73838 49982 73890 50034
rect 2046 49870 2098 49922
rect 46734 49870 46786 49922
rect 50430 49870 50482 49922
rect 76302 49870 76354 49922
rect 46622 49758 46674 49810
rect 47182 49758 47234 49810
rect 50654 49758 50706 49810
rect 73390 49758 73442 49810
rect 73614 49758 73666 49810
rect 74062 49758 74114 49810
rect 3278 49646 3330 49698
rect 3726 49646 3778 49698
rect 48190 49646 48242 49698
rect 48750 49646 48802 49698
rect 50318 49646 50370 49698
rect 51550 49646 51602 49698
rect 51998 49646 52050 49698
rect 72606 49646 72658 49698
rect 73950 49646 74002 49698
rect 75182 49646 75234 49698
rect 76862 49646 76914 49698
rect 48302 49534 48354 49586
rect 50878 49534 50930 49586
rect 51438 49534 51490 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 3278 49086 3330 49138
rect 48078 49086 48130 49138
rect 49422 49086 49474 49138
rect 50654 49086 50706 49138
rect 51214 49086 51266 49138
rect 66670 49086 66722 49138
rect 67118 49086 67170 49138
rect 68350 49086 68402 49138
rect 69470 49086 69522 49138
rect 74958 49086 75010 49138
rect 49198 48974 49250 49026
rect 49870 48974 49922 49026
rect 68574 48974 68626 49026
rect 69358 48974 69410 49026
rect 1934 48862 1986 48914
rect 70030 48862 70082 48914
rect 76302 48862 76354 48914
rect 3838 48750 3890 48802
rect 4174 48750 4226 48802
rect 49646 48750 49698 48802
rect 49758 48750 49810 48802
rect 50542 48750 50594 48802
rect 67230 48750 67282 48802
rect 67902 48750 67954 48802
rect 68014 48750 68066 48802
rect 68126 48750 68178 48802
rect 73054 48750 73106 48802
rect 77310 48750 77362 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 48526 48414 48578 48466
rect 49646 48414 49698 48466
rect 68910 48414 68962 48466
rect 48414 48302 48466 48354
rect 3054 48190 3106 48242
rect 4846 48190 4898 48242
rect 49870 48190 49922 48242
rect 50094 48190 50146 48242
rect 50318 48190 50370 48242
rect 74958 48190 75010 48242
rect 76750 48190 76802 48242
rect 2046 48078 2098 48130
rect 3726 48078 3778 48130
rect 5406 48078 5458 48130
rect 47742 48078 47794 48130
rect 49758 48078 49810 48130
rect 74510 48078 74562 48130
rect 75966 48078 76018 48130
rect 77870 48078 77922 48130
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 49534 47630 49586 47682
rect 3054 47406 3106 47458
rect 74958 47406 75010 47458
rect 1934 47294 1986 47346
rect 47070 47294 47122 47346
rect 47406 47294 47458 47346
rect 48078 47294 48130 47346
rect 49646 47294 49698 47346
rect 50206 47294 50258 47346
rect 76078 47294 76130 47346
rect 3502 47182 3554 47234
rect 48414 47182 48466 47234
rect 48862 47182 48914 47234
rect 74398 47182 74450 47234
rect 77198 47182 77250 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 46398 46734 46450 46786
rect 47742 46734 47794 46786
rect 3054 46622 3106 46674
rect 45950 46622 46002 46674
rect 46734 46622 46786 46674
rect 47518 46622 47570 46674
rect 74958 46622 75010 46674
rect 2046 46510 2098 46562
rect 3614 46510 3666 46562
rect 48190 46510 48242 46562
rect 74510 46510 74562 46562
rect 75966 46510 76018 46562
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 3054 45838 3106 45890
rect 46062 45838 46114 45890
rect 46958 45838 47010 45890
rect 74958 45838 75010 45890
rect 1934 45726 1986 45778
rect 47182 45726 47234 45778
rect 76078 45726 76130 45778
rect 3502 45614 3554 45666
rect 45726 45614 45778 45666
rect 47742 45614 47794 45666
rect 48190 45614 48242 45666
rect 74398 45614 74450 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 44382 45278 44434 45330
rect 45614 45278 45666 45330
rect 46174 45166 46226 45218
rect 47406 45166 47458 45218
rect 3054 45054 3106 45106
rect 43934 45054 43986 45106
rect 44718 45054 44770 45106
rect 45390 45054 45442 45106
rect 46510 45054 46562 45106
rect 47182 45054 47234 45106
rect 74958 45054 75010 45106
rect 2046 44942 2098 44994
rect 3614 44942 3666 44994
rect 47854 44942 47906 44994
rect 48302 44942 48354 44994
rect 74510 44942 74562 44994
rect 75966 44942 76018 44994
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 3054 44270 3106 44322
rect 74958 44270 75010 44322
rect 1934 44158 1986 44210
rect 43710 44158 43762 44210
rect 44046 44158 44098 44210
rect 44606 44158 44658 44210
rect 45502 44158 45554 44210
rect 46398 44158 46450 44210
rect 76078 44158 76130 44210
rect 3502 44046 3554 44098
rect 45838 44046 45890 44098
rect 46734 44046 46786 44098
rect 74398 44046 74450 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 43038 43710 43090 43762
rect 44494 43710 44546 43762
rect 3054 43486 3106 43538
rect 42590 43486 42642 43538
rect 43374 43486 43426 43538
rect 44270 43486 44322 43538
rect 74958 43486 75010 43538
rect 1934 43374 1986 43426
rect 3614 43374 3666 43426
rect 44942 43374 44994 43426
rect 74510 43374 74562 43426
rect 76078 43374 76130 43426
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 3054 42702 3106 42754
rect 43486 42702 43538 42754
rect 74958 42702 75010 42754
rect 1934 42590 1986 42642
rect 3502 42590 3554 42642
rect 42366 42590 42418 42642
rect 42702 42590 42754 42642
rect 44270 42590 44322 42642
rect 76078 42590 76130 42642
rect 41918 42478 41970 42530
rect 43710 42478 43762 42530
rect 74398 42478 74450 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 41806 42142 41858 42194
rect 43150 42030 43202 42082
rect 3054 41918 3106 41970
rect 42142 41918 42194 41970
rect 42926 41918 42978 41970
rect 74958 41918 75010 41970
rect 1934 41806 1986 41858
rect 3614 41806 3666 41858
rect 43598 41806 43650 41858
rect 74510 41806 74562 41858
rect 76078 41806 76130 41858
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 3054 41134 3106 41186
rect 74958 41134 75010 41186
rect 1934 41022 1986 41074
rect 41022 41022 41074 41074
rect 41358 41022 41410 41074
rect 42142 41022 42194 41074
rect 76078 41022 76130 41074
rect 3502 40910 3554 40962
rect 40126 40910 40178 40962
rect 40574 40910 40626 40962
rect 42478 40910 42530 40962
rect 42926 40910 42978 40962
rect 74398 40910 74450 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 40350 40574 40402 40626
rect 42366 40574 42418 40626
rect 39454 40462 39506 40514
rect 41918 40462 41970 40514
rect 3054 40350 3106 40402
rect 3614 40350 3666 40402
rect 39790 40350 39842 40402
rect 40686 40350 40738 40402
rect 41582 40350 41634 40402
rect 42814 40350 42866 40402
rect 74510 40350 74562 40402
rect 74958 40350 75010 40402
rect 76078 40350 76130 40402
rect 1934 40238 1986 40290
rect 39006 40238 39058 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 1934 39566 1986 39618
rect 3054 39566 3106 39618
rect 74958 39566 75010 39618
rect 76078 39566 76130 39618
rect 3614 39454 3666 39506
rect 38894 39454 38946 39506
rect 39230 39454 39282 39506
rect 39790 39454 39842 39506
rect 40686 39454 40738 39506
rect 41022 39454 41074 39506
rect 38446 39342 38498 39394
rect 40126 39342 40178 39394
rect 41470 39342 41522 39394
rect 74510 39342 74562 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 1934 38894 1986 38946
rect 38334 38894 38386 38946
rect 39678 38894 39730 38946
rect 74510 38894 74562 38946
rect 76078 38894 76130 38946
rect 3054 38782 3106 38834
rect 3614 38782 3666 38834
rect 38670 38782 38722 38834
rect 39454 38782 39506 38834
rect 74958 38782 75010 38834
rect 37886 38670 37938 38722
rect 40350 38670 40402 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 1934 38110 1986 38162
rect 76078 38110 76130 38162
rect 3054 37998 3106 38050
rect 38894 37998 38946 38050
rect 74958 37998 75010 38050
rect 37998 37886 38050 37938
rect 40014 37886 40066 37938
rect 3614 37774 3666 37826
rect 37662 37774 37714 37826
rect 39118 37774 39170 37826
rect 39566 37774 39618 37826
rect 74510 37774 74562 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 1934 37326 1986 37378
rect 36990 37326 37042 37378
rect 38446 37326 38498 37378
rect 74510 37326 74562 37378
rect 76078 37326 76130 37378
rect 3054 37214 3106 37266
rect 36542 37214 36594 37266
rect 37326 37214 37378 37266
rect 38110 37214 38162 37266
rect 39342 37214 39394 37266
rect 74958 37214 75010 37266
rect 3614 37102 3666 37154
rect 38894 37102 38946 37154
rect 39118 36990 39170 37042
rect 39454 36990 39506 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 1934 36542 1986 36594
rect 76078 36542 76130 36594
rect 3054 36430 3106 36482
rect 36542 36430 36594 36482
rect 74958 36430 75010 36482
rect 35870 36318 35922 36370
rect 37550 36318 37602 36370
rect 3614 36206 3666 36258
rect 35422 36206 35474 36258
rect 36318 36206 36370 36258
rect 37886 36206 37938 36258
rect 74510 36206 74562 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 1934 35758 1986 35810
rect 34750 35758 34802 35810
rect 35646 35758 35698 35810
rect 36990 35758 37042 35810
rect 74510 35758 74562 35810
rect 76078 35758 76130 35810
rect 3054 35646 3106 35698
rect 4846 35646 4898 35698
rect 34974 35646 35026 35698
rect 35982 35646 36034 35698
rect 36654 35646 36706 35698
rect 37886 35646 37938 35698
rect 38334 35646 38386 35698
rect 74958 35646 75010 35698
rect 76750 35646 76802 35698
rect 3726 35534 3778 35586
rect 5406 35534 5458 35586
rect 37438 35534 37490 35586
rect 77870 35534 77922 35586
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 1934 34974 1986 35026
rect 3614 34974 3666 35026
rect 37438 34974 37490 35026
rect 76078 34974 76130 35026
rect 3054 34862 3106 34914
rect 35310 34862 35362 34914
rect 36094 34862 36146 34914
rect 74958 34862 75010 34914
rect 33854 34750 33906 34802
rect 34302 34750 34354 34802
rect 34638 34750 34690 34802
rect 36430 34750 36482 34802
rect 74510 34750 74562 34802
rect 4062 34638 4114 34690
rect 35534 34638 35586 34690
rect 77198 34638 77250 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 1934 34190 1986 34242
rect 33742 34190 33794 34242
rect 35086 34190 35138 34242
rect 74510 34190 74562 34242
rect 76078 34190 76130 34242
rect 3054 34078 3106 34130
rect 34078 34078 34130 34130
rect 34862 34078 34914 34130
rect 36206 34078 36258 34130
rect 74958 34078 75010 34130
rect 3614 33966 3666 34018
rect 35758 33966 35810 34018
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 1934 33406 1986 33458
rect 34862 33406 34914 33458
rect 76078 33406 76130 33458
rect 3054 33294 3106 33346
rect 33182 33294 33234 33346
rect 34078 33294 34130 33346
rect 74958 33294 75010 33346
rect 3614 33182 3666 33234
rect 32958 33182 33010 33234
rect 32510 33070 32562 33122
rect 34414 33070 34466 33122
rect 74510 33070 74562 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 34414 32734 34466 32786
rect 1934 32622 1986 32674
rect 32286 32622 32338 32674
rect 33966 32622 34018 32674
rect 74510 32622 74562 32674
rect 76078 32622 76130 32674
rect 3054 32510 3106 32562
rect 32510 32510 32562 32562
rect 33630 32510 33682 32562
rect 74958 32510 75010 32562
rect 3614 32398 3666 32450
rect 31838 32398 31890 32450
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 1934 31838 1986 31890
rect 33518 31838 33570 31890
rect 76078 31838 76130 31890
rect 3054 31726 3106 31778
rect 31950 31726 32002 31778
rect 32846 31726 32898 31778
rect 33966 31726 34018 31778
rect 74958 31726 75010 31778
rect 3614 31502 3666 31554
rect 30718 31502 30770 31554
rect 31166 31502 31218 31554
rect 31614 31502 31666 31554
rect 33070 31502 33122 31554
rect 74510 31502 74562 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 1934 31054 1986 31106
rect 30046 31054 30098 31106
rect 30942 31054 30994 31106
rect 32286 31054 32338 31106
rect 74510 31054 74562 31106
rect 76078 31054 76130 31106
rect 3054 30942 3106 30994
rect 4846 30942 4898 30994
rect 30382 30942 30434 30994
rect 31278 30942 31330 30994
rect 32062 30942 32114 30994
rect 32734 30942 32786 30994
rect 74958 30942 75010 30994
rect 76750 30942 76802 30994
rect 3726 30830 3778 30882
rect 5406 30830 5458 30882
rect 29374 30830 29426 30882
rect 77870 30830 77922 30882
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 1934 30270 1986 30322
rect 32174 30270 32226 30322
rect 3054 30158 3106 30210
rect 3614 30158 3666 30210
rect 74958 30158 75010 30210
rect 76078 30158 76130 30210
rect 29598 30046 29650 30098
rect 29934 30046 29986 30098
rect 30494 30046 30546 30098
rect 31390 30046 31442 30098
rect 31726 30046 31778 30098
rect 74510 30046 74562 30098
rect 4062 29934 4114 29986
rect 28814 29934 28866 29986
rect 30830 29934 30882 29986
rect 77198 29934 77250 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 1934 29486 1986 29538
rect 28926 29486 28978 29538
rect 30382 29486 30434 29538
rect 74510 29486 74562 29538
rect 76078 29486 76130 29538
rect 3054 29374 3106 29426
rect 28478 29374 28530 29426
rect 29262 29374 29314 29426
rect 30046 29374 30098 29426
rect 31054 29374 31106 29426
rect 74958 29374 75010 29426
rect 3614 29262 3666 29314
rect 31502 29262 31554 29314
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 1934 28702 1986 28754
rect 76078 28702 76130 28754
rect 3054 28590 3106 28642
rect 3614 28590 3666 28642
rect 27806 28590 27858 28642
rect 74510 28590 74562 28642
rect 74958 28590 75010 28642
rect 28254 28478 28306 28530
rect 28590 28478 28642 28530
rect 29598 28478 29650 28530
rect 29934 28366 29986 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 29374 28030 29426 28082
rect 1934 27918 1986 27970
rect 27582 27918 27634 27970
rect 28926 27918 28978 27970
rect 74510 27918 74562 27970
rect 76078 27918 76130 27970
rect 3054 27806 3106 27858
rect 27806 27806 27858 27858
rect 28590 27806 28642 27858
rect 29822 27806 29874 27858
rect 74958 27806 75010 27858
rect 3614 27694 3666 27746
rect 27134 27694 27186 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 1934 27134 1986 27186
rect 76078 27134 76130 27186
rect 3054 27022 3106 27074
rect 3614 27022 3666 27074
rect 74958 27022 75010 27074
rect 26462 26910 26514 26962
rect 27246 26910 27298 26962
rect 27918 26910 27970 26962
rect 28814 26910 28866 26962
rect 74510 26910 74562 26962
rect 26910 26798 26962 26850
rect 28254 26798 28306 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 1934 26350 1986 26402
rect 26238 26350 26290 26402
rect 27694 26350 27746 26402
rect 74510 26350 74562 26402
rect 76078 26350 76130 26402
rect 2942 26238 2994 26290
rect 4846 26238 4898 26290
rect 25790 26238 25842 26290
rect 26574 26238 26626 26290
rect 27358 26238 27410 26290
rect 74958 26238 75010 26290
rect 76974 26238 77026 26290
rect 3726 26126 3778 26178
rect 5406 26126 5458 26178
rect 25006 26126 25058 26178
rect 77870 26126 77922 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 1934 25566 1986 25618
rect 76078 25566 76130 25618
rect 3054 25454 3106 25506
rect 25566 25454 25618 25506
rect 26462 25454 26514 25506
rect 27582 25454 27634 25506
rect 74958 25454 75010 25506
rect 4062 25342 4114 25394
rect 24334 25342 24386 25394
rect 24670 25342 24722 25394
rect 25230 25342 25282 25394
rect 27134 25342 27186 25394
rect 3614 25230 3666 25282
rect 26686 25230 26738 25282
rect 74510 25230 74562 25282
rect 77198 25230 77250 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 1934 24782 1986 24834
rect 23662 24782 23714 24834
rect 24894 24782 24946 24834
rect 26126 24782 26178 24834
rect 76078 24782 76130 24834
rect 3054 24670 3106 24722
rect 22766 24670 22818 24722
rect 23102 24670 23154 24722
rect 23998 24670 24050 24722
rect 24558 24670 24610 24722
rect 25902 24670 25954 24722
rect 74510 24670 74562 24722
rect 74958 24670 75010 24722
rect 3614 24558 3666 24610
rect 26574 24558 26626 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 1934 23998 1986 24050
rect 76078 23998 76130 24050
rect 3054 23886 3106 23938
rect 74958 23886 75010 23938
rect 23998 23774 24050 23826
rect 25342 23774 25394 23826
rect 3614 23662 3666 23714
rect 23102 23662 23154 23714
rect 23662 23662 23714 23714
rect 24894 23662 24946 23714
rect 25678 23662 25730 23714
rect 26126 23662 26178 23714
rect 74510 23662 74562 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 1934 23214 1986 23266
rect 22430 23214 22482 23266
rect 23886 23214 23938 23266
rect 74510 23214 74562 23266
rect 76078 23214 76130 23266
rect 3054 23102 3106 23154
rect 22766 23102 22818 23154
rect 23662 23102 23714 23154
rect 74958 23102 75010 23154
rect 3614 22990 3666 23042
rect 24334 22990 24386 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 1934 22430 1986 22482
rect 76078 22430 76130 22482
rect 3054 22318 3106 22370
rect 23102 22318 23154 22370
rect 74958 22318 75010 22370
rect 22430 22206 22482 22258
rect 3614 22094 3666 22146
rect 22094 22094 22146 22146
rect 23326 22094 23378 22146
rect 23774 22094 23826 22146
rect 24334 22094 24386 22146
rect 74510 22094 74562 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 22654 21758 22706 21810
rect 1934 21646 1986 21698
rect 21758 21646 21810 21698
rect 23998 21646 24050 21698
rect 74510 21646 74562 21698
rect 76078 21646 76130 21698
rect 2942 21534 2994 21586
rect 4846 21534 4898 21586
rect 22094 21534 22146 21586
rect 23102 21534 23154 21586
rect 23662 21534 23714 21586
rect 24446 21534 24498 21586
rect 74958 21534 75010 21586
rect 76974 21534 77026 21586
rect 3726 21422 3778 21474
rect 5406 21422 5458 21474
rect 77870 21422 77922 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 1934 20862 1986 20914
rect 3614 20862 3666 20914
rect 76078 20862 76130 20914
rect 3054 20750 3106 20802
rect 21870 20750 21922 20802
rect 22766 20750 22818 20802
rect 23214 20750 23266 20802
rect 74958 20750 75010 20802
rect 4062 20638 4114 20690
rect 21646 20638 21698 20690
rect 20974 20526 21026 20578
rect 23550 20526 23602 20578
rect 74510 20526 74562 20578
rect 77198 20526 77250 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 19966 20190 20018 20242
rect 21198 20190 21250 20242
rect 1934 20078 1986 20130
rect 76078 20078 76130 20130
rect 3054 19966 3106 20018
rect 19518 19966 19570 20018
rect 20302 19966 20354 20018
rect 20862 19966 20914 20018
rect 21646 19966 21698 20018
rect 74958 19966 75010 20018
rect 3614 19854 3666 19906
rect 74510 19854 74562 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 1934 19294 1986 19346
rect 76078 19294 76130 19346
rect 3054 19182 3106 19234
rect 18958 19182 19010 19234
rect 74958 19182 75010 19234
rect 19630 19070 19682 19122
rect 19966 19070 20018 19122
rect 20526 19070 20578 19122
rect 21646 19070 21698 19122
rect 21982 19070 22034 19122
rect 74510 19070 74562 19122
rect 3614 18958 3666 19010
rect 18286 18958 18338 19010
rect 18734 18958 18786 19010
rect 20862 18958 20914 19010
rect 22430 18958 22482 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 21534 18622 21586 18674
rect 56254 18622 56306 18674
rect 1934 18510 1986 18562
rect 18622 18510 18674 18562
rect 21086 18510 21138 18562
rect 55582 18510 55634 18562
rect 3054 18398 3106 18450
rect 18958 18398 19010 18450
rect 20750 18398 20802 18450
rect 55806 18398 55858 18450
rect 56030 18398 56082 18450
rect 56254 18398 56306 18450
rect 74510 18398 74562 18450
rect 74958 18398 75010 18450
rect 76078 18398 76130 18450
rect 3614 18286 3666 18338
rect 18174 18286 18226 18338
rect 19742 18286 19794 18338
rect 20190 18286 20242 18338
rect 54574 18286 54626 18338
rect 55022 18286 55074 18338
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 20750 17838 20802 17890
rect 56254 17838 56306 17890
rect 1934 17726 1986 17778
rect 26238 17726 26290 17778
rect 55694 17726 55746 17778
rect 76078 17726 76130 17778
rect 3054 17614 3106 17666
rect 17166 17614 17218 17666
rect 20190 17614 20242 17666
rect 20302 17614 20354 17666
rect 20526 17614 20578 17666
rect 54126 17614 54178 17666
rect 55022 17614 55074 17666
rect 55582 17614 55634 17666
rect 56142 17614 56194 17666
rect 74958 17614 75010 17666
rect 17950 17502 18002 17554
rect 18510 17502 18562 17554
rect 18846 17502 18898 17554
rect 20862 17502 20914 17554
rect 25902 17502 25954 17554
rect 74510 17502 74562 17554
rect 3614 17390 3666 17442
rect 16382 17390 16434 17442
rect 17614 17390 17666 17442
rect 19294 17390 19346 17442
rect 21534 17390 21586 17442
rect 21982 17390 22034 17442
rect 24110 17390 24162 17442
rect 25006 17390 25058 17442
rect 25342 17390 25394 17442
rect 26126 17390 26178 17442
rect 53678 17390 53730 17442
rect 55134 17390 55186 17442
rect 55358 17390 55410 17442
rect 56702 17390 56754 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 19966 17054 20018 17106
rect 21086 17054 21138 17106
rect 24446 17054 24498 17106
rect 1934 16942 1986 16994
rect 15710 16942 15762 16994
rect 16606 16942 16658 16994
rect 18510 16942 18562 16994
rect 19518 16942 19570 16994
rect 26014 16942 26066 16994
rect 74510 16942 74562 16994
rect 76078 16942 76130 16994
rect 3054 16830 3106 16882
rect 4846 16830 4898 16882
rect 5406 16830 5458 16882
rect 16046 16830 16098 16882
rect 16942 16830 16994 16882
rect 18174 16830 18226 16882
rect 19182 16830 19234 16882
rect 20414 16830 20466 16882
rect 23662 16830 23714 16882
rect 24894 16830 24946 16882
rect 25678 16830 25730 16882
rect 25902 16830 25954 16882
rect 26238 16830 26290 16882
rect 26686 16830 26738 16882
rect 54574 16830 54626 16882
rect 74958 16830 75010 16882
rect 76750 16830 76802 16882
rect 77870 16830 77922 16882
rect 3726 16718 3778 16770
rect 17614 16718 17666 16770
rect 22318 16718 22370 16770
rect 22990 16718 23042 16770
rect 23214 16718 23266 16770
rect 22878 16606 22930 16658
rect 23438 16606 23490 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 18734 16270 18786 16322
rect 22878 16270 22930 16322
rect 23214 16270 23266 16322
rect 1934 16158 1986 16210
rect 3614 16158 3666 16210
rect 76078 16158 76130 16210
rect 3054 16046 3106 16098
rect 18062 16046 18114 16098
rect 18286 16046 18338 16098
rect 18510 16046 18562 16098
rect 18846 16046 18898 16098
rect 22654 16046 22706 16098
rect 74510 16046 74562 16098
rect 74958 16046 75010 16098
rect 15822 15934 15874 15986
rect 16158 15934 16210 15986
rect 19406 15934 19458 15986
rect 20190 15934 20242 15986
rect 4062 15822 4114 15874
rect 16718 15822 16770 15874
rect 17166 15822 17218 15874
rect 19742 15822 19794 15874
rect 23886 15822 23938 15874
rect 24334 15822 24386 15874
rect 77198 15822 77250 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 1934 15374 1986 15426
rect 14702 15374 14754 15426
rect 18174 15374 18226 15426
rect 56366 15374 56418 15426
rect 74510 15374 74562 15426
rect 76078 15374 76130 15426
rect 3054 15262 3106 15314
rect 15038 15262 15090 15314
rect 16382 15262 16434 15314
rect 56030 15262 56082 15314
rect 74958 15262 75010 15314
rect 3614 15150 3666 15202
rect 15486 15150 15538 15202
rect 17726 15150 17778 15202
rect 19070 15150 19122 15202
rect 55470 15150 55522 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 55358 14702 55410 14754
rect 1934 14590 1986 14642
rect 54126 14590 54178 14642
rect 76078 14590 76130 14642
rect 3054 14478 3106 14530
rect 54910 14478 54962 14530
rect 55134 14478 55186 14530
rect 56142 14478 56194 14530
rect 56814 14478 56866 14530
rect 74958 14478 75010 14530
rect 14366 14366 14418 14418
rect 3614 14254 3666 14306
rect 14030 14254 14082 14306
rect 14814 14254 14866 14306
rect 53678 14254 53730 14306
rect 55022 14254 55074 14306
rect 56366 14254 56418 14306
rect 74510 14254 74562 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 1934 13806 1986 13858
rect 12462 13806 12514 13858
rect 13358 13806 13410 13858
rect 55694 13806 55746 13858
rect 57822 13806 57874 13858
rect 74510 13806 74562 13858
rect 76078 13806 76130 13858
rect 3054 13694 3106 13746
rect 12798 13694 12850 13746
rect 13694 13694 13746 13746
rect 14142 13694 14194 13746
rect 54574 13694 54626 13746
rect 55358 13694 55410 13746
rect 57486 13694 57538 13746
rect 74958 13694 75010 13746
rect 3614 13582 3666 13634
rect 12014 13582 12066 13634
rect 56702 13582 56754 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 1934 13022 1986 13074
rect 55022 13022 55074 13074
rect 74510 13022 74562 13074
rect 76078 13022 76130 13074
rect 3054 12910 3106 12962
rect 74958 12910 75010 12962
rect 3614 12686 3666 12738
rect 12014 12686 12066 12738
rect 12910 12686 12962 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 1934 12238 1986 12290
rect 11342 12238 11394 12290
rect 12238 12238 12290 12290
rect 13470 12238 13522 12290
rect 74510 12238 74562 12290
rect 76078 12238 76130 12290
rect 3054 12126 3106 12178
rect 4846 12126 4898 12178
rect 11678 12126 11730 12178
rect 12574 12126 12626 12178
rect 13246 12126 13298 12178
rect 74958 12126 75010 12178
rect 76750 12126 76802 12178
rect 3726 12014 3778 12066
rect 13918 12014 13970 12066
rect 77870 12014 77922 12066
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 1934 11454 1986 11506
rect 3614 11454 3666 11506
rect 4062 11454 4114 11506
rect 76078 11454 76130 11506
rect 3054 11342 3106 11394
rect 12574 11342 12626 11394
rect 13582 11342 13634 11394
rect 74958 11342 75010 11394
rect 10670 11230 10722 11282
rect 11006 11230 11058 11282
rect 11566 11230 11618 11282
rect 12798 11230 12850 11282
rect 74510 11230 74562 11282
rect 11902 11118 11954 11170
rect 77198 11118 77250 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 1934 10670 1986 10722
rect 10110 10670 10162 10722
rect 11454 10670 11506 10722
rect 74510 10670 74562 10722
rect 76078 10670 76130 10722
rect 3054 10558 3106 10610
rect 10446 10558 10498 10610
rect 11118 10558 11170 10610
rect 74958 10558 75010 10610
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 1934 9886 1986 9938
rect 76078 9886 76130 9938
rect 3054 9774 3106 9826
rect 9662 9774 9714 9826
rect 74958 9774 75010 9826
rect 9438 9662 9490 9714
rect 10558 9662 10610 9714
rect 10894 9550 10946 9602
rect 74510 9550 74562 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 1934 9102 1986 9154
rect 8654 9102 8706 9154
rect 10222 9102 10274 9154
rect 74510 9102 74562 9154
rect 76078 9102 76130 9154
rect 3054 8990 3106 9042
rect 8990 8990 9042 9042
rect 9886 8990 9938 9042
rect 74958 8990 75010 9042
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 1934 8318 1986 8370
rect 76078 8318 76130 8370
rect 3054 8206 3106 8258
rect 74958 8206 75010 8258
rect 8094 8094 8146 8146
rect 8430 8094 8482 8146
rect 9102 8094 9154 8146
rect 9438 7982 9490 8034
rect 74510 7982 74562 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 1934 7534 1986 7586
rect 6526 7534 6578 7586
rect 7422 7534 7474 7586
rect 8766 7534 8818 7586
rect 74510 7534 74562 7586
rect 76078 7534 76130 7586
rect 3054 7422 3106 7474
rect 4846 7422 4898 7474
rect 6862 7422 6914 7474
rect 7646 7422 7698 7474
rect 8430 7422 8482 7474
rect 74958 7422 75010 7474
rect 76750 7422 76802 7474
rect 3726 7310 3778 7362
rect 18062 7310 18114 7362
rect 77870 7310 77922 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 1934 6750 1986 6802
rect 16270 6750 16322 6802
rect 19518 6750 19570 6802
rect 23662 6750 23714 6802
rect 27022 6750 27074 6802
rect 70030 6750 70082 6802
rect 3054 6638 3106 6690
rect 6302 6638 6354 6690
rect 6974 6638 7026 6690
rect 7870 6638 7922 6690
rect 68686 6638 68738 6690
rect 69358 6638 69410 6690
rect 74958 6638 75010 6690
rect 76078 6638 76130 6690
rect 6078 6526 6130 6578
rect 7310 6526 7362 6578
rect 17278 6526 17330 6578
rect 18510 6526 18562 6578
rect 22430 6526 22482 6578
rect 28030 6526 28082 6578
rect 66782 6526 66834 6578
rect 77198 6526 77250 6578
rect 8206 6414 8258 6466
rect 8654 6414 8706 6466
rect 20638 6414 20690 6466
rect 21870 6414 21922 6466
rect 26574 6414 26626 6466
rect 31054 6414 31106 6466
rect 74510 6414 74562 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 53006 6078 53058 6130
rect 54238 6078 54290 6130
rect 55022 6078 55074 6130
rect 55358 6078 55410 6130
rect 57374 6078 57426 6130
rect 58158 6078 58210 6130
rect 58718 6078 58770 6130
rect 59166 6078 59218 6130
rect 59614 6078 59666 6130
rect 60286 6078 60338 6130
rect 61182 6078 61234 6130
rect 61518 6078 61570 6130
rect 62078 6078 62130 6130
rect 64206 6078 64258 6130
rect 65326 6078 65378 6130
rect 65774 6078 65826 6130
rect 66334 6078 66386 6130
rect 66782 6078 66834 6130
rect 1934 5966 1986 6018
rect 4622 5966 4674 6018
rect 6862 5966 6914 6018
rect 8654 5966 8706 6018
rect 15934 5966 15986 6018
rect 20302 5966 20354 6018
rect 21982 5966 22034 6018
rect 23102 5966 23154 6018
rect 28702 5966 28754 6018
rect 30382 5966 30434 6018
rect 32398 5966 32450 6018
rect 35198 5966 35250 6018
rect 47294 5966 47346 6018
rect 76078 5966 76130 6018
rect 3054 5854 3106 5906
rect 4958 5854 5010 5906
rect 18398 5854 18450 5906
rect 50542 5854 50594 5906
rect 51214 5854 51266 5906
rect 67342 5854 67394 5906
rect 70142 5854 70194 5906
rect 70814 5854 70866 5906
rect 74958 5854 75010 5906
rect 76750 5854 76802 5906
rect 4174 5742 4226 5794
rect 5518 5742 5570 5794
rect 7758 5742 7810 5794
rect 11118 5742 11170 5794
rect 11902 5742 11954 5794
rect 13470 5742 13522 5794
rect 13918 5742 13970 5794
rect 14478 5742 14530 5794
rect 16718 5742 16770 5794
rect 17950 5742 18002 5794
rect 18958 5742 19010 5794
rect 20974 5742 21026 5794
rect 24222 5742 24274 5794
rect 27358 5742 27410 5794
rect 29374 5742 29426 5794
rect 31614 5742 31666 5794
rect 33518 5742 33570 5794
rect 34638 5742 34690 5794
rect 36318 5742 36370 5794
rect 38782 5742 38834 5794
rect 40238 5742 40290 5794
rect 42254 5742 42306 5794
rect 45390 5742 45442 5794
rect 46734 5742 46786 5794
rect 48414 5742 48466 5794
rect 49646 5742 49698 5794
rect 51662 5742 51714 5794
rect 55806 5742 55858 5794
rect 56366 5742 56418 5794
rect 68014 5742 68066 5794
rect 69246 5742 69298 5794
rect 73390 5742 73442 5794
rect 73838 5742 73890 5794
rect 74510 5742 74562 5794
rect 77870 5742 77922 5794
rect 73502 5630 73554 5682
rect 73838 5630 73890 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 1934 5182 1986 5234
rect 7646 5182 7698 5234
rect 9662 5182 9714 5234
rect 11566 5182 11618 5234
rect 16718 5182 16770 5234
rect 18622 5182 18674 5234
rect 20862 5182 20914 5234
rect 21982 5182 22034 5234
rect 24670 5182 24722 5234
rect 25454 5182 25506 5234
rect 27582 5182 27634 5234
rect 29486 5182 29538 5234
rect 31278 5182 31330 5234
rect 34526 5182 34578 5234
rect 35310 5182 35362 5234
rect 39678 5182 39730 5234
rect 40462 5182 40514 5234
rect 43710 5182 43762 5234
rect 46958 5182 47010 5234
rect 48750 5182 48802 5234
rect 51998 5182 52050 5234
rect 55918 5182 55970 5234
rect 59950 5182 60002 5234
rect 62078 5182 62130 5234
rect 67790 5182 67842 5234
rect 70142 5182 70194 5234
rect 73278 5182 73330 5234
rect 74062 5182 74114 5234
rect 3054 5070 3106 5122
rect 14478 5070 14530 5122
rect 21646 5070 21698 5122
rect 22766 5070 22818 5122
rect 30830 5070 30882 5122
rect 37438 5070 37490 5122
rect 44830 5070 44882 5122
rect 49646 5070 49698 5122
rect 50766 5070 50818 5122
rect 51326 5070 51378 5122
rect 54462 5070 54514 5122
rect 55246 5070 55298 5122
rect 57374 5070 57426 5122
rect 58494 5070 58546 5122
rect 59278 5070 59330 5122
rect 61406 5070 61458 5122
rect 64542 5070 64594 5122
rect 66334 5070 66386 5122
rect 67118 5070 67170 5122
rect 69358 5070 69410 5122
rect 71598 5070 71650 5122
rect 76526 5070 76578 5122
rect 4622 4958 4674 5010
rect 6414 4958 6466 5010
rect 8430 4958 8482 5010
rect 10446 4958 10498 5010
rect 12462 4958 12514 5010
rect 13694 4958 13746 5010
rect 14030 4958 14082 5010
rect 15822 4958 15874 5010
rect 17838 4958 17890 5010
rect 19518 4958 19570 5010
rect 23774 4958 23826 5010
rect 26686 4958 26738 5010
rect 28366 4958 28418 5010
rect 29934 4958 29986 5010
rect 32286 4958 32338 5010
rect 33742 4958 33794 5010
rect 36318 4958 36370 5010
rect 38670 4958 38722 5010
rect 41470 4958 41522 5010
rect 42590 4958 42642 5010
rect 45614 4958 45666 5010
rect 47630 4958 47682 5010
rect 53566 4958 53618 5010
rect 63422 4958 63474 5010
rect 65438 4958 65490 5010
rect 72270 4958 72322 5010
rect 75070 4958 75122 5010
rect 4958 4846 5010 4898
rect 6750 4846 6802 4898
rect 37998 4846 38050 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 4622 4510 4674 4562
rect 16830 4510 16882 4562
rect 69470 4510 69522 4562
rect 6750 4398 6802 4450
rect 7982 4398 8034 4450
rect 11230 4398 11282 4450
rect 12686 4398 12738 4450
rect 14366 4398 14418 4450
rect 19854 4398 19906 4450
rect 21870 4398 21922 4450
rect 24782 4398 24834 4450
rect 28702 4398 28754 4450
rect 29822 4398 29874 4450
rect 32734 4398 32786 4450
rect 35534 4398 35586 4450
rect 38110 4398 38162 4450
rect 40126 4398 40178 4450
rect 41694 4398 41746 4450
rect 44606 4398 44658 4450
rect 45726 4398 45778 4450
rect 50542 4398 50594 4450
rect 70814 4398 70866 4450
rect 74398 4398 74450 4450
rect 76414 4398 76466 4450
rect 4846 4286 4898 4338
rect 9662 4286 9714 4338
rect 26014 4286 26066 4338
rect 33518 4286 33570 4338
rect 51550 4286 51602 4338
rect 53342 4286 53394 4338
rect 56142 4286 56194 4338
rect 57486 4286 57538 4338
rect 59390 4286 59442 4338
rect 61070 4286 61122 4338
rect 63870 4286 63922 4338
rect 64542 4286 64594 4338
rect 65662 4286 65714 4338
rect 68238 4286 68290 4338
rect 68910 4286 68962 4338
rect 5742 4174 5794 4226
rect 8990 4174 9042 4226
rect 10446 4174 10498 4226
rect 13582 4174 13634 4226
rect 17614 4174 17666 4226
rect 18062 4174 18114 4226
rect 18846 4174 18898 4226
rect 20750 4174 20802 4226
rect 22654 4174 22706 4226
rect 23438 4174 23490 4226
rect 25566 4174 25618 4226
rect 26798 4174 26850 4226
rect 27470 4174 27522 4226
rect 30606 4174 30658 4226
rect 31502 4174 31554 4226
rect 33966 4174 34018 4226
rect 34526 4174 34578 4226
rect 36542 4174 36594 4226
rect 37326 4174 37378 4226
rect 39118 4174 39170 4226
rect 42814 4174 42866 4226
rect 43598 4174 43650 4226
rect 46846 4174 46898 4226
rect 47518 4174 47570 4226
rect 48750 4174 48802 4226
rect 49534 4174 49586 4226
rect 52222 4174 52274 4226
rect 54014 4174 54066 4226
rect 55470 4174 55522 4226
rect 58158 4174 58210 4226
rect 59950 4174 60002 4226
rect 61742 4174 61794 4226
rect 62974 4174 63026 4226
rect 66110 4174 66162 4226
rect 67342 4174 67394 4226
rect 70254 4174 70306 4226
rect 71934 4174 71986 4226
rect 72718 4174 72770 4226
rect 73390 4174 73442 4226
rect 75406 4174 75458 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 16830 3726 16882 3778
rect 4958 3614 5010 3666
rect 8878 3614 8930 3666
rect 9550 3614 9602 3666
rect 12574 3614 12626 3666
rect 19742 3614 19794 3666
rect 21310 3614 21362 3666
rect 24334 3614 24386 3666
rect 28478 3614 28530 3666
rect 32174 3614 32226 3666
rect 36318 3614 36370 3666
rect 37886 3614 37938 3666
rect 39006 3614 39058 3666
rect 41806 3614 41858 3666
rect 44270 3614 44322 3666
rect 44942 3614 44994 3666
rect 46846 3614 46898 3666
rect 48862 3614 48914 3666
rect 51102 3614 51154 3666
rect 51550 3614 51602 3666
rect 52110 3614 52162 3666
rect 53566 3614 53618 3666
rect 57374 3614 57426 3666
rect 59166 3614 59218 3666
rect 61294 3614 61346 3666
rect 63086 3614 63138 3666
rect 65214 3614 65266 3666
rect 68350 3614 68402 3666
rect 71262 3614 71314 3666
rect 72382 3614 72434 3666
rect 75630 3614 75682 3666
rect 76974 3614 77026 3666
rect 22542 3502 22594 3554
rect 36990 3502 37042 3554
rect 52782 3502 52834 3554
rect 54574 3502 54626 3554
rect 56702 3502 56754 3554
rect 58494 3502 58546 3554
rect 60622 3502 60674 3554
rect 62414 3502 62466 3554
rect 64542 3502 64594 3554
rect 67454 3502 67506 3554
rect 76302 3502 76354 3554
rect 3950 3390 4002 3442
rect 5742 3390 5794 3442
rect 6862 3390 6914 3442
rect 7870 3390 7922 3442
rect 9998 3390 10050 3442
rect 10894 3390 10946 3442
rect 11678 3390 11730 3442
rect 13806 3390 13858 3442
rect 14702 3390 14754 3442
rect 17614 3390 17666 3442
rect 23438 3390 23490 3442
rect 25342 3390 25394 3442
rect 27470 3390 27522 3442
rect 29150 3390 29202 3442
rect 29710 3390 29762 3442
rect 31390 3390 31442 3442
rect 33182 3390 33234 3442
rect 34414 3390 34466 3442
rect 35198 3390 35250 3442
rect 38334 3390 38386 3442
rect 39790 3390 39842 3442
rect 41246 3390 41298 3442
rect 42814 3390 42866 3442
rect 43710 3390 43762 3442
rect 45950 3390 46002 3442
rect 48190 3390 48242 3442
rect 49870 3390 49922 3442
rect 55694 3390 55746 3442
rect 66446 3390 66498 3442
rect 69582 3390 69634 3442
rect 70142 3390 70194 3442
rect 73390 3390 73442 3442
rect 75070 3390 75122 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 2044 75794 2100 75806
rect 75628 75796 75684 75806
rect 2044 75742 2046 75794
rect 2098 75742 2100 75794
rect 1932 74786 1988 74798
rect 1932 74734 1934 74786
rect 1986 74734 1988 74786
rect 1932 73220 1988 74734
rect 2044 74564 2100 75742
rect 75516 75794 75684 75796
rect 75516 75742 75630 75794
rect 75682 75742 75684 75794
rect 75516 75740 75684 75742
rect 3052 75684 3108 75694
rect 3500 75684 3556 75694
rect 3052 75682 3556 75684
rect 3052 75630 3054 75682
rect 3106 75630 3502 75682
rect 3554 75630 3556 75682
rect 3052 75628 3556 75630
rect 3052 75618 3108 75628
rect 3052 74900 3108 74910
rect 3052 74806 3108 74844
rect 2044 74498 2100 74508
rect 3276 74228 3332 74238
rect 3276 74226 3444 74228
rect 3276 74174 3278 74226
rect 3330 74174 3444 74226
rect 3276 74172 3444 74174
rect 3276 74162 3332 74172
rect 2268 74004 2324 74014
rect 2268 73910 2324 73948
rect 3052 73332 3108 73342
rect 3388 73332 3444 74172
rect 3500 73556 3556 75628
rect 74956 75682 75012 75694
rect 74956 75630 74958 75682
rect 75010 75630 75012 75682
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 73724 75124 73780 75134
rect 3500 73490 3556 73500
rect 3612 74900 3668 74910
rect 3612 74786 3668 74844
rect 3612 74734 3614 74786
rect 3666 74734 3668 74786
rect 3388 73276 3556 73332
rect 3052 73238 3108 73276
rect 1932 73154 1988 73164
rect 2044 73218 2100 73230
rect 2044 73166 2046 73218
rect 2098 73166 2100 73218
rect 1932 72436 1988 72446
rect 1820 72434 1988 72436
rect 1820 72382 1934 72434
rect 1986 72382 1988 72434
rect 1820 72380 1988 72382
rect 1820 70532 1876 72380
rect 1932 72370 1988 72380
rect 2044 71876 2100 73166
rect 3052 72546 3108 72558
rect 3052 72494 3054 72546
rect 3106 72494 3108 72546
rect 3052 72324 3108 72494
rect 3052 72258 3108 72268
rect 2044 71810 2100 71820
rect 3052 71764 3108 71774
rect 1820 70466 1876 70476
rect 2044 71650 2100 71662
rect 2044 71598 2046 71650
rect 2098 71598 2100 71650
rect 1932 70308 1988 70318
rect 1820 70252 1932 70308
rect 1708 69300 1764 69310
rect 1708 67060 1764 69244
rect 1820 67844 1876 70252
rect 1932 70176 1988 70252
rect 2044 69860 2100 71598
rect 2044 69794 2100 69804
rect 2156 70866 2212 70878
rect 2156 70814 2158 70866
rect 2210 70814 2212 70866
rect 2156 70756 2212 70814
rect 2156 69188 2212 70700
rect 2268 69300 2324 69310
rect 2268 69206 2324 69244
rect 2156 69122 2212 69132
rect 3052 69188 3108 71708
rect 3276 71090 3332 71102
rect 3276 71038 3278 71090
rect 3330 71038 3332 71090
rect 3276 70980 3332 71038
rect 3388 70980 3444 70990
rect 3276 70924 3388 70980
rect 3388 70914 3444 70924
rect 3276 70082 3332 70094
rect 3276 70030 3278 70082
rect 3330 70030 3332 70082
rect 3276 69972 3332 70030
rect 3388 69972 3444 69982
rect 3276 69916 3388 69972
rect 3388 69906 3444 69916
rect 3276 69522 3332 69534
rect 3276 69470 3278 69522
rect 3330 69470 3332 69522
rect 3276 69412 3332 69470
rect 3276 69356 3444 69412
rect 3052 69122 3108 69132
rect 2268 68740 2324 68750
rect 1820 67778 1876 67788
rect 2156 68684 2268 68740
rect 2156 67396 2212 68684
rect 2268 68646 2324 68684
rect 3164 68514 3220 68526
rect 3164 68462 3166 68514
rect 3218 68462 3220 68514
rect 2156 67330 2212 67340
rect 2268 67732 2324 67742
rect 3164 67732 3220 68462
rect 3388 68292 3444 69356
rect 3500 68516 3556 73276
rect 3612 72660 3668 74734
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 3836 74002 3892 74014
rect 3836 73950 3838 74002
rect 3890 73950 3892 74002
rect 3836 73332 3892 73950
rect 4172 74004 4228 74014
rect 4172 73910 4228 73948
rect 73612 73892 73668 73902
rect 73500 73890 73668 73892
rect 73500 73838 73614 73890
rect 73666 73838 73668 73890
rect 73500 73836 73668 73838
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 68908 73556 68964 73566
rect 68908 73462 68964 73500
rect 69020 73444 69076 73454
rect 69020 73350 69076 73388
rect 3612 72594 3668 72604
rect 3724 73218 3780 73230
rect 3724 73166 3726 73218
rect 3778 73166 3780 73218
rect 3724 72548 3780 73166
rect 3724 72482 3780 72492
rect 3612 72322 3668 72334
rect 3612 72270 3614 72322
rect 3666 72270 3668 72322
rect 3612 71764 3668 72270
rect 3836 72212 3892 73276
rect 4844 73330 4900 73342
rect 4844 73278 4846 73330
rect 4898 73278 4900 73330
rect 4844 73220 4900 73278
rect 72492 73332 72548 73342
rect 4844 73154 4900 73164
rect 5404 73220 5460 73230
rect 5404 73126 5460 73164
rect 69692 73218 69748 73230
rect 69692 73166 69694 73218
rect 69746 73166 69748 73218
rect 68460 73108 68516 73118
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 3836 72146 3892 72156
rect 3948 72324 4004 72334
rect 3612 71698 3668 71708
rect 3724 71650 3780 71662
rect 3724 71598 3726 71650
rect 3778 71598 3780 71650
rect 3724 71204 3780 71598
rect 3724 71138 3780 71148
rect 3836 70980 3892 70990
rect 3724 70756 3780 70766
rect 3724 70662 3780 70700
rect 3724 70308 3780 70318
rect 3724 70214 3780 70252
rect 3724 69186 3780 69198
rect 3724 69134 3726 69186
rect 3778 69134 3780 69186
rect 3724 68740 3780 69134
rect 3724 68674 3780 68684
rect 3836 68628 3892 70924
rect 3948 70308 4004 72268
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 4844 71762 4900 71774
rect 4844 71710 4846 71762
rect 4898 71710 4900 71762
rect 4844 71652 4900 71710
rect 4844 71586 4900 71596
rect 5404 71652 5460 71662
rect 5404 71558 5460 71596
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 3948 70242 4004 70252
rect 4060 69972 4116 69982
rect 3836 68562 3892 68572
rect 3948 68738 4004 68750
rect 3948 68686 3950 68738
rect 4002 68686 4004 68738
rect 3948 68516 4004 68686
rect 3500 68460 3780 68516
rect 3388 68236 3668 68292
rect 3500 68066 3556 68078
rect 3500 68014 3502 68066
rect 3554 68014 3556 68066
rect 3276 67956 3332 67966
rect 3500 67956 3556 68014
rect 3276 67954 3556 67956
rect 3276 67902 3278 67954
rect 3330 67902 3556 67954
rect 3276 67900 3556 67902
rect 3276 67890 3332 67900
rect 3164 67676 3444 67732
rect 1708 66994 1764 67004
rect 2156 67170 2212 67182
rect 2156 67118 2158 67170
rect 2210 67118 2212 67170
rect 2156 67060 2212 67118
rect 2044 66162 2100 66174
rect 2044 66110 2046 66162
rect 2098 66110 2100 66162
rect 2044 66052 2100 66110
rect 1932 65604 1988 65614
rect 1820 65602 1988 65604
rect 1820 65550 1934 65602
rect 1986 65550 1988 65602
rect 1820 65548 1988 65550
rect 1820 65380 1876 65548
rect 1932 65538 1988 65548
rect 1820 63140 1876 65324
rect 1820 63074 1876 63084
rect 1932 64708 1988 64718
rect 1932 64594 1988 64652
rect 1932 64542 1934 64594
rect 1986 64542 1988 64594
rect 1932 62692 1988 64542
rect 2044 64484 2100 65996
rect 2156 65156 2212 67004
rect 2268 65828 2324 67676
rect 3388 67228 3444 67676
rect 3612 67620 3668 68236
rect 3724 67732 3780 68460
rect 3836 67956 3892 67966
rect 3948 67956 4004 68460
rect 3836 67954 4004 67956
rect 3836 67902 3838 67954
rect 3890 67902 4004 67954
rect 3836 67900 4004 67902
rect 3836 67890 3892 67900
rect 3724 67676 4004 67732
rect 3612 67564 3892 67620
rect 3388 67172 3668 67228
rect 3276 66948 3332 66958
rect 3276 66946 3556 66948
rect 3276 66894 3278 66946
rect 3330 66894 3556 66946
rect 3276 66892 3556 66894
rect 3276 66882 3332 66892
rect 3276 66386 3332 66398
rect 3276 66334 3278 66386
rect 3330 66334 3332 66386
rect 3276 65940 3332 66334
rect 3276 65884 3444 65940
rect 2268 65762 2324 65772
rect 3388 65492 3444 65884
rect 3388 65426 3444 65436
rect 3276 65378 3332 65390
rect 3276 65326 3278 65378
rect 3330 65326 3332 65378
rect 3276 65268 3332 65326
rect 3276 65212 3444 65268
rect 2156 65090 2212 65100
rect 3388 65156 3444 65212
rect 3388 65090 3444 65100
rect 3276 64820 3332 64830
rect 3276 64818 3444 64820
rect 3276 64766 3278 64818
rect 3330 64766 3444 64818
rect 3276 64764 3444 64766
rect 3276 64754 3332 64764
rect 2044 64418 2100 64428
rect 3388 64372 3444 64764
rect 3500 64596 3556 66892
rect 3612 66164 3668 67172
rect 3724 67060 3780 67070
rect 3724 66966 3780 67004
rect 3836 66948 3892 67564
rect 3948 67228 4004 67676
rect 4060 67620 4116 69916
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 66780 69412 66836 69422
rect 4172 69300 4228 69310
rect 4172 69206 4228 69244
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 5292 68514 5348 68526
rect 5292 68462 5294 68514
rect 5346 68462 5348 68514
rect 5292 68404 5348 68462
rect 5292 68338 5348 68348
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 4284 68066 4340 68078
rect 4284 68014 4286 68066
rect 4338 68014 4340 68066
rect 4172 67732 4228 67742
rect 4172 67638 4228 67676
rect 4060 67554 4116 67564
rect 3948 67172 4116 67228
rect 3836 66882 3892 66892
rect 3612 66098 3668 66108
rect 3724 66052 3780 66062
rect 3724 65958 3780 65996
rect 3724 65380 3780 65390
rect 3724 65286 3780 65324
rect 3500 64530 3556 64540
rect 3724 64482 3780 64494
rect 3724 64430 3726 64482
rect 3778 64430 3780 64482
rect 3388 64316 3668 64372
rect 1932 62626 1988 62636
rect 2044 64260 2100 64270
rect 2044 64034 2100 64204
rect 2044 63982 2046 64034
rect 2098 63982 2100 64034
rect 1932 62468 1988 62478
rect 1820 62412 1932 62468
rect 1820 60452 1876 62412
rect 1932 62336 1988 62412
rect 2044 61796 2100 63982
rect 3612 63924 3668 64316
rect 3724 64260 3780 64430
rect 3724 64194 3780 64204
rect 3948 64034 4004 64046
rect 3948 63982 3950 64034
rect 4002 63982 4004 64034
rect 3612 63868 3780 63924
rect 3276 63810 3332 63822
rect 3276 63758 3278 63810
rect 3330 63758 3332 63810
rect 3276 63476 3332 63758
rect 3276 63420 3444 63476
rect 3388 63364 3444 63420
rect 3388 63308 3668 63364
rect 3276 63252 3332 63262
rect 3276 63250 3556 63252
rect 3276 63198 3278 63250
rect 3330 63198 3556 63250
rect 3276 63196 3556 63198
rect 3276 63186 3332 63196
rect 2044 61730 2100 61740
rect 2156 63026 2212 63038
rect 2156 62974 2158 63026
rect 2210 62974 2212 63026
rect 2156 62916 2212 62974
rect 1820 60386 1876 60396
rect 2044 61458 2100 61470
rect 2044 61406 2046 61458
rect 2098 61406 2100 61458
rect 2044 61348 2100 61406
rect 2044 59780 2100 61292
rect 2156 61124 2212 62860
rect 3276 62244 3332 62254
rect 3276 62242 3444 62244
rect 3276 62190 3278 62242
rect 3330 62190 3444 62242
rect 3276 62188 3444 62190
rect 3276 62178 3332 62188
rect 3276 61684 3332 61694
rect 3276 61590 3332 61628
rect 3388 61124 3444 62188
rect 3500 62132 3556 63196
rect 3500 62066 3556 62076
rect 3612 61460 3668 63308
rect 3724 63028 3780 63868
rect 3948 63812 4004 63982
rect 3836 63252 3892 63262
rect 3948 63252 4004 63756
rect 3836 63250 4004 63252
rect 3836 63198 3838 63250
rect 3890 63198 4004 63250
rect 3836 63196 4004 63198
rect 3836 63186 3892 63196
rect 3724 62962 3780 62972
rect 3724 62468 3780 62478
rect 3724 62374 3780 62412
rect 3612 61394 3668 61404
rect 3724 61348 3780 61358
rect 3724 61254 3780 61292
rect 3388 61068 3892 61124
rect 2156 61058 2212 61068
rect 2044 59714 2100 59724
rect 2156 60898 2212 60910
rect 2156 60846 2158 60898
rect 2210 60846 2212 60898
rect 2156 60676 2212 60846
rect 1932 59332 1988 59342
rect 1820 59276 1932 59332
rect 1820 57092 1876 59276
rect 1932 59200 1988 59276
rect 2156 58436 2212 60620
rect 3276 60676 3332 60686
rect 3724 60676 3780 60686
rect 3276 60674 3668 60676
rect 3276 60622 3278 60674
rect 3330 60622 3668 60674
rect 3276 60620 3668 60622
rect 3276 60610 3332 60620
rect 3276 60114 3332 60126
rect 3276 60062 3278 60114
rect 3330 60062 3332 60114
rect 2156 58370 2212 58380
rect 2268 59890 2324 59902
rect 2268 59838 2270 59890
rect 2322 59838 2324 59890
rect 2268 59780 2324 59838
rect 3276 59780 3332 60062
rect 3276 59724 3556 59780
rect 2044 58322 2100 58334
rect 2044 58270 2046 58322
rect 2098 58270 2100 58322
rect 2044 58212 2100 58270
rect 1820 57026 1876 57036
rect 1932 57762 1988 57774
rect 1932 57710 1934 57762
rect 1986 57710 1988 57762
rect 1932 57540 1988 57710
rect 1820 56196 1876 56206
rect 1820 54404 1876 56140
rect 1932 55748 1988 57484
rect 2044 56420 2100 58156
rect 2268 57764 2324 59724
rect 3276 59108 3332 59118
rect 3276 59106 3444 59108
rect 3276 59054 3278 59106
rect 3330 59054 3444 59106
rect 3276 59052 3444 59054
rect 3276 59042 3332 59052
rect 3276 58546 3332 58558
rect 3276 58494 3278 58546
rect 3330 58494 3332 58546
rect 3276 58212 3332 58494
rect 3388 58324 3444 59052
rect 3500 58772 3556 59724
rect 3500 58706 3556 58716
rect 3612 58660 3668 60620
rect 3724 60582 3780 60620
rect 3836 60004 3892 61068
rect 3836 59938 3892 59948
rect 3724 59778 3780 59790
rect 3724 59726 3726 59778
rect 3778 59726 3780 59778
rect 3724 59332 3780 59726
rect 3724 59266 3780 59276
rect 3948 59330 4004 59342
rect 3948 59278 3950 59330
rect 4002 59278 4004 59330
rect 3612 58594 3668 58604
rect 3948 59108 4004 59278
rect 3836 58548 3892 58558
rect 3948 58548 4004 59052
rect 3836 58546 4004 58548
rect 3836 58494 3838 58546
rect 3890 58494 4004 58546
rect 3836 58492 4004 58494
rect 3836 58482 3892 58492
rect 3388 58268 3892 58324
rect 3276 58156 3668 58212
rect 2268 57698 2324 57708
rect 3164 57538 3220 57550
rect 3164 57486 3166 57538
rect 3218 57486 3220 57538
rect 2268 56756 2324 56766
rect 2044 56354 2100 56364
rect 2156 56700 2268 56756
rect 1932 55682 1988 55692
rect 2156 55524 2212 56700
rect 2268 56662 2324 56700
rect 3164 56308 3220 57486
rect 3612 57092 3668 58156
rect 3724 57540 3780 57550
rect 3724 57446 3780 57484
rect 3724 57092 3780 57102
rect 3612 57036 3724 57092
rect 3724 57026 3780 57036
rect 3276 56980 3332 56990
rect 3276 56978 3444 56980
rect 3276 56926 3278 56978
rect 3330 56926 3444 56978
rect 3276 56924 3444 56926
rect 3276 56914 3332 56924
rect 3388 56756 3444 56924
rect 3836 56868 3892 58268
rect 3836 56802 3892 56812
rect 3724 56756 3780 56766
rect 3388 56700 3668 56756
rect 3164 56252 3444 56308
rect 2268 56196 2324 56206
rect 3388 56196 3444 56252
rect 3388 56140 3556 56196
rect 2268 56102 2324 56140
rect 3276 55972 3332 55982
rect 3276 55970 3444 55972
rect 3276 55918 3278 55970
rect 3330 55918 3444 55970
rect 3276 55916 3444 55918
rect 3276 55906 3332 55916
rect 2156 55458 2212 55468
rect 3276 55412 3332 55422
rect 3276 55318 3332 55356
rect 1820 54338 1876 54348
rect 2044 55186 2100 55198
rect 2044 55134 2046 55186
rect 2098 55134 2100 55186
rect 2044 55076 2100 55134
rect 2044 53844 2100 55020
rect 2044 53778 2100 53788
rect 2156 54740 2212 54750
rect 2156 54626 2212 54684
rect 2156 54574 2158 54626
rect 2210 54574 2212 54626
rect 2044 53618 2100 53630
rect 2044 53566 2046 53618
rect 2098 53566 2100 53618
rect 2044 53508 2100 53566
rect 1932 53058 1988 53070
rect 1932 53006 1934 53058
rect 1986 53006 1988 53058
rect 1932 52836 1988 53006
rect 1932 51716 1988 52780
rect 2044 52388 2100 53452
rect 2156 53060 2212 54574
rect 3388 54628 3444 55916
rect 3500 55188 3556 56140
rect 3500 55122 3556 55132
rect 3388 54562 3444 54572
rect 3612 54516 3668 56700
rect 3724 56662 3780 56700
rect 3724 56196 3780 56206
rect 3724 56102 3780 56140
rect 4060 55468 4116 67172
rect 4284 65380 4340 68014
rect 64876 67956 64932 67966
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 63532 67060 63588 67070
rect 63532 66966 63588 67004
rect 63420 66948 63476 66958
rect 63420 66854 63476 66892
rect 63980 66948 64036 66958
rect 63980 66854 64036 66892
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 64876 66388 64932 67900
rect 66780 67956 66836 69356
rect 67116 68516 67172 68526
rect 67116 68422 67172 68460
rect 67676 68516 67732 68526
rect 67676 68422 67732 68460
rect 67788 68404 67844 68414
rect 68460 68404 68516 73052
rect 68796 73108 68852 73118
rect 68796 73106 68964 73108
rect 68796 73054 68798 73106
rect 68850 73054 68964 73106
rect 68796 73052 68964 73054
rect 68796 73042 68852 73052
rect 68908 72436 68964 73052
rect 69356 72436 69412 72446
rect 68908 72380 69356 72436
rect 68572 69524 68628 69534
rect 68572 68738 68628 69468
rect 68572 68686 68574 68738
rect 68626 68686 68628 68738
rect 68572 68674 68628 68686
rect 67788 68402 68404 68404
rect 67788 68350 67790 68402
rect 67842 68350 68404 68402
rect 67788 68348 68404 68350
rect 68460 68348 68628 68404
rect 67788 68338 67844 68348
rect 67900 68180 67956 68190
rect 66780 67954 67060 67956
rect 66780 67902 66782 67954
rect 66834 67902 67060 67954
rect 66780 67900 67060 67902
rect 66780 67890 66836 67900
rect 66332 67620 66388 67630
rect 66332 67526 66388 67564
rect 67004 67170 67060 67900
rect 67900 67954 67956 68124
rect 67900 67902 67902 67954
rect 67954 67902 67956 67954
rect 67900 67890 67956 67902
rect 67228 67730 67284 67742
rect 67228 67678 67230 67730
rect 67282 67678 67284 67730
rect 67228 67620 67284 67678
rect 67228 67554 67284 67564
rect 67340 67618 67396 67630
rect 68012 67620 68068 67630
rect 67340 67566 67342 67618
rect 67394 67566 67396 67618
rect 67004 67118 67006 67170
rect 67058 67118 67060 67170
rect 67004 67106 67060 67118
rect 65660 67060 65716 67070
rect 64540 66386 64932 66388
rect 64540 66334 64878 66386
rect 64930 66334 64932 66386
rect 64540 66332 64932 66334
rect 63308 66164 63364 66174
rect 63308 66070 63364 66108
rect 63868 66164 63924 66174
rect 63868 66070 63924 66108
rect 63420 66052 63476 66062
rect 63420 65958 63476 65996
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 62076 65604 62132 65614
rect 4284 65314 4340 65324
rect 4956 65492 5012 65502
rect 4284 65156 4340 65166
rect 4172 64708 4228 64718
rect 4172 64614 4228 64652
rect 4172 62916 4228 62926
rect 4172 62822 4228 62860
rect 4284 62244 4340 65100
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 4956 63924 5012 65436
rect 62076 65490 62132 65548
rect 64540 65602 64596 66332
rect 64876 66322 64932 66332
rect 65548 67058 65716 67060
rect 65548 67006 65662 67058
rect 65714 67006 65716 67058
rect 65548 67004 65716 67006
rect 65548 66050 65604 67004
rect 65660 66994 65716 67004
rect 65884 67060 65940 67070
rect 65884 66966 65940 67004
rect 65772 66946 65828 66958
rect 65772 66894 65774 66946
rect 65826 66894 65828 66946
rect 65772 66276 65828 66894
rect 66108 66946 66164 66958
rect 66108 66894 66110 66946
rect 66162 66894 66164 66946
rect 66108 66836 66164 66894
rect 66108 66770 66164 66780
rect 66332 66836 66388 66846
rect 66892 66836 66948 66846
rect 66332 66834 66948 66836
rect 66332 66782 66334 66834
rect 66386 66782 66894 66834
rect 66946 66782 66948 66834
rect 66332 66780 66948 66782
rect 66332 66770 66388 66780
rect 66892 66770 66948 66780
rect 67340 66834 67396 67566
rect 67788 67618 68068 67620
rect 67788 67566 68014 67618
rect 68066 67566 68068 67618
rect 67788 67564 68068 67566
rect 67340 66782 67342 66834
rect 67394 66782 67396 66834
rect 67340 66770 67396 66782
rect 67452 67172 67508 67182
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 65772 66210 65828 66220
rect 65884 66500 65940 66510
rect 65884 66274 65940 66444
rect 66892 66388 66948 66398
rect 66892 66294 66948 66332
rect 67452 66388 67508 67116
rect 67676 67060 67732 67070
rect 67452 66322 67508 66332
rect 67564 66948 67620 66958
rect 65884 66222 65886 66274
rect 65938 66222 65940 66274
rect 65548 65998 65550 66050
rect 65602 65998 65604 66050
rect 65548 65716 65604 65998
rect 64540 65550 64542 65602
rect 64594 65550 64596 65602
rect 64540 65538 64596 65550
rect 65436 65660 65604 65716
rect 65660 66050 65716 66062
rect 65660 65998 65662 66050
rect 65714 65998 65716 66050
rect 62076 65438 62078 65490
rect 62130 65438 62132 65490
rect 62076 65426 62132 65438
rect 65436 65492 65492 65660
rect 65660 65604 65716 65998
rect 65772 66052 65828 66062
rect 65772 65958 65828 65996
rect 65884 65828 65940 66222
rect 66220 66276 66276 66286
rect 66780 66276 66836 66286
rect 66220 66274 66836 66276
rect 66220 66222 66222 66274
rect 66274 66222 66782 66274
rect 66834 66222 66836 66274
rect 66220 66220 66836 66222
rect 66220 66210 66276 66220
rect 66780 66210 66836 66220
rect 67004 66276 67060 66286
rect 65436 65426 65492 65436
rect 65548 65548 65716 65604
rect 65772 65772 65940 65828
rect 61964 65380 62020 65390
rect 61964 65286 62020 65324
rect 62524 65380 62580 65390
rect 62524 65286 62580 65324
rect 64652 65268 64708 65278
rect 65436 65268 65492 65278
rect 64652 65266 65492 65268
rect 64652 65214 64654 65266
rect 64706 65214 65438 65266
rect 65490 65214 65492 65266
rect 64652 65212 65492 65214
rect 64652 65202 64708 65212
rect 65436 65202 65492 65212
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 65436 64932 65492 64942
rect 65548 64932 65604 65548
rect 65772 65490 65828 65772
rect 65884 65604 65940 65614
rect 65884 65510 65940 65548
rect 65772 65438 65774 65490
rect 65826 65438 65828 65490
rect 65772 64932 65828 65438
rect 66108 65492 66164 65502
rect 66108 65398 66164 65436
rect 66668 65492 66724 65502
rect 65996 65378 66052 65390
rect 65996 65326 65998 65378
rect 66050 65326 66052 65378
rect 65996 65268 66052 65326
rect 65996 65212 66612 65268
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 66444 65044 66500 65054
rect 65548 64876 65716 64932
rect 64652 64820 64708 64830
rect 63756 64708 63812 64718
rect 63756 64614 63812 64652
rect 64316 64708 64372 64718
rect 64316 64614 64372 64652
rect 60732 64596 60788 64606
rect 60732 64502 60788 64540
rect 61740 64596 61796 64606
rect 61740 64502 61796 64540
rect 61852 64484 61908 64494
rect 61852 64390 61908 64428
rect 62300 64482 62356 64494
rect 64204 64484 64260 64494
rect 62300 64430 62302 64482
rect 62354 64430 62356 64482
rect 61740 64372 61796 64382
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 4956 63858 5012 63868
rect 59052 64148 59108 64158
rect 5292 63812 5348 63822
rect 5292 63718 5348 63756
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 4284 62178 4340 62188
rect 4844 62132 4900 62142
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 4844 60900 4900 62076
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 58492 61684 58548 61694
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 58492 61012 58548 61628
rect 59052 61346 59108 64092
rect 61180 64036 61236 64046
rect 61180 63942 61236 63980
rect 61068 63924 61124 63934
rect 61068 63830 61124 63868
rect 61628 63924 61684 63934
rect 61628 63830 61684 63868
rect 59276 63812 59332 63822
rect 59276 63252 59332 63756
rect 59276 63120 59332 63196
rect 59836 63252 59892 63262
rect 59836 63158 59892 63196
rect 61404 63028 61460 63038
rect 61404 62934 61460 62972
rect 59388 62916 59444 62926
rect 59388 62822 59444 62860
rect 61516 62914 61572 62926
rect 61516 62862 61518 62914
rect 61570 62862 61572 62914
rect 61516 62580 61572 62862
rect 61516 62514 61572 62524
rect 61628 62468 61684 62478
rect 61740 62468 61796 64316
rect 62300 64148 62356 64430
rect 62300 63924 62356 64092
rect 63868 64482 64260 64484
rect 63868 64430 64206 64482
rect 64258 64430 64260 64482
rect 63868 64428 64260 64430
rect 62300 63830 62356 63868
rect 62524 64034 62580 64046
rect 62524 63982 62526 64034
rect 62578 63982 62580 64034
rect 62524 63812 62580 63982
rect 63532 64036 63588 64046
rect 63532 63942 63588 63980
rect 61964 63028 62020 63038
rect 61964 62934 62020 62972
rect 61628 62466 61796 62468
rect 61628 62414 61630 62466
rect 61682 62414 61796 62466
rect 61628 62412 61796 62414
rect 59724 62356 59780 62366
rect 59724 62262 59780 62300
rect 61180 62356 61236 62366
rect 61628 62356 61684 62412
rect 61180 62354 61684 62356
rect 61180 62302 61182 62354
rect 61234 62302 61684 62354
rect 61180 62300 61684 62302
rect 62524 62354 62580 63756
rect 63308 63922 63364 63934
rect 63308 63870 63310 63922
rect 63362 63870 63364 63922
rect 63196 63140 63252 63150
rect 63308 63140 63364 63870
rect 62972 63138 63364 63140
rect 62972 63086 63198 63138
rect 63250 63086 63364 63138
rect 62972 63084 63364 63086
rect 63420 63810 63476 63822
rect 63420 63758 63422 63810
rect 63474 63758 63476 63810
rect 63420 63140 63476 63758
rect 63756 63812 63812 63822
rect 63644 63252 63700 63262
rect 63756 63252 63812 63756
rect 63868 63362 63924 64428
rect 64204 64418 64260 64428
rect 64652 64036 64708 64764
rect 65436 64706 65492 64876
rect 65436 64654 65438 64706
rect 65490 64654 65492 64706
rect 65100 64482 65156 64494
rect 65100 64430 65102 64482
rect 65154 64430 65156 64482
rect 65100 64260 65156 64430
rect 65100 64194 65156 64204
rect 65212 64482 65268 64494
rect 65212 64430 65214 64482
rect 65266 64430 65268 64482
rect 64652 64034 65044 64036
rect 64652 63982 64654 64034
rect 64706 63982 65044 64034
rect 64652 63980 65044 63982
rect 64652 63970 64708 63980
rect 63980 63700 64036 63710
rect 64540 63700 64596 63710
rect 63980 63698 64596 63700
rect 63980 63646 63982 63698
rect 64034 63646 64542 63698
rect 64594 63646 64596 63698
rect 63980 63644 64596 63646
rect 63980 63634 64036 63644
rect 64540 63634 64596 63644
rect 63868 63310 63870 63362
rect 63922 63310 63924 63362
rect 63868 63298 63924 63310
rect 63644 63250 63812 63252
rect 63644 63198 63646 63250
rect 63698 63198 63812 63250
rect 63644 63196 63812 63198
rect 63644 63186 63700 63196
rect 63756 63140 63812 63196
rect 64988 63250 65044 63980
rect 64988 63198 64990 63250
rect 65042 63198 65044 63250
rect 64988 63186 65044 63198
rect 63420 63084 63588 63140
rect 63756 63084 64148 63140
rect 62748 62580 62804 62590
rect 62748 62486 62804 62524
rect 62972 62578 63028 63084
rect 62972 62526 62974 62578
rect 63026 62526 63028 62578
rect 62972 62514 63028 62526
rect 63196 62580 63252 63084
rect 62524 62302 62526 62354
rect 62578 62302 62580 62354
rect 61180 62290 61236 62300
rect 62524 62290 62580 62302
rect 59612 62244 59668 62254
rect 59612 62150 59668 62188
rect 60172 62244 60228 62254
rect 60172 62150 60228 62188
rect 61740 62244 61796 62254
rect 61740 62150 61796 62188
rect 62300 62244 62356 62282
rect 62300 62178 62356 62188
rect 62860 62242 62916 62254
rect 62860 62190 62862 62242
rect 62914 62190 62916 62242
rect 60284 61458 60340 61470
rect 60284 61406 60286 61458
rect 60338 61406 60340 61458
rect 59052 61294 59054 61346
rect 59106 61294 59108 61346
rect 58492 61010 58884 61012
rect 58492 60958 58494 61010
rect 58546 60958 58884 61010
rect 58492 60956 58884 60958
rect 58492 60946 58548 60956
rect 4844 60834 4900 60844
rect 57596 60788 57652 60798
rect 57596 60694 57652 60732
rect 57484 60676 57540 60686
rect 57484 60582 57540 60620
rect 58044 60676 58100 60686
rect 58044 60582 58100 60620
rect 57148 60564 57204 60574
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 56812 59890 56868 59902
rect 56812 59838 56814 59890
rect 56866 59838 56868 59890
rect 4172 59780 4228 59790
rect 4172 59686 4228 59724
rect 56364 59780 56420 59790
rect 56812 59780 56868 59838
rect 57148 59890 57204 60508
rect 58828 60114 58884 60956
rect 59052 60564 59108 61294
rect 59836 61348 59892 61358
rect 59836 61254 59892 61292
rect 60284 61348 60340 61406
rect 61516 61458 61572 61470
rect 61516 61406 61518 61458
rect 61570 61406 61572 61458
rect 60284 61282 60340 61292
rect 60396 61346 60452 61358
rect 60396 61294 60398 61346
rect 60450 61294 60452 61346
rect 60396 61012 60452 61294
rect 61516 61348 61572 61406
rect 61516 61282 61572 61292
rect 61628 61348 61684 61358
rect 62188 61348 62244 61358
rect 61628 61346 62020 61348
rect 61628 61294 61630 61346
rect 61682 61294 62020 61346
rect 61628 61292 62020 61294
rect 61628 61282 61684 61292
rect 60396 60946 60452 60956
rect 59724 60898 59780 60910
rect 59724 60846 59726 60898
rect 59778 60846 59780 60898
rect 59052 60498 59108 60508
rect 59388 60786 59444 60798
rect 59388 60734 59390 60786
rect 59442 60734 59444 60786
rect 59388 60564 59444 60734
rect 59724 60676 59780 60846
rect 60732 60900 60788 60910
rect 60732 60806 60788 60844
rect 61068 60900 61124 60910
rect 60956 60788 61012 60798
rect 60956 60694 61012 60732
rect 59724 60610 59780 60620
rect 60396 60676 60452 60686
rect 59388 60498 59444 60508
rect 58828 60062 58830 60114
rect 58882 60062 58884 60114
rect 58828 60050 58884 60062
rect 59948 60116 60004 60126
rect 57148 59838 57150 59890
rect 57202 59838 57204 59890
rect 57148 59826 57204 59838
rect 57820 60004 57876 60014
rect 56364 59778 56868 59780
rect 56364 59726 56366 59778
rect 56418 59726 56868 59778
rect 56364 59724 56868 59726
rect 56364 59668 56420 59724
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 55804 59612 56420 59668
rect 5292 59106 5348 59118
rect 5292 59054 5294 59106
rect 5346 59054 5348 59106
rect 4476 58828 4740 58838
rect 4284 58772 4340 58782
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 4172 58212 4228 58222
rect 4172 58118 4228 58156
rect 4284 57652 4340 58716
rect 4284 57586 4340 57596
rect 4956 58660 5012 58670
rect 4956 57540 5012 58604
rect 5292 58212 5348 59054
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 5292 58146 5348 58156
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 54572 57652 54628 57662
rect 54572 57558 54628 57596
rect 55132 57652 55188 57662
rect 55132 57558 55188 57596
rect 4956 57474 5012 57484
rect 55244 57426 55300 57438
rect 55244 57374 55246 57426
rect 55298 57374 55300 57426
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 4620 57092 4676 57102
rect 4620 55972 4676 57036
rect 55244 56868 55300 57374
rect 55244 56802 55300 56812
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 53228 56084 53284 56094
rect 53228 55990 53284 56028
rect 55356 56082 55412 56094
rect 55356 56030 55358 56082
rect 55410 56030 55412 56082
rect 4620 55906 4676 55916
rect 53116 55972 53172 55982
rect 53116 55878 53172 55916
rect 53676 55972 53732 55982
rect 54796 55972 54852 55982
rect 53676 55878 53732 55916
rect 54572 55970 54852 55972
rect 54572 55918 54798 55970
rect 54850 55918 54852 55970
rect 54572 55916 54852 55918
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 3948 55412 4004 55422
rect 4060 55412 5012 55468
rect 3724 55076 3780 55086
rect 3724 54982 3780 55020
rect 3724 54740 3780 54750
rect 3724 54646 3780 54684
rect 3612 54450 3668 54460
rect 3276 54404 3332 54414
rect 3276 54402 3556 54404
rect 3276 54350 3278 54402
rect 3330 54350 3556 54402
rect 3276 54348 3556 54350
rect 3276 54338 3332 54348
rect 3276 53844 3332 53854
rect 3276 53842 3444 53844
rect 3276 53790 3278 53842
rect 3330 53790 3444 53842
rect 3276 53788 3444 53790
rect 3276 53778 3332 53788
rect 3388 53732 3444 53788
rect 3388 53666 3444 53676
rect 2156 52994 2212 53004
rect 3500 52948 3556 54348
rect 3724 53508 3780 53518
rect 3724 53414 3780 53452
rect 3500 52882 3556 52892
rect 3276 52836 3332 52846
rect 3724 52836 3780 52846
rect 3276 52834 3444 52836
rect 3276 52782 3278 52834
rect 3330 52782 3444 52834
rect 3276 52780 3444 52782
rect 3276 52770 3332 52780
rect 3388 52724 3444 52780
rect 3724 52742 3780 52780
rect 3948 52836 4004 55356
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 3948 52770 4004 52780
rect 3388 52658 3444 52668
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 2044 52322 2100 52332
rect 3276 52276 3332 52286
rect 3276 52274 3444 52276
rect 3276 52222 3278 52274
rect 3330 52222 3444 52274
rect 3276 52220 3444 52222
rect 3276 52210 3332 52220
rect 1932 51650 1988 51660
rect 2044 52050 2100 52062
rect 2044 51998 2046 52050
rect 2098 51998 2100 52050
rect 2044 51940 2100 51998
rect 3388 52052 3444 52220
rect 3388 51986 3444 51996
rect 3724 52162 3780 52174
rect 3724 52110 3726 52162
rect 3778 52110 3780 52162
rect 2044 51044 2100 51884
rect 3724 51940 3780 52110
rect 3724 51874 3780 51884
rect 2044 50978 2100 50988
rect 2156 51490 2212 51502
rect 2156 51438 2158 51490
rect 2210 51438 2212 51490
rect 2156 51268 2212 51438
rect 1932 50596 1988 50606
rect 1932 50482 1988 50540
rect 1932 50430 1934 50482
rect 1986 50430 1988 50482
rect 1932 49812 1988 50430
rect 2156 50484 2212 51212
rect 3276 51268 3332 51278
rect 3724 51268 3780 51278
rect 3276 51266 3668 51268
rect 3276 51214 3278 51266
rect 3330 51214 3668 51266
rect 3276 51212 3668 51214
rect 3276 51202 3332 51212
rect 3276 50708 3332 50718
rect 3276 50706 3556 50708
rect 3276 50654 3278 50706
rect 3330 50654 3556 50706
rect 3276 50652 3556 50654
rect 3276 50642 3332 50652
rect 2156 50418 2212 50428
rect 1932 49746 1988 49756
rect 2044 49922 2100 49934
rect 2044 49870 2046 49922
rect 2098 49870 2100 49922
rect 2044 49700 2100 49870
rect 3500 49812 3556 50652
rect 3612 49924 3668 51212
rect 3724 51174 3780 51212
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4956 50708 5012 55412
rect 54460 55412 54516 55422
rect 52332 55300 52388 55310
rect 50652 55186 50708 55198
rect 50652 55134 50654 55186
rect 50706 55134 50708 55186
rect 50652 55076 50708 55134
rect 50764 55188 50820 55198
rect 50764 55094 50820 55132
rect 50652 55010 50708 55020
rect 51212 55076 51268 55086
rect 51212 54982 51268 55020
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 52220 54628 52276 54638
rect 52220 54534 52276 54572
rect 51548 54516 51604 54526
rect 51548 54422 51604 54460
rect 52108 54516 52164 54526
rect 52108 54422 52164 54460
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 48188 53732 48244 53742
rect 52220 53732 52276 53742
rect 52332 53732 52388 55244
rect 54236 55300 54292 55310
rect 54236 55206 54292 55244
rect 54460 55186 54516 55356
rect 54572 55300 54628 55916
rect 54796 55906 54852 55916
rect 55356 55636 55412 56030
rect 55580 56084 55636 56094
rect 55580 55990 55636 56028
rect 55692 56082 55748 56094
rect 55692 56030 55694 56082
rect 55746 56030 55748 56082
rect 54572 55234 54628 55244
rect 54684 55580 55412 55636
rect 54460 55134 54462 55186
rect 54514 55134 54516 55186
rect 53676 55076 53732 55086
rect 53676 55074 53844 55076
rect 53676 55022 53678 55074
rect 53730 55022 53844 55074
rect 53676 55020 53844 55022
rect 53676 55010 53732 55020
rect 53788 54740 53844 55020
rect 53900 54740 53956 54750
rect 53788 54684 53900 54740
rect 53900 54626 53956 54684
rect 53900 54574 53902 54626
rect 53954 54574 53956 54626
rect 53900 54562 53956 54574
rect 52780 54404 52836 54414
rect 52780 54310 52836 54348
rect 53340 54404 53396 54414
rect 53340 54310 53396 54348
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 47740 52948 47796 52958
rect 47740 52854 47796 52892
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 48188 52276 48244 53676
rect 51772 53730 52388 53732
rect 51772 53678 52222 53730
rect 52274 53678 52388 53730
rect 51772 53676 52388 53678
rect 52892 54290 52948 54302
rect 52892 54238 52894 54290
rect 52946 54238 52948 54290
rect 52892 53732 52948 54238
rect 54012 54292 54068 54302
rect 54012 54290 54292 54292
rect 54012 54238 54014 54290
rect 54066 54238 54292 54290
rect 54012 54236 54292 54238
rect 54012 54226 54068 54236
rect 54236 53954 54292 54236
rect 54236 53902 54238 53954
rect 54290 53902 54292 53954
rect 54236 53890 54292 53902
rect 54460 53842 54516 55134
rect 54684 54514 54740 55580
rect 55020 55412 55076 55422
rect 54908 54628 54964 54638
rect 54908 54534 54964 54572
rect 54684 54462 54686 54514
rect 54738 54462 54740 54514
rect 54684 53956 54740 54462
rect 55020 54514 55076 55356
rect 55244 55300 55300 55310
rect 55356 55300 55412 55580
rect 55468 55970 55524 55982
rect 55468 55918 55470 55970
rect 55522 55918 55524 55970
rect 55468 55468 55524 55918
rect 55468 55412 55636 55468
rect 55244 55298 55412 55300
rect 55244 55246 55246 55298
rect 55298 55246 55412 55298
rect 55244 55244 55412 55246
rect 55244 55234 55300 55244
rect 55468 55188 55524 55198
rect 55468 55094 55524 55132
rect 55356 55076 55412 55086
rect 55020 54462 55022 54514
rect 55074 54462 55076 54514
rect 55020 54450 55076 54462
rect 55132 55074 55412 55076
rect 55132 55022 55358 55074
rect 55410 55022 55412 55074
rect 55132 55020 55412 55022
rect 54796 54404 54852 54414
rect 54796 54310 54852 54348
rect 54684 53890 54740 53900
rect 54460 53790 54462 53842
rect 54514 53790 54516 53842
rect 54460 53778 54516 53790
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 48300 52948 48356 52958
rect 48300 52854 48356 52892
rect 50540 52948 50596 52958
rect 51772 52948 51828 53676
rect 52220 53666 52276 53676
rect 52892 53666 52948 53676
rect 54684 53732 54740 53742
rect 54684 53638 54740 53676
rect 53564 53620 53620 53630
rect 53564 53618 53732 53620
rect 53564 53566 53566 53618
rect 53618 53566 53732 53618
rect 53564 53564 53732 53566
rect 53564 53554 53620 53564
rect 53452 53506 53508 53518
rect 53452 53454 53454 53506
rect 53506 53454 53508 53506
rect 51996 53060 52052 53070
rect 51996 53058 52388 53060
rect 51996 53006 51998 53058
rect 52050 53006 52388 53058
rect 51996 53004 52388 53006
rect 51996 52994 52052 53004
rect 50540 52854 50596 52892
rect 51324 52946 51828 52948
rect 51324 52894 51774 52946
rect 51826 52894 51828 52946
rect 51324 52892 51828 52894
rect 50428 52836 50484 52846
rect 50428 52742 50484 52780
rect 50988 52836 51044 52846
rect 50988 52742 51044 52780
rect 48412 52724 48468 52734
rect 49532 52724 49588 52734
rect 48412 52722 48580 52724
rect 48412 52670 48414 52722
rect 48466 52670 48580 52722
rect 48412 52668 48580 52670
rect 48412 52658 48468 52668
rect 48300 52276 48356 52286
rect 48188 52220 48300 52276
rect 48300 52144 48356 52220
rect 48412 51940 48468 51950
rect 48412 51846 48468 51884
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 48524 51492 48580 52668
rect 48860 52276 48916 52286
rect 48860 52182 48916 52220
rect 49532 52274 49588 52668
rect 51324 52276 51380 52892
rect 51772 52882 51828 52892
rect 49532 52222 49534 52274
rect 49586 52222 49588 52274
rect 48524 51426 48580 51436
rect 48972 52052 49028 52062
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 4956 50642 5012 50652
rect 48972 50708 49028 51996
rect 49532 51602 49588 52222
rect 50876 52274 51380 52276
rect 50876 52222 51326 52274
rect 51378 52222 51380 52274
rect 50876 52220 51380 52222
rect 50876 52162 50932 52220
rect 51324 52210 51380 52220
rect 52332 52836 52388 53004
rect 50876 52110 50878 52162
rect 50930 52110 50932 52162
rect 50876 52098 50932 52110
rect 52332 52162 52388 52780
rect 52892 52946 52948 52958
rect 52892 52894 52894 52946
rect 52946 52894 52948 52946
rect 52668 52276 52724 52286
rect 52668 52182 52724 52220
rect 52332 52110 52334 52162
rect 52386 52110 52388 52162
rect 49532 51550 49534 51602
rect 49586 51550 49588 51602
rect 49532 51538 49588 51550
rect 49644 51938 49700 51950
rect 50540 51940 50596 51950
rect 51996 51940 52052 51950
rect 49644 51886 49646 51938
rect 49698 51886 49700 51938
rect 49644 51380 49700 51886
rect 49644 51314 49700 51324
rect 50428 51938 50596 51940
rect 50428 51886 50542 51938
rect 50594 51886 50596 51938
rect 50428 51884 50596 51886
rect 50428 50932 50484 51884
rect 50540 51874 50596 51884
rect 51884 51938 52052 51940
rect 51884 51886 51998 51938
rect 52050 51886 52052 51938
rect 51884 51884 52052 51886
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 51884 51604 51940 51884
rect 51996 51874 52052 51884
rect 52108 51938 52164 51950
rect 52108 51886 52110 51938
rect 52162 51886 52164 51938
rect 52108 51828 52164 51886
rect 52220 51940 52276 51950
rect 52220 51846 52276 51884
rect 52108 51762 52164 51772
rect 51884 51472 51940 51548
rect 52108 51490 52164 51502
rect 52108 51438 52110 51490
rect 52162 51438 52164 51490
rect 52108 51380 52164 51438
rect 52108 51314 52164 51324
rect 52332 51378 52388 52110
rect 52556 52164 52612 52174
rect 52332 51326 52334 51378
rect 52386 51326 52388 51378
rect 52332 51314 52388 51326
rect 52444 51828 52500 51838
rect 51996 51266 52052 51278
rect 51996 51214 51998 51266
rect 52050 51214 52052 51266
rect 50428 50876 50932 50932
rect 49420 50708 49476 50718
rect 48972 50706 49476 50708
rect 48972 50654 48974 50706
rect 49026 50654 49422 50706
rect 49474 50654 49476 50706
rect 48972 50652 49476 50654
rect 48972 50642 49028 50652
rect 49420 50642 49476 50652
rect 50540 50708 50596 50718
rect 50876 50708 50932 50876
rect 50540 50706 50820 50708
rect 50540 50654 50542 50706
rect 50594 50654 50820 50706
rect 50540 50652 50820 50654
rect 50540 50642 50596 50652
rect 3724 50596 3780 50606
rect 3724 50502 3780 50540
rect 49532 50484 49588 50494
rect 49532 50390 49588 50428
rect 50428 50482 50484 50494
rect 50428 50430 50430 50482
rect 50482 50430 50484 50482
rect 50428 50372 50484 50430
rect 50652 50484 50708 50494
rect 50652 50390 50708 50428
rect 50204 50316 50428 50372
rect 50764 50372 50820 50652
rect 50876 50706 51044 50708
rect 50876 50654 50878 50706
rect 50930 50654 51044 50706
rect 50876 50652 51044 50654
rect 50876 50642 50932 50652
rect 50764 50316 50932 50372
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 50204 50036 50260 50316
rect 50428 50306 50484 50316
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 49868 50034 50260 50036
rect 49868 49982 50206 50034
rect 50258 49982 50260 50034
rect 49868 49980 50260 49982
rect 3612 49858 3668 49868
rect 46732 49924 46788 49934
rect 46732 49830 46788 49868
rect 3500 49746 3556 49756
rect 46620 49812 46676 49822
rect 46620 49718 46676 49756
rect 47180 49812 47236 49822
rect 47180 49718 47236 49756
rect 49420 49812 49476 49822
rect 2044 49028 2100 49644
rect 3276 49700 3332 49710
rect 3724 49700 3780 49710
rect 3276 49698 3444 49700
rect 3276 49646 3278 49698
rect 3330 49646 3444 49698
rect 3276 49644 3444 49646
rect 3276 49634 3332 49644
rect 3388 49252 3444 49644
rect 3724 49606 3780 49644
rect 48188 49700 48244 49710
rect 48188 49606 48244 49644
rect 48748 49700 48804 49710
rect 48748 49606 48804 49644
rect 48300 49586 48356 49598
rect 48300 49534 48302 49586
rect 48354 49534 48356 49586
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 3388 49186 3444 49196
rect 48076 49252 48132 49262
rect 3276 49140 3332 49150
rect 3276 49046 3332 49084
rect 48076 49138 48132 49196
rect 48076 49086 48078 49138
rect 48130 49086 48132 49138
rect 48076 49074 48132 49086
rect 2044 48962 2100 48972
rect 1932 48914 1988 48926
rect 1932 48862 1934 48914
rect 1986 48862 1988 48914
rect 1932 48804 1988 48862
rect 1932 48356 1988 48748
rect 3836 48802 3892 48814
rect 3836 48750 3838 48802
rect 3890 48750 3892 48802
rect 3836 48356 3892 48750
rect 4172 48804 4228 48814
rect 4172 48710 4228 48748
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 1932 48290 1988 48300
rect 3052 48300 3892 48356
rect 3052 48242 3108 48300
rect 3052 48190 3054 48242
rect 3106 48190 3108 48242
rect 3052 48178 3108 48190
rect 2044 48130 2100 48142
rect 2044 48078 2046 48130
rect 2098 48078 2100 48130
rect 1932 47346 1988 47358
rect 1932 47294 1934 47346
rect 1986 47294 1988 47346
rect 1932 46340 1988 47294
rect 2044 47012 2100 48078
rect 3724 48130 3780 48142
rect 3724 48078 3726 48130
rect 3778 48078 3780 48130
rect 3724 47684 3780 48078
rect 3724 47618 3780 47628
rect 3052 47460 3108 47470
rect 3052 47458 3556 47460
rect 3052 47406 3054 47458
rect 3106 47406 3556 47458
rect 3052 47404 3556 47406
rect 3052 47394 3108 47404
rect 3500 47236 3556 47404
rect 3500 47234 3780 47236
rect 3500 47182 3502 47234
rect 3554 47182 3780 47234
rect 3500 47180 3780 47182
rect 3500 47170 3556 47180
rect 2044 46946 2100 46956
rect 3052 46676 3108 46686
rect 3052 46582 3108 46620
rect 3612 46676 3668 46686
rect 1932 46274 1988 46284
rect 2044 46562 2100 46574
rect 2044 46510 2046 46562
rect 2098 46510 2100 46562
rect 1932 45778 1988 45790
rect 1932 45726 1934 45778
rect 1986 45726 1988 45778
rect 1932 44996 1988 45726
rect 2044 45668 2100 46510
rect 3612 46562 3668 46620
rect 3612 46510 3614 46562
rect 3666 46510 3668 46562
rect 3052 45890 3108 45902
rect 3052 45838 3054 45890
rect 3106 45838 3108 45890
rect 3052 45668 3108 45838
rect 3500 45668 3556 45678
rect 3052 45666 3556 45668
rect 3052 45614 3502 45666
rect 3554 45614 3556 45666
rect 3052 45612 3556 45614
rect 2044 45602 2100 45612
rect 3500 45332 3556 45612
rect 3500 45266 3556 45276
rect 3612 45220 3668 46510
rect 3724 45668 3780 47180
rect 3836 46788 3892 48300
rect 4844 48242 4900 48254
rect 4844 48190 4846 48242
rect 4898 48190 4900 48242
rect 4844 48132 4900 48190
rect 48300 48244 48356 49534
rect 48412 49252 48468 49262
rect 48412 48354 48468 49196
rect 49420 49138 49476 49756
rect 49420 49086 49422 49138
rect 49474 49086 49476 49138
rect 49420 49074 49476 49086
rect 49196 49028 49252 49038
rect 49868 49028 49924 49980
rect 50204 49970 50260 49980
rect 50428 49924 50484 49934
rect 50428 49830 50484 49868
rect 49196 49026 49364 49028
rect 49196 48974 49198 49026
rect 49250 48974 49364 49026
rect 49196 48972 49364 48974
rect 49196 48962 49252 48972
rect 48524 48804 48580 48814
rect 48524 48466 48580 48748
rect 48524 48414 48526 48466
rect 48578 48414 48580 48466
rect 48524 48402 48580 48414
rect 48412 48302 48414 48354
rect 48466 48302 48468 48354
rect 48412 48290 48468 48302
rect 48300 48178 48356 48188
rect 4844 48066 4900 48076
rect 5404 48132 5460 48142
rect 5404 48038 5460 48076
rect 47068 48132 47124 48142
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 47068 47346 47124 48076
rect 47740 48130 47796 48142
rect 47740 48078 47742 48130
rect 47794 48078 47796 48130
rect 47068 47294 47070 47346
rect 47122 47294 47124 47346
rect 47068 47282 47124 47294
rect 47404 47348 47460 47358
rect 47404 47254 47460 47292
rect 47740 47348 47796 48078
rect 49308 48132 49364 48972
rect 49532 49026 49924 49028
rect 49532 48974 49870 49026
rect 49922 48974 49924 49026
rect 49532 48972 49924 48974
rect 49532 48468 49588 48972
rect 49868 48962 49924 48972
rect 50092 49812 50148 49822
rect 49644 48804 49700 48814
rect 49644 48710 49700 48748
rect 49756 48802 49812 48814
rect 49756 48750 49758 48802
rect 49810 48750 49812 48802
rect 49644 48468 49700 48478
rect 49532 48466 49700 48468
rect 49532 48414 49646 48466
rect 49698 48414 49700 48466
rect 49532 48412 49700 48414
rect 49756 48468 49812 48750
rect 49756 48412 50036 48468
rect 49644 48402 49700 48412
rect 49868 48244 49924 48254
rect 49868 48150 49924 48188
rect 49308 48076 49588 48132
rect 49532 47682 49588 48076
rect 49532 47630 49534 47682
rect 49586 47630 49588 47682
rect 49532 47618 49588 47630
rect 49756 48130 49812 48142
rect 49756 48078 49758 48130
rect 49810 48078 49812 48130
rect 47740 47282 47796 47292
rect 48076 47348 48132 47358
rect 48076 47254 48132 47292
rect 48860 47348 48916 47358
rect 48412 47236 48468 47246
rect 48412 47142 48468 47180
rect 48860 47234 48916 47292
rect 49644 47348 49700 47358
rect 49644 47254 49700 47292
rect 48860 47182 48862 47234
rect 48914 47182 48916 47234
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 3836 46722 3892 46732
rect 46396 46788 46452 46798
rect 46396 46694 46452 46732
rect 47740 46788 47796 46798
rect 47740 46694 47796 46732
rect 45948 46676 46004 46686
rect 45948 46582 46004 46620
rect 46732 46676 46788 46686
rect 46732 46582 46788 46620
rect 47516 46676 47572 46686
rect 47516 46582 47572 46620
rect 48188 46676 48244 46686
rect 48188 46564 48244 46620
rect 48188 46562 48468 46564
rect 48188 46510 48190 46562
rect 48242 46510 48468 46562
rect 48188 46508 48468 46510
rect 48188 46498 48244 46508
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 46060 45892 46116 45902
rect 46060 45798 46116 45836
rect 46956 45892 47012 45902
rect 46956 45798 47012 45836
rect 47740 45892 47796 45902
rect 47180 45780 47236 45790
rect 47180 45686 47236 45724
rect 3724 45602 3780 45612
rect 45724 45668 45780 45678
rect 45724 45574 45780 45612
rect 47740 45668 47796 45836
rect 48188 45668 48244 45678
rect 47740 45666 48244 45668
rect 47740 45614 47742 45666
rect 47794 45614 48190 45666
rect 48242 45614 48244 45666
rect 47740 45612 48244 45614
rect 45612 45556 45668 45566
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 44380 45332 44436 45342
rect 44380 45238 44436 45276
rect 45612 45330 45668 45500
rect 45612 45278 45614 45330
rect 45666 45278 45668 45330
rect 45612 45266 45668 45278
rect 3612 45154 3668 45164
rect 46172 45220 46228 45230
rect 46172 45126 46228 45164
rect 47404 45220 47460 45230
rect 47404 45126 47460 45164
rect 3052 45106 3108 45118
rect 3052 45054 3054 45106
rect 3106 45054 3108 45106
rect 1932 44930 1988 44940
rect 2044 44994 2100 45006
rect 2044 44942 2046 44994
rect 2098 44942 2100 44994
rect 2044 44324 2100 44942
rect 3052 44996 3108 45054
rect 43932 45108 43988 45118
rect 43932 45014 43988 45052
rect 44716 45108 44772 45118
rect 44716 45014 44772 45052
rect 45388 45108 45444 45118
rect 3052 44930 3108 44940
rect 3612 44996 3668 45006
rect 3612 44902 3668 44940
rect 43708 44996 43764 45006
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 2044 44258 2100 44268
rect 3052 44322 3108 44334
rect 3052 44270 3054 44322
rect 3106 44270 3108 44322
rect 1932 44210 1988 44222
rect 1932 44158 1934 44210
rect 1986 44158 1988 44210
rect 1932 43652 1988 44158
rect 3052 44100 3108 44270
rect 43708 44210 43764 44940
rect 45388 44548 45444 45052
rect 46508 45108 46564 45118
rect 46508 45014 46564 45052
rect 47180 45108 47236 45118
rect 47180 45014 47236 45052
rect 45388 44482 45444 44492
rect 46732 44548 46788 44558
rect 43708 44158 43710 44210
rect 43762 44158 43764 44210
rect 43708 44146 43764 44158
rect 44044 44212 44100 44222
rect 44044 44118 44100 44156
rect 44604 44212 44660 44222
rect 44604 44118 44660 44156
rect 45500 44212 45556 44222
rect 45500 44118 45556 44156
rect 46396 44212 46452 44222
rect 3052 44034 3108 44044
rect 3500 44100 3556 44110
rect 3500 44006 3556 44044
rect 43036 44100 43092 44110
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 43036 43762 43092 44044
rect 45836 44100 45892 44110
rect 45836 44006 45892 44044
rect 43036 43710 43038 43762
rect 43090 43710 43092 43762
rect 43036 43698 43092 43710
rect 44492 43764 44548 43802
rect 44492 43698 44548 43708
rect 1932 43586 1988 43596
rect 3052 43538 3108 43550
rect 3052 43486 3054 43538
rect 3106 43486 3108 43538
rect 1932 43426 1988 43438
rect 1932 43374 1934 43426
rect 1986 43374 1988 43426
rect 1932 42980 1988 43374
rect 3052 43428 3108 43486
rect 42588 43540 42644 43550
rect 42588 43446 42644 43484
rect 43372 43540 43428 43550
rect 43372 43446 43428 43484
rect 44268 43540 44324 43550
rect 44268 43446 44324 43484
rect 44940 43540 44996 43550
rect 3052 43362 3108 43372
rect 3612 43428 3668 43438
rect 3612 43334 3668 43372
rect 42364 43428 42420 43438
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 1932 42914 1988 42924
rect 3052 42754 3108 42766
rect 3052 42702 3054 42754
rect 3106 42702 3108 42754
rect 1932 42642 1988 42654
rect 1932 42590 1934 42642
rect 1986 42590 1988 42642
rect 1932 42308 1988 42590
rect 3052 42644 3108 42702
rect 3052 42578 3108 42588
rect 3500 42644 3556 42654
rect 3500 42550 3556 42588
rect 41804 42644 41860 42654
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 1932 42242 1988 42252
rect 41804 42194 41860 42588
rect 42364 42642 42420 43372
rect 44940 43426 44996 43484
rect 44940 43374 44942 43426
rect 44994 43374 44996 43426
rect 43484 42754 43540 42766
rect 43484 42702 43486 42754
rect 43538 42702 43540 42754
rect 42364 42590 42366 42642
rect 42418 42590 42420 42642
rect 42364 42578 42420 42590
rect 42700 42644 42756 42654
rect 42700 42550 42756 42588
rect 43484 42644 43540 42702
rect 41916 42532 41972 42542
rect 41916 42438 41972 42476
rect 41804 42142 41806 42194
rect 41858 42142 41860 42194
rect 41804 42130 41860 42142
rect 43148 42084 43204 42094
rect 43148 41990 43204 42028
rect 3052 41970 3108 41982
rect 3052 41918 3054 41970
rect 3106 41918 3108 41970
rect 1932 41858 1988 41870
rect 1932 41806 1934 41858
rect 1986 41806 1988 41858
rect 1932 41636 1988 41806
rect 3052 41860 3108 41918
rect 42140 41970 42196 41982
rect 42140 41918 42142 41970
rect 42194 41918 42196 41970
rect 3052 41794 3108 41804
rect 3612 41860 3668 41870
rect 3612 41766 3668 41804
rect 41020 41860 41076 41870
rect 1932 41570 1988 41580
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 3052 41186 3108 41198
rect 3052 41134 3054 41186
rect 3106 41134 3108 41186
rect 1932 41074 1988 41086
rect 1932 41022 1934 41074
rect 1986 41022 1988 41074
rect 1932 40964 1988 41022
rect 1932 40898 1988 40908
rect 3052 40964 3108 41134
rect 41020 41074 41076 41804
rect 42140 41860 42196 41918
rect 42140 41794 42196 41804
rect 42924 41970 42980 41982
rect 42924 41918 42926 41970
rect 42978 41918 42980 41970
rect 42924 41860 42980 41918
rect 41020 41022 41022 41074
rect 41074 41022 41076 41074
rect 41020 41010 41076 41022
rect 41356 41074 41412 41086
rect 41356 41022 41358 41074
rect 41410 41022 41412 41074
rect 3052 40898 3108 40908
rect 3500 40964 3556 40974
rect 3500 40870 3556 40908
rect 40124 40962 40180 40974
rect 40124 40910 40126 40962
rect 40178 40910 40180 40962
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 39452 40514 39508 40526
rect 39452 40462 39454 40514
rect 39506 40462 39508 40514
rect 3052 40404 3108 40414
rect 3052 40310 3108 40348
rect 3612 40404 3668 40414
rect 3612 40310 3668 40348
rect 39452 40404 39508 40462
rect 39452 40338 39508 40348
rect 39788 40402 39844 40414
rect 39788 40350 39790 40402
rect 39842 40350 39844 40402
rect 1932 40292 1988 40302
rect 1932 40198 1988 40236
rect 39004 40290 39060 40302
rect 39004 40238 39006 40290
rect 39058 40238 39060 40290
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 1932 39620 1988 39630
rect 1932 39526 1988 39564
rect 3052 39618 3108 39630
rect 3052 39566 3054 39618
rect 3106 39566 3108 39618
rect 3052 39508 3108 39566
rect 3052 39442 3108 39452
rect 3612 39508 3668 39518
rect 3612 39414 3668 39452
rect 38892 39508 38948 39518
rect 38892 39414 38948 39452
rect 38444 39396 38500 39406
rect 38444 39302 38500 39340
rect 39004 39396 39060 40238
rect 39788 39956 39844 40350
rect 39788 39890 39844 39900
rect 40124 39956 40180 40910
rect 40348 40964 40404 40974
rect 40348 40626 40404 40908
rect 40348 40574 40350 40626
rect 40402 40574 40404 40626
rect 40348 40562 40404 40574
rect 40572 40962 40628 40974
rect 40572 40910 40574 40962
rect 40626 40910 40628 40962
rect 40572 40628 40628 40910
rect 40572 40562 40628 40572
rect 41356 40628 41412 41022
rect 42140 41074 42196 41086
rect 42140 41022 42142 41074
rect 42194 41022 42196 41074
rect 41356 40562 41412 40572
rect 41804 40628 41860 40638
rect 40684 40404 40740 40414
rect 40684 40310 40740 40348
rect 41580 40404 41636 40414
rect 40124 39890 40180 39900
rect 40684 39956 40740 39966
rect 39004 39330 39060 39340
rect 39228 39508 39284 39518
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 1932 38948 1988 38958
rect 1932 38854 1988 38892
rect 38332 38946 38388 38958
rect 38332 38894 38334 38946
rect 38386 38894 38388 38946
rect 3052 38836 3108 38846
rect 3052 38742 3108 38780
rect 3612 38836 3668 38846
rect 3612 38742 3668 38780
rect 38332 38836 38388 38894
rect 38332 38770 38388 38780
rect 38668 38836 38724 38846
rect 38668 38742 38724 38780
rect 37884 38724 37940 38734
rect 37884 38630 37940 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 1932 38276 1988 38286
rect 1932 38162 1988 38220
rect 1932 38110 1934 38162
rect 1986 38110 1988 38162
rect 1932 38098 1988 38110
rect 3052 38050 3108 38062
rect 3052 37998 3054 38050
rect 3106 37998 3108 38050
rect 3052 37828 3108 37998
rect 38892 38050 38948 38062
rect 38892 37998 38894 38050
rect 38946 37998 38948 38050
rect 37996 37940 38052 37950
rect 37996 37846 38052 37884
rect 38892 37940 38948 37998
rect 3052 37762 3108 37772
rect 3612 37828 3668 37838
rect 3612 37734 3668 37772
rect 37660 37828 37716 37838
rect 37660 37734 37716 37772
rect 19836 37660 20100 37670
rect 1932 37604 1988 37614
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 1932 37378 1988 37548
rect 1932 37326 1934 37378
rect 1986 37326 1988 37378
rect 1932 37314 1988 37326
rect 36988 37378 37044 37390
rect 36988 37326 36990 37378
rect 37042 37326 37044 37378
rect 3052 37266 3108 37278
rect 3052 37214 3054 37266
rect 3106 37214 3108 37266
rect 3052 37044 3108 37214
rect 36540 37268 36596 37278
rect 36540 37174 36596 37212
rect 3052 36978 3108 36988
rect 3612 37154 3668 37166
rect 3612 37102 3614 37154
rect 3666 37102 3668 37154
rect 3612 37044 3668 37102
rect 3612 36978 3668 36988
rect 36988 37044 37044 37326
rect 38444 37380 38500 37390
rect 38444 37286 38500 37324
rect 36988 36978 37044 36988
rect 37324 37268 37380 37278
rect 1932 36932 1988 36942
rect 1932 36594 1988 36876
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 1932 36542 1934 36594
rect 1986 36542 1988 36594
rect 1932 36530 1988 36542
rect 3052 36482 3108 36494
rect 3052 36430 3054 36482
rect 3106 36430 3108 36482
rect 1932 36260 1988 36270
rect 1932 35810 1988 36204
rect 3052 36260 3108 36430
rect 36540 36482 36596 36494
rect 36540 36430 36542 36482
rect 36594 36430 36596 36482
rect 35868 36372 35924 36382
rect 35868 36278 35924 36316
rect 36540 36372 36596 36430
rect 3052 36194 3108 36204
rect 3612 36260 3668 36270
rect 3612 36166 3668 36204
rect 35420 36258 35476 36270
rect 35420 36206 35422 36258
rect 35474 36206 35476 36258
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 1932 35758 1934 35810
rect 1986 35758 1988 35810
rect 1932 35746 1988 35758
rect 3052 35812 3108 35822
rect 3052 35698 3108 35756
rect 3052 35646 3054 35698
rect 3106 35646 3108 35698
rect 3052 35634 3108 35646
rect 3612 35812 3668 35822
rect 1932 35588 1988 35598
rect 1932 35026 1988 35532
rect 1932 34974 1934 35026
rect 1986 34974 1988 35026
rect 1932 34962 1988 34974
rect 3612 35026 3668 35756
rect 34748 35810 34804 35822
rect 34748 35758 34750 35810
rect 34802 35758 34804 35810
rect 4844 35698 4900 35710
rect 4844 35646 4846 35698
rect 4898 35646 4900 35698
rect 3612 34974 3614 35026
rect 3666 34974 3668 35026
rect 3612 34962 3668 34974
rect 3724 35586 3780 35598
rect 3724 35534 3726 35586
rect 3778 35534 3780 35586
rect 3052 34914 3108 34926
rect 3052 34862 3054 34914
rect 3106 34862 3108 34914
rect 3052 34692 3108 34862
rect 3724 34916 3780 35534
rect 4844 35588 4900 35646
rect 4844 35522 4900 35532
rect 5404 35588 5460 35598
rect 5404 35494 5460 35532
rect 34300 35588 34356 35598
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 3724 34850 3780 34860
rect 33852 34804 33908 34814
rect 33852 34710 33908 34748
rect 34300 34802 34356 35532
rect 34300 34750 34302 34802
rect 34354 34750 34356 34802
rect 34300 34738 34356 34750
rect 34636 34804 34692 34814
rect 34636 34710 34692 34748
rect 3052 34626 3108 34636
rect 4060 34692 4116 34702
rect 4060 34598 4116 34636
rect 34748 34692 34804 35758
rect 34748 34626 34804 34636
rect 34972 35700 35028 35710
rect 35420 35700 35476 36206
rect 36316 36260 36372 36270
rect 36316 36166 36372 36204
rect 35644 35812 35700 35822
rect 35644 35718 35700 35756
rect 34972 35698 35476 35700
rect 34972 35646 34974 35698
rect 35026 35646 35476 35698
rect 34972 35644 35476 35646
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 1932 34244 1988 34254
rect 1932 34150 1988 34188
rect 33740 34242 33796 34254
rect 33740 34190 33742 34242
rect 33794 34190 33796 34242
rect 3052 34130 3108 34142
rect 3052 34078 3054 34130
rect 3106 34078 3108 34130
rect 3052 34020 3108 34078
rect 3052 33954 3108 33964
rect 3612 34020 3668 34030
rect 3612 33926 3668 33964
rect 33740 34020 33796 34190
rect 34076 34132 34132 34142
rect 34076 34038 34132 34076
rect 34860 34132 34916 34142
rect 33740 33954 33796 33964
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 1932 33572 1988 33582
rect 1932 33458 1988 33516
rect 1932 33406 1934 33458
rect 1986 33406 1988 33458
rect 1932 33394 1988 33406
rect 34860 33458 34916 34076
rect 34860 33406 34862 33458
rect 34914 33406 34916 33458
rect 3052 33346 3108 33358
rect 3052 33294 3054 33346
rect 3106 33294 3108 33346
rect 3052 33236 3108 33294
rect 32508 33348 32564 33358
rect 3052 33170 3108 33180
rect 3612 33236 3668 33246
rect 3612 33142 3668 33180
rect 32508 33124 32564 33292
rect 33180 33348 33236 33358
rect 33180 33254 33236 33292
rect 34076 33348 34132 33358
rect 34132 33292 34356 33348
rect 34076 33254 34132 33292
rect 32956 33236 33012 33246
rect 32956 33142 33012 33180
rect 32396 33122 32564 33124
rect 32396 33070 32510 33122
rect 32562 33070 32564 33122
rect 32396 33068 32564 33070
rect 19836 32956 20100 32966
rect 1932 32900 1988 32910
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 1932 32674 1988 32844
rect 1932 32622 1934 32674
rect 1986 32622 1988 32674
rect 1932 32610 1988 32622
rect 32284 32674 32340 32686
rect 32284 32622 32286 32674
rect 32338 32622 32340 32674
rect 3052 32562 3108 32574
rect 3052 32510 3054 32562
rect 3106 32510 3108 32562
rect 3052 32340 3108 32510
rect 31836 32564 31892 32574
rect 3052 32274 3108 32284
rect 3612 32450 3668 32462
rect 3612 32398 3614 32450
rect 3666 32398 3668 32450
rect 3612 32340 3668 32398
rect 3612 32274 3668 32284
rect 31836 32450 31892 32508
rect 31836 32398 31838 32450
rect 31890 32398 31892 32450
rect 1932 32228 1988 32238
rect 1932 31890 1988 32172
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 1932 31838 1934 31890
rect 1986 31838 1988 31890
rect 1932 31826 1988 31838
rect 3052 31778 3108 31790
rect 3052 31726 3054 31778
rect 3106 31726 3108 31778
rect 1932 31556 1988 31566
rect 1932 31106 1988 31500
rect 3052 31556 3108 31726
rect 31164 31668 31220 31678
rect 3052 31490 3108 31500
rect 3612 31556 3668 31566
rect 3612 31462 3668 31500
rect 30716 31554 30772 31566
rect 30716 31502 30718 31554
rect 30770 31502 30772 31554
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 1932 31054 1934 31106
rect 1986 31054 1988 31106
rect 1932 31042 1988 31054
rect 3052 31108 3108 31118
rect 3052 30994 3108 31052
rect 3052 30942 3054 30994
rect 3106 30942 3108 30994
rect 3052 30930 3108 30942
rect 3612 31108 3668 31118
rect 1932 30884 1988 30894
rect 1932 30322 1988 30828
rect 1932 30270 1934 30322
rect 1986 30270 1988 30322
rect 1932 30258 1988 30270
rect 3052 30210 3108 30222
rect 3052 30158 3054 30210
rect 3106 30158 3108 30210
rect 3052 29988 3108 30158
rect 3612 30210 3668 31052
rect 30044 31106 30100 31118
rect 30044 31054 30046 31106
rect 30098 31054 30100 31106
rect 4844 30994 4900 31006
rect 4844 30942 4846 30994
rect 4898 30942 4900 30994
rect 3612 30158 3614 30210
rect 3666 30158 3668 30210
rect 3612 30146 3668 30158
rect 3724 30882 3780 30894
rect 3724 30830 3726 30882
rect 3778 30830 3780 30882
rect 3724 30212 3780 30830
rect 4844 30884 4900 30942
rect 4844 30818 4900 30828
rect 5404 30884 5460 30894
rect 5404 30790 5460 30828
rect 29372 30882 29428 30894
rect 29372 30830 29374 30882
rect 29426 30830 29428 30882
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 3724 30146 3780 30156
rect 28812 30100 28868 30110
rect 3052 29922 3108 29932
rect 4060 29988 4116 29998
rect 28812 29988 28868 30044
rect 29372 30100 29428 30830
rect 29372 30034 29428 30044
rect 29596 30884 29652 30894
rect 29596 30098 29652 30828
rect 29596 30046 29598 30098
rect 29650 30046 29652 30098
rect 29596 30034 29652 30046
rect 29932 30100 29988 30110
rect 29932 30006 29988 30044
rect 4060 29894 4116 29932
rect 28700 29986 28868 29988
rect 28700 29934 28814 29986
rect 28866 29934 28868 29986
rect 28700 29932 28868 29934
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 1932 29540 1988 29550
rect 1932 29446 1988 29484
rect 3052 29426 3108 29438
rect 3052 29374 3054 29426
rect 3106 29374 3108 29426
rect 3052 29316 3108 29374
rect 28476 29428 28532 29438
rect 28476 29334 28532 29372
rect 3052 29250 3108 29260
rect 3612 29316 3668 29326
rect 3612 29222 3668 29260
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 1932 28868 1988 28878
rect 1932 28754 1988 28812
rect 1932 28702 1934 28754
rect 1986 28702 1988 28754
rect 1932 28690 1988 28702
rect 3052 28644 3108 28654
rect 3052 28550 3108 28588
rect 3612 28644 3668 28654
rect 27804 28644 27860 28654
rect 3612 28550 3668 28588
rect 27692 28642 27860 28644
rect 27692 28590 27806 28642
rect 27858 28590 27860 28642
rect 27692 28588 27860 28590
rect 27692 28532 27748 28588
rect 27804 28578 27860 28588
rect 28252 28644 28308 28654
rect 19836 28252 20100 28262
rect 1932 28196 1988 28206
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 1932 27970 1988 28140
rect 1932 27918 1934 27970
rect 1986 27918 1988 27970
rect 1932 27906 1988 27918
rect 27580 27970 27636 27982
rect 27580 27918 27582 27970
rect 27634 27918 27636 27970
rect 3052 27858 3108 27870
rect 3052 27806 3054 27858
rect 3106 27806 3108 27858
rect 3052 27748 3108 27806
rect 27132 27860 27188 27870
rect 3052 27682 3108 27692
rect 3612 27748 3668 27758
rect 27132 27748 27188 27804
rect 3612 27654 3668 27692
rect 27020 27746 27188 27748
rect 27020 27694 27134 27746
rect 27186 27694 27188 27746
rect 27020 27692 27188 27694
rect 1932 27524 1988 27534
rect 1932 27186 1988 27468
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 1932 27134 1934 27186
rect 1986 27134 1988 27186
rect 1932 27122 1988 27134
rect 3052 27076 3108 27086
rect 3052 26982 3108 27020
rect 3612 27076 3668 27086
rect 3612 26982 3668 27020
rect 26908 27076 26964 27086
rect 26460 26964 26516 26974
rect 26460 26870 26516 26908
rect 1932 26852 1988 26862
rect 1932 26402 1988 26796
rect 26908 26850 26964 27020
rect 26908 26798 26910 26850
rect 26962 26798 26964 26850
rect 26908 26786 26964 26798
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 1932 26350 1934 26402
rect 1986 26350 1988 26402
rect 1932 26338 1988 26350
rect 26236 26402 26292 26414
rect 26236 26350 26238 26402
rect 26290 26350 26292 26402
rect 2940 26290 2996 26302
rect 2940 26238 2942 26290
rect 2994 26238 2996 26290
rect 1932 26180 1988 26190
rect 1932 25618 1988 26124
rect 1932 25566 1934 25618
rect 1986 25566 1988 25618
rect 1932 25554 1988 25566
rect 2940 25284 2996 26238
rect 4844 26290 4900 26302
rect 4844 26238 4846 26290
rect 4898 26238 4900 26290
rect 3724 26178 3780 26190
rect 3724 26126 3726 26178
rect 3778 26126 3780 26178
rect 3052 25506 3108 25518
rect 3052 25454 3054 25506
rect 3106 25454 3108 25506
rect 3052 25396 3108 25454
rect 3724 25508 3780 26126
rect 4844 26180 4900 26238
rect 25788 26292 25844 26302
rect 25788 26198 25844 26236
rect 4844 26114 4900 26124
rect 5404 26180 5460 26190
rect 5404 26086 5460 26124
rect 24332 26180 24388 26190
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 3724 25442 3780 25452
rect 3052 25330 3108 25340
rect 4060 25396 4116 25406
rect 4060 25302 4116 25340
rect 24332 25394 24388 26124
rect 25004 26178 25060 26190
rect 25004 26126 25006 26178
rect 25058 26126 25060 26178
rect 24332 25342 24334 25394
rect 24386 25342 24388 25394
rect 24332 25330 24388 25342
rect 24668 25394 24724 25406
rect 24668 25342 24670 25394
rect 24722 25342 24724 25394
rect 2940 25218 2996 25228
rect 3612 25284 3668 25294
rect 3612 25190 3668 25228
rect 24668 25172 24724 25342
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 24668 25106 24724 25116
rect 25004 25172 25060 26126
rect 25564 25508 25620 25518
rect 25564 25414 25620 25452
rect 25228 25396 25284 25406
rect 25228 25302 25284 25340
rect 26236 25284 26292 26350
rect 26572 26292 26628 26302
rect 26572 26198 26628 26236
rect 27020 25844 27076 27692
rect 27132 27682 27188 27692
rect 27580 27748 27636 27918
rect 27580 27682 27636 27692
rect 27692 27524 27748 28476
rect 28252 28530 28308 28588
rect 28252 28478 28254 28530
rect 28306 28478 28308 28530
rect 28252 28466 28308 28478
rect 28588 28532 28644 28542
rect 28588 28438 28644 28476
rect 27804 27860 27860 27870
rect 27804 27766 27860 27804
rect 28588 27860 28644 27870
rect 28588 27766 28644 27804
rect 27580 27468 27748 27524
rect 27244 26964 27300 26974
rect 27020 25778 27076 25788
rect 27132 26292 27188 26302
rect 26460 25508 26516 25518
rect 26516 25452 26628 25508
rect 26460 25376 26516 25452
rect 26236 25218 26292 25228
rect 25004 25106 25060 25116
rect 25900 25172 25956 25182
rect 19836 25050 20100 25060
rect 1932 24836 1988 24846
rect 1932 24742 1988 24780
rect 23660 24834 23716 24846
rect 23660 24782 23662 24834
rect 23714 24782 23716 24834
rect 3052 24722 3108 24734
rect 3052 24670 3054 24722
rect 3106 24670 3108 24722
rect 3052 24500 3108 24670
rect 22764 24724 22820 24734
rect 22764 24630 22820 24668
rect 23100 24724 23156 24734
rect 23100 24630 23156 24668
rect 3052 24434 3108 24444
rect 3612 24610 3668 24622
rect 3612 24558 3614 24610
rect 3666 24558 3668 24610
rect 3612 24500 3668 24558
rect 3612 24434 3668 24444
rect 23660 24500 23716 24782
rect 24892 24834 24948 24846
rect 24892 24782 24894 24834
rect 24946 24782 24948 24834
rect 23996 24724 24052 24734
rect 24556 24724 24612 24734
rect 24052 24722 24612 24724
rect 24052 24670 24558 24722
rect 24610 24670 24612 24722
rect 24052 24668 24612 24670
rect 23996 24592 24052 24668
rect 23660 24434 23716 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 1932 24164 1988 24174
rect 1932 24050 1988 24108
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23986 1988 23998
rect 3052 23938 3108 23950
rect 3052 23886 3054 23938
rect 3106 23886 3108 23938
rect 3052 23716 3108 23886
rect 23996 23826 24052 23838
rect 23996 23774 23998 23826
rect 24050 23774 24052 23826
rect 3052 23650 3108 23660
rect 3612 23716 3668 23726
rect 3612 23622 3668 23660
rect 23100 23714 23156 23726
rect 23100 23662 23102 23714
rect 23154 23662 23156 23714
rect 19836 23548 20100 23558
rect 1932 23492 1988 23502
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 1932 23266 1988 23436
rect 1932 23214 1934 23266
rect 1986 23214 1988 23266
rect 1932 23202 1988 23214
rect 22428 23266 22484 23278
rect 22428 23214 22430 23266
rect 22482 23214 22484 23266
rect 3052 23154 3108 23166
rect 3052 23102 3054 23154
rect 3106 23102 3108 23154
rect 3052 23044 3108 23102
rect 3052 22978 3108 22988
rect 3612 23044 3668 23054
rect 3612 22950 3668 22988
rect 22428 23044 22484 23214
rect 22764 23156 22820 23166
rect 22764 23062 22820 23100
rect 23100 23156 23156 23662
rect 23660 23716 23716 23726
rect 23660 23622 23716 23660
rect 23884 23268 23940 23278
rect 23884 23174 23940 23212
rect 23100 23090 23156 23100
rect 23660 23156 23716 23166
rect 23716 23100 23828 23156
rect 23660 23024 23716 23100
rect 22428 22978 22484 22988
rect 1932 22820 1988 22830
rect 1932 22482 1988 22764
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 1932 22430 1934 22482
rect 1986 22430 1988 22482
rect 1932 22418 1988 22430
rect 3052 22370 3108 22382
rect 3052 22318 3054 22370
rect 3106 22318 3108 22370
rect 1932 22148 1988 22158
rect 1932 21698 1988 22092
rect 3052 22148 3108 22318
rect 23100 22370 23156 22382
rect 23100 22318 23102 22370
rect 23154 22318 23156 22370
rect 22428 22258 22484 22270
rect 22428 22206 22430 22258
rect 22482 22206 22484 22258
rect 3052 22082 3108 22092
rect 3612 22148 3668 22158
rect 3612 22054 3668 22092
rect 22092 22148 22148 22158
rect 22092 22054 22148 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 22428 21812 22484 22206
rect 22652 21812 22708 21822
rect 22428 21756 22652 21812
rect 22652 21718 22708 21756
rect 23100 21812 23156 22318
rect 23324 22148 23380 22158
rect 23324 22054 23380 22092
rect 23772 22146 23828 23100
rect 23996 23044 24052 23774
rect 24332 23044 24388 23054
rect 23996 23042 24388 23044
rect 23996 22990 24334 23042
rect 24386 22990 24388 23042
rect 23996 22988 24388 22990
rect 24332 22932 24388 22988
rect 24332 22866 24388 22876
rect 24332 22148 24388 22158
rect 23772 22094 23774 22146
rect 23826 22094 23828 22146
rect 23100 21746 23156 21756
rect 1932 21646 1934 21698
rect 1986 21646 1988 21698
rect 1932 21634 1988 21646
rect 21756 21698 21812 21710
rect 21756 21646 21758 21698
rect 21810 21646 21812 21698
rect 2940 21586 2996 21598
rect 2940 21534 2942 21586
rect 2994 21534 2996 21586
rect 1932 21476 1988 21486
rect 1932 20914 1988 21420
rect 1932 20862 1934 20914
rect 1986 20862 1988 20914
rect 1932 20850 1988 20862
rect 2940 20916 2996 21534
rect 4844 21586 4900 21598
rect 4844 21534 4846 21586
rect 4898 21534 4900 21586
rect 3724 21474 3780 21486
rect 3724 21422 3726 21474
rect 3778 21422 3780 21474
rect 2940 20850 2996 20860
rect 3612 20916 3668 20926
rect 3612 20822 3668 20860
rect 3052 20802 3108 20814
rect 3052 20750 3054 20802
rect 3106 20750 3108 20802
rect 3052 20692 3108 20750
rect 3724 20804 3780 21422
rect 4844 21476 4900 21534
rect 4844 21410 4900 21420
rect 5404 21476 5460 21486
rect 5404 21382 5460 21420
rect 19628 21476 19684 21486
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 3724 20738 3780 20748
rect 3052 20626 3108 20636
rect 4060 20692 4116 20702
rect 4060 20598 4116 20636
rect 19628 20244 19684 21420
rect 21756 20916 21812 21646
rect 22092 21588 22148 21598
rect 22092 21494 22148 21532
rect 23100 21588 23156 21598
rect 21756 20850 21812 20860
rect 20972 20804 21028 20814
rect 20972 20578 21028 20748
rect 21868 20804 21924 20814
rect 21868 20710 21924 20748
rect 22764 20804 22820 20814
rect 22764 20710 22820 20748
rect 21644 20692 21700 20702
rect 21644 20598 21700 20636
rect 20972 20526 20974 20578
rect 21026 20526 21028 20578
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19964 20244 20020 20254
rect 19628 20242 20020 20244
rect 19628 20190 19966 20242
rect 20018 20190 20020 20242
rect 19628 20188 20020 20190
rect 19964 20178 20020 20188
rect 1932 20132 1988 20142
rect 1932 20038 1988 20076
rect 3052 20018 3108 20030
rect 3052 19966 3054 20018
rect 3106 19966 3108 20018
rect 3052 19908 3108 19966
rect 19516 20020 19572 20030
rect 19516 19926 19572 19964
rect 20300 20020 20356 20030
rect 3052 19842 3108 19852
rect 3612 19908 3668 19918
rect 3612 19814 3668 19852
rect 19628 19908 19684 19918
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 1932 19460 1988 19470
rect 1932 19346 1988 19404
rect 1932 19294 1934 19346
rect 1986 19294 1988 19346
rect 1932 19282 1988 19294
rect 3052 19234 3108 19246
rect 3052 19182 3054 19234
rect 3106 19182 3108 19234
rect 3052 18900 3108 19182
rect 18956 19234 19012 19246
rect 18956 19182 18958 19234
rect 19010 19182 19012 19234
rect 3052 18834 3108 18844
rect 3612 19010 3668 19022
rect 3612 18958 3614 19010
rect 3666 18958 3668 19010
rect 3612 18900 3668 18958
rect 18284 19012 18340 19022
rect 18284 18918 18340 18956
rect 18732 19010 18788 19022
rect 18732 18958 18734 19010
rect 18786 18958 18788 19010
rect 3612 18834 3668 18844
rect 18732 18900 18788 18958
rect 18732 18834 18788 18844
rect 18956 19012 19012 19182
rect 19628 19122 19684 19852
rect 19628 19070 19630 19122
rect 19682 19070 19684 19122
rect 19628 19058 19684 19070
rect 19964 19122 20020 19134
rect 19964 19070 19966 19122
rect 20018 19070 20020 19122
rect 19964 19012 20020 19070
rect 19964 18956 20244 19012
rect 1932 18788 1988 18798
rect 1932 18562 1988 18732
rect 18956 18676 19012 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 18732 18620 19012 18676
rect 1932 18510 1934 18562
rect 1986 18510 1988 18562
rect 1932 18498 1988 18510
rect 18620 18562 18676 18574
rect 18620 18510 18622 18562
rect 18674 18510 18676 18562
rect 3052 18450 3108 18462
rect 3052 18398 3054 18450
rect 3106 18398 3108 18450
rect 3052 18340 3108 18398
rect 3052 18274 3108 18284
rect 3612 18340 3668 18350
rect 3612 18246 3668 18284
rect 18172 18338 18228 18350
rect 18172 18286 18174 18338
rect 18226 18286 18228 18338
rect 1932 18116 1988 18126
rect 1932 17778 1988 18060
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17726 1934 17778
rect 1986 17726 1988 17778
rect 1932 17714 1988 17726
rect 3052 17666 3108 17678
rect 3052 17614 3054 17666
rect 3106 17614 3108 17666
rect 1932 17444 1988 17454
rect 1932 16994 1988 17388
rect 3052 17332 3108 17614
rect 17164 17668 17220 17678
rect 17164 17666 17780 17668
rect 17164 17614 17166 17666
rect 17218 17614 17780 17666
rect 17164 17612 17780 17614
rect 17164 17602 17220 17612
rect 17724 17556 17780 17612
rect 17948 17556 18004 17566
rect 18172 17556 18228 18286
rect 18620 18340 18676 18510
rect 18620 18274 18676 18284
rect 18508 17556 18564 17566
rect 17724 17554 18564 17556
rect 17724 17502 17950 17554
rect 18002 17502 18510 17554
rect 18562 17502 18564 17554
rect 17724 17500 18564 17502
rect 17948 17490 18004 17500
rect 3052 17266 3108 17276
rect 3612 17442 3668 17454
rect 3612 17390 3614 17442
rect 3666 17390 3668 17442
rect 3612 17332 3668 17390
rect 3612 17266 3668 17276
rect 16380 17442 16436 17454
rect 16380 17390 16382 17442
rect 16434 17390 16436 17442
rect 1932 16942 1934 16994
rect 1986 16942 1988 16994
rect 1932 16930 1988 16942
rect 3052 16996 3108 17006
rect 3052 16882 3108 16940
rect 3052 16830 3054 16882
rect 3106 16830 3108 16882
rect 3052 16818 3108 16830
rect 3612 16996 3668 17006
rect 1932 16772 1988 16782
rect 1932 16210 1988 16716
rect 1932 16158 1934 16210
rect 1986 16158 1988 16210
rect 1932 16146 1988 16158
rect 3612 16210 3668 16940
rect 15708 16994 15764 17006
rect 15708 16942 15710 16994
rect 15762 16942 15764 16994
rect 4844 16884 4900 16894
rect 4844 16790 4900 16828
rect 5404 16884 5460 16894
rect 5404 16790 5460 16828
rect 3612 16158 3614 16210
rect 3666 16158 3668 16210
rect 3612 16146 3668 16158
rect 3724 16770 3780 16782
rect 3724 16718 3726 16770
rect 3778 16718 3780 16770
rect 3052 16098 3108 16110
rect 3052 16046 3054 16098
rect 3106 16046 3108 16098
rect 3052 15876 3108 16046
rect 3724 16100 3780 16718
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 3724 16034 3780 16044
rect 3052 15810 3108 15820
rect 4060 15876 4116 15886
rect 4060 15782 4116 15820
rect 15708 15876 15764 16942
rect 15820 16884 15876 16894
rect 15820 15986 15876 16828
rect 16044 16884 16100 16894
rect 16044 16790 16100 16828
rect 16380 16884 16436 17390
rect 17612 17442 17668 17454
rect 17612 17390 17614 17442
rect 17666 17390 17668 17442
rect 17612 17332 17668 17390
rect 17612 17266 17668 17276
rect 16604 16996 16660 17006
rect 16604 16902 16660 16940
rect 16380 16818 16436 16828
rect 16716 16884 16772 16894
rect 15820 15934 15822 15986
rect 15874 15934 15876 15986
rect 15820 15922 15876 15934
rect 16156 15988 16212 15998
rect 16156 15986 16324 15988
rect 16156 15934 16158 15986
rect 16210 15934 16324 15986
rect 16156 15932 16324 15934
rect 16156 15922 16212 15932
rect 15708 15810 15764 15820
rect 1932 15428 1988 15438
rect 1932 15334 1988 15372
rect 14700 15426 14756 15438
rect 14700 15374 14702 15426
rect 14754 15374 14756 15426
rect 3052 15314 3108 15326
rect 3052 15262 3054 15314
rect 3106 15262 3108 15314
rect 3052 15204 3108 15262
rect 3052 15138 3108 15148
rect 3612 15204 3668 15214
rect 3612 15110 3668 15148
rect 14700 15204 14756 15374
rect 14700 15138 14756 15148
rect 15036 15314 15092 15326
rect 15036 15262 15038 15314
rect 15090 15262 15092 15314
rect 15036 15204 15092 15262
rect 16268 15316 16324 15932
rect 16716 15874 16772 16828
rect 16716 15822 16718 15874
rect 16770 15822 16772 15874
rect 16380 15316 16436 15326
rect 16268 15260 16380 15316
rect 16380 15222 16436 15260
rect 15036 15138 15092 15148
rect 15484 15204 15540 15214
rect 15484 15110 15540 15148
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 1932 14756 1988 14766
rect 1932 14642 1988 14700
rect 1932 14590 1934 14642
rect 1986 14590 1988 14642
rect 1932 14578 1988 14590
rect 3052 14530 3108 14542
rect 3052 14478 3054 14530
rect 3106 14478 3108 14530
rect 3052 14308 3108 14478
rect 14364 14418 14420 14430
rect 14364 14366 14366 14418
rect 14418 14366 14420 14418
rect 3052 14242 3108 14252
rect 3612 14308 3668 14318
rect 3612 14214 3668 14252
rect 14028 14308 14084 14318
rect 14028 14214 14084 14252
rect 14364 14308 14420 14366
rect 14364 14242 14420 14252
rect 14812 14308 14868 14318
rect 14812 14214 14868 14252
rect 1932 14084 1988 14094
rect 1932 13858 1988 14028
rect 1932 13806 1934 13858
rect 1986 13806 1988 13858
rect 1932 13794 1988 13806
rect 12460 13858 12516 13870
rect 12460 13806 12462 13858
rect 12514 13806 12516 13858
rect 3052 13746 3108 13758
rect 3052 13694 3054 13746
rect 3106 13694 3108 13746
rect 3052 13636 3108 13694
rect 3052 13570 3108 13580
rect 3612 13636 3668 13646
rect 3612 13542 3668 13580
rect 12012 13634 12068 13646
rect 12012 13582 12014 13634
rect 12066 13582 12068 13634
rect 12012 13524 12068 13582
rect 12012 13458 12068 13468
rect 1932 13412 1988 13422
rect 1932 13074 1988 13356
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 1932 13022 1934 13074
rect 1986 13022 1988 13074
rect 1932 13010 1988 13022
rect 3052 12962 3108 12974
rect 3052 12910 3054 12962
rect 3106 12910 3108 12962
rect 1932 12740 1988 12750
rect 1932 12290 1988 12684
rect 3052 12740 3108 12910
rect 3052 12674 3108 12684
rect 3612 12740 3668 12750
rect 3612 12646 3668 12684
rect 12012 12738 12068 12750
rect 12012 12686 12014 12738
rect 12066 12686 12068 12738
rect 1932 12238 1934 12290
rect 1986 12238 1988 12290
rect 1932 12226 1988 12238
rect 3052 12292 3108 12302
rect 3052 12178 3108 12236
rect 3052 12126 3054 12178
rect 3106 12126 3108 12178
rect 3052 12114 3108 12126
rect 3612 12292 3668 12302
rect 1932 12068 1988 12078
rect 1932 11506 1988 12012
rect 1932 11454 1934 11506
rect 1986 11454 1988 11506
rect 1932 11442 1988 11454
rect 3052 11508 3108 11518
rect 3052 11394 3108 11452
rect 3612 11506 3668 12236
rect 11340 12290 11396 12302
rect 11340 12238 11342 12290
rect 11394 12238 11396 12290
rect 4844 12178 4900 12190
rect 4844 12126 4846 12178
rect 4898 12126 4900 12178
rect 3612 11454 3614 11506
rect 3666 11454 3668 11506
rect 3612 11442 3668 11454
rect 3724 12066 3780 12078
rect 3724 12014 3726 12066
rect 3778 12014 3780 12066
rect 3052 11342 3054 11394
rect 3106 11342 3108 11394
rect 3052 11330 3108 11342
rect 3724 11396 3780 12014
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4060 11508 4116 11518
rect 4060 11414 4116 11452
rect 3724 11330 3780 11340
rect 4844 11284 4900 12126
rect 11340 11508 11396 12238
rect 11676 12180 11732 12190
rect 12012 12180 12068 12686
rect 12460 12740 12516 13806
rect 13356 13858 13412 13870
rect 13356 13806 13358 13858
rect 13410 13806 13412 13858
rect 12796 13746 12852 13758
rect 12796 13694 12798 13746
rect 12850 13694 12852 13746
rect 12796 13524 12852 13694
rect 13356 13636 13412 13806
rect 13692 13748 13748 13758
rect 13692 13654 13748 13692
rect 14140 13748 14196 13758
rect 14140 13654 14196 13692
rect 13356 13570 13412 13580
rect 12796 13458 12852 13468
rect 14028 13524 14084 13534
rect 12460 12674 12516 12684
rect 12908 12738 12964 12750
rect 12908 12686 12910 12738
rect 12962 12686 12964 12738
rect 12236 12292 12292 12302
rect 12236 12198 12292 12236
rect 11676 12178 12068 12180
rect 11676 12126 11678 12178
rect 11730 12126 12068 12178
rect 11676 12124 12068 12126
rect 12572 12180 12628 12190
rect 11676 12114 11732 12124
rect 11340 11442 11396 11452
rect 11788 11396 11844 12124
rect 12572 12086 12628 12124
rect 12908 12180 12964 12686
rect 13468 12292 13524 12302
rect 13468 12198 13524 12236
rect 12908 12114 12964 12124
rect 13244 12180 13300 12190
rect 13244 12086 13300 12124
rect 13916 12180 13972 12190
rect 13916 12066 13972 12124
rect 13916 12014 13918 12066
rect 13970 12014 13972 12066
rect 11788 11330 11844 11340
rect 12572 11396 12628 11406
rect 4844 11218 4900 11228
rect 10668 11284 10724 11294
rect 10668 11190 10724 11228
rect 11004 11284 11060 11294
rect 11564 11284 11620 11294
rect 11004 11282 11620 11284
rect 11004 11230 11006 11282
rect 11058 11230 11566 11282
rect 11618 11230 11620 11282
rect 11004 11228 11620 11230
rect 11004 11218 11060 11228
rect 1932 10724 1988 10734
rect 1932 10630 1988 10668
rect 3052 10724 3108 10734
rect 3052 10610 3108 10668
rect 10108 10724 10164 10734
rect 10108 10630 10164 10668
rect 11452 10724 11508 10734
rect 11452 10630 11508 10668
rect 3052 10558 3054 10610
rect 3106 10558 3108 10610
rect 3052 10546 3108 10558
rect 10444 10612 10500 10622
rect 11116 10612 11172 10622
rect 10444 10610 11172 10612
rect 10444 10558 10446 10610
rect 10498 10558 11118 10610
rect 11170 10558 11172 10610
rect 10444 10556 11172 10558
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 1932 10052 1988 10062
rect 1932 9938 1988 9996
rect 1932 9886 1934 9938
rect 1986 9886 1988 9938
rect 1932 9874 1988 9886
rect 3052 9826 3108 9838
rect 3052 9774 3054 9826
rect 3106 9774 3108 9826
rect 3052 9716 3108 9774
rect 9660 9826 9716 9838
rect 9660 9774 9662 9826
rect 9714 9774 9716 9826
rect 3052 9650 3108 9660
rect 9436 9716 9492 9726
rect 9436 9622 9492 9660
rect 9660 9716 9716 9774
rect 1932 9380 1988 9390
rect 1932 9154 1988 9324
rect 1932 9102 1934 9154
rect 1986 9102 1988 9154
rect 1932 9090 1988 9102
rect 3052 9156 3108 9166
rect 3052 9042 3108 9100
rect 8652 9156 8708 9166
rect 8652 9062 8708 9100
rect 3052 8990 3054 9042
rect 3106 8990 3108 9042
rect 3052 8978 3108 8990
rect 8988 9044 9044 9054
rect 1932 8708 1988 8718
rect 1932 8370 1988 8652
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 8988 8428 9044 8988
rect 1932 8318 1934 8370
rect 1986 8318 1988 8370
rect 1932 8306 1988 8318
rect 8876 8372 9044 8428
rect 3052 8258 3108 8270
rect 3052 8206 3054 8258
rect 3106 8206 3108 8258
rect 3052 8148 3108 8206
rect 3052 8082 3108 8092
rect 8092 8148 8148 8158
rect 8092 8054 8148 8092
rect 8428 8148 8484 8158
rect 8428 8054 8484 8092
rect 1932 8036 1988 8046
rect 1932 7586 1988 7980
rect 1932 7534 1934 7586
rect 1986 7534 1988 7586
rect 1932 7522 1988 7534
rect 3052 7588 3108 7598
rect 3052 7474 3108 7532
rect 6524 7586 6580 7598
rect 6524 7534 6526 7586
rect 6578 7534 6580 7586
rect 3052 7422 3054 7474
rect 3106 7422 3108 7474
rect 3052 7410 3108 7422
rect 4844 7474 4900 7486
rect 4844 7422 4846 7474
rect 4898 7422 4900 7474
rect 1932 7364 1988 7374
rect 1932 6802 1988 7308
rect 3724 7362 3780 7374
rect 3724 7310 3726 7362
rect 3778 7310 3780 7362
rect 1932 6750 1934 6802
rect 1986 6750 1988 6802
rect 1932 6738 1988 6750
rect 3052 6804 3108 6814
rect 3052 6690 3108 6748
rect 3052 6638 3054 6690
rect 3106 6638 3108 6690
rect 3052 6626 3108 6638
rect 3724 6692 3780 7310
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 3724 6626 3780 6636
rect 4844 6580 4900 7422
rect 6524 6804 6580 7534
rect 7420 7588 7476 7598
rect 7420 7494 7476 7532
rect 8764 7588 8820 7598
rect 8764 7494 8820 7532
rect 6524 6738 6580 6748
rect 6860 7474 6916 7486
rect 6860 7422 6862 7474
rect 6914 7422 6916 7474
rect 6860 6804 6916 7422
rect 6860 6738 6916 6748
rect 7644 7476 7700 7486
rect 4844 6514 4900 6524
rect 5740 6692 5796 6702
rect 1932 6020 1988 6030
rect 1932 5926 1988 5964
rect 3052 6020 3108 6030
rect 3052 5906 3108 5964
rect 4620 6020 4676 6030
rect 4620 5926 4676 5964
rect 3052 5854 3054 5906
rect 3106 5854 3108 5906
rect 3052 5842 3108 5854
rect 4956 5906 5012 5918
rect 4956 5854 4958 5906
rect 5010 5854 5012 5906
rect 4172 5794 4228 5806
rect 4172 5742 4174 5794
rect 4226 5742 4228 5794
rect 1932 5348 1988 5358
rect 1932 5234 1988 5292
rect 1932 5182 1934 5234
rect 1986 5182 1988 5234
rect 1932 5170 1988 5182
rect 3052 5122 3108 5134
rect 3052 5070 3054 5122
rect 3106 5070 3108 5122
rect 3052 4564 3108 5070
rect 4172 4788 4228 5742
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4620 5236 4676 5246
rect 4620 5012 4676 5180
rect 4956 5124 5012 5854
rect 5516 5794 5572 5806
rect 5516 5742 5518 5794
rect 5570 5742 5572 5794
rect 5516 5236 5572 5742
rect 5516 5170 5572 5180
rect 4956 5068 5124 5124
rect 5068 5012 5124 5068
rect 4620 5010 4900 5012
rect 4620 4958 4622 5010
rect 4674 4958 4900 5010
rect 4620 4956 4900 4958
rect 4620 4946 4676 4956
rect 4172 4722 4228 4732
rect 3052 4498 3108 4508
rect 4620 4564 4676 4574
rect 4620 4470 4676 4508
rect 4844 4338 4900 4956
rect 4956 4900 5012 4910
rect 4956 4806 5012 4844
rect 4844 4286 4846 4338
rect 4898 4286 4900 4338
rect 4844 4274 4900 4286
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4956 3668 5012 3678
rect 5068 3668 5124 4956
rect 4956 3666 5124 3668
rect 4956 3614 4958 3666
rect 5010 3614 5124 3666
rect 4956 3612 5124 3614
rect 5292 4788 5348 4798
rect 4956 3602 5012 3612
rect 3948 3444 4004 3454
rect 3948 3350 4004 3388
rect 5292 800 5348 4732
rect 5740 4226 5796 6636
rect 6300 6692 6356 6702
rect 6300 6598 6356 6636
rect 6972 6692 7028 6702
rect 6972 6598 7028 6636
rect 7308 6692 7364 6702
rect 6076 6580 6132 6590
rect 6076 6486 6132 6524
rect 7308 6578 7364 6636
rect 7308 6526 7310 6578
rect 7362 6526 7364 6578
rect 7308 6514 7364 6526
rect 6860 6018 6916 6030
rect 6860 5966 6862 6018
rect 6914 5966 6916 6018
rect 6412 5012 6468 5022
rect 6412 4918 6468 4956
rect 6748 4898 6804 4910
rect 6748 4846 6750 4898
rect 6802 4846 6804 4898
rect 6748 4676 6804 4846
rect 6860 4788 6916 5966
rect 6860 4722 6916 4732
rect 7308 6020 7364 6030
rect 6748 4610 6804 4620
rect 5740 4174 5742 4226
rect 5794 4174 5796 4226
rect 5740 4162 5796 4174
rect 6748 4450 6804 4462
rect 6748 4398 6750 4450
rect 6802 4398 6804 4450
rect 5740 3444 5796 3454
rect 6748 3444 6804 4398
rect 6860 3444 6916 3454
rect 5740 3332 5796 3388
rect 6636 3442 6916 3444
rect 6636 3390 6862 3442
rect 6914 3390 6916 3442
rect 6636 3388 6916 3390
rect 5740 3276 6020 3332
rect 5964 800 6020 3276
rect 6636 800 6692 3388
rect 6860 3378 6916 3388
rect 7308 800 7364 5964
rect 7644 5234 7700 7420
rect 8428 7476 8484 7486
rect 8428 7382 8484 7420
rect 7868 6804 7924 6814
rect 7868 6690 7924 6748
rect 7868 6638 7870 6690
rect 7922 6638 7924 6690
rect 7756 5796 7812 5806
rect 7868 5796 7924 6638
rect 8204 6466 8260 6478
rect 8204 6414 8206 6466
rect 8258 6414 8260 6466
rect 8204 6132 8260 6414
rect 8204 6066 8260 6076
rect 8652 6466 8708 6478
rect 8652 6414 8654 6466
rect 8706 6414 8708 6466
rect 8652 6020 8708 6414
rect 8652 5888 8708 5964
rect 7756 5794 7924 5796
rect 7756 5742 7758 5794
rect 7810 5742 7924 5794
rect 7756 5740 7924 5742
rect 7756 5730 7812 5740
rect 7644 5182 7646 5234
rect 7698 5182 7700 5234
rect 7644 5170 7700 5182
rect 8428 5012 8484 5022
rect 8316 5010 8484 5012
rect 8316 4958 8430 5010
rect 8482 4958 8484 5010
rect 8316 4956 8484 4958
rect 7980 4450 8036 4462
rect 7980 4398 7982 4450
rect 8034 4398 8036 4450
rect 7980 3668 8036 4398
rect 7980 3602 8036 3612
rect 8092 4228 8148 4238
rect 7868 3444 7924 3454
rect 7868 3350 7924 3388
rect 8092 3332 8148 4172
rect 8316 4228 8372 4956
rect 8428 4946 8484 4956
rect 8316 4162 8372 4172
rect 7980 3276 8148 3332
rect 8652 3668 8708 3678
rect 7980 800 8036 3276
rect 8652 800 8708 3612
rect 8876 3666 8932 8372
rect 8988 8148 9044 8158
rect 9100 8148 9156 8158
rect 9044 8146 9156 8148
rect 9044 8094 9102 8146
rect 9154 8094 9156 8146
rect 9044 8092 9156 8094
rect 8988 4226 9044 8092
rect 9100 8082 9156 8092
rect 9436 8036 9492 8046
rect 9436 7942 9492 7980
rect 9660 5234 9716 9660
rect 10220 9156 10276 9166
rect 10220 9062 10276 9100
rect 9884 9044 9940 9054
rect 9884 8950 9940 8988
rect 10444 8428 10500 10556
rect 11116 10546 11172 10556
rect 10556 9716 10612 9726
rect 10556 9622 10612 9660
rect 10892 9604 10948 9614
rect 10892 9510 10948 9548
rect 10444 8372 10612 8428
rect 9660 5182 9662 5234
rect 9714 5182 9716 5234
rect 9660 5170 9716 5182
rect 10444 5012 10500 5022
rect 10108 4956 10444 5012
rect 9660 4340 9716 4350
rect 9660 4246 9716 4284
rect 8988 4174 8990 4226
rect 9042 4174 9044 4226
rect 8988 4162 9044 4174
rect 8876 3614 8878 3666
rect 8930 3614 8932 3666
rect 8876 3602 8932 3614
rect 9548 3668 9604 3678
rect 9548 3574 9604 3612
rect 9324 3444 9380 3454
rect 9324 800 9380 3388
rect 9996 3444 10052 3454
rect 9996 3350 10052 3388
rect 10108 3220 10164 4956
rect 10444 4880 10500 4956
rect 10444 4228 10500 4238
rect 10556 4228 10612 8372
rect 11116 5794 11172 5806
rect 11116 5742 11118 5794
rect 11170 5742 11172 5794
rect 11116 5012 11172 5742
rect 11116 4946 11172 4956
rect 11228 5796 11284 5806
rect 11228 4452 11284 5740
rect 11564 5234 11620 11228
rect 11900 11172 11956 11182
rect 11900 11078 11956 11116
rect 11900 5796 11956 5806
rect 11900 5702 11956 5740
rect 11564 5182 11566 5234
rect 11618 5182 11620 5234
rect 11564 5170 11620 5182
rect 10444 4226 10612 4228
rect 10444 4174 10446 4226
rect 10498 4174 10612 4226
rect 10444 4172 10612 4174
rect 10668 4450 11284 4452
rect 10668 4398 11230 4450
rect 11282 4398 11284 4450
rect 10668 4396 11284 4398
rect 10444 4162 10500 4172
rect 9996 3164 10164 3220
rect 9996 800 10052 3164
rect 10668 800 10724 4396
rect 11228 4386 11284 4396
rect 11340 5012 11396 5022
rect 10892 3444 10948 3454
rect 10892 3350 10948 3388
rect 11340 800 11396 4956
rect 12460 5012 12516 5022
rect 12460 4788 12516 4956
rect 12460 4722 12516 4732
rect 12572 3666 12628 11340
rect 13580 11396 13636 11406
rect 13580 11302 13636 11340
rect 12796 11284 12852 11294
rect 12796 11190 12852 11228
rect 13916 8428 13972 12014
rect 13580 8372 13972 8428
rect 12572 3614 12574 3666
rect 12626 3614 12628 3666
rect 12572 3602 12628 3614
rect 12684 5796 12740 5806
rect 12684 4450 12740 5740
rect 13468 5794 13524 5806
rect 13468 5742 13470 5794
rect 13522 5742 13524 5794
rect 13468 5012 13524 5742
rect 13468 4946 13524 4956
rect 12684 4398 12686 4450
rect 12738 4398 12740 4450
rect 11676 3444 11732 3454
rect 11732 3388 12068 3444
rect 11676 3312 11732 3388
rect 12012 800 12068 3388
rect 12684 800 12740 4398
rect 13580 4226 13636 8372
rect 13916 5796 13972 5806
rect 13916 5702 13972 5740
rect 13580 4174 13582 4226
rect 13634 4174 13636 4226
rect 13580 4162 13636 4174
rect 13692 5012 13748 5022
rect 13692 3780 13748 4956
rect 14028 5010 14084 13468
rect 16716 8428 16772 15822
rect 16940 16882 16996 16894
rect 16940 16830 16942 16882
rect 16994 16830 16996 16882
rect 16940 15876 16996 16830
rect 18172 16882 18228 16894
rect 18172 16830 18174 16882
rect 18226 16830 18228 16882
rect 17612 16770 17668 16782
rect 17612 16718 17614 16770
rect 17666 16718 17668 16770
rect 17164 15876 17220 15886
rect 16940 15874 17220 15876
rect 16940 15822 17166 15874
rect 17218 15822 17220 15874
rect 16940 15820 17220 15822
rect 17164 15428 17220 15820
rect 17612 15428 17668 16718
rect 18060 16100 18116 16110
rect 18172 16100 18228 16830
rect 18060 16098 18228 16100
rect 18060 16046 18062 16098
rect 18114 16046 18228 16098
rect 18060 16044 18228 16046
rect 18284 16100 18340 16110
rect 18396 16100 18452 17500
rect 18508 17490 18564 17500
rect 18732 17108 18788 18620
rect 18956 18450 19012 18462
rect 18956 18398 18958 18450
rect 19010 18398 19012 18450
rect 18844 17556 18900 17566
rect 18844 17462 18900 17500
rect 18732 17042 18788 17052
rect 18956 17332 19012 18398
rect 20188 18452 20244 18956
rect 19740 18340 19796 18350
rect 19628 18338 19796 18340
rect 19628 18286 19742 18338
rect 19794 18286 19796 18338
rect 19628 18284 19796 18286
rect 19292 17442 19348 17454
rect 19292 17390 19294 17442
rect 19346 17390 19348 17442
rect 19292 17332 19348 17390
rect 19628 17332 19684 18284
rect 19740 18274 19796 18284
rect 20188 18338 20244 18396
rect 20188 18286 20190 18338
rect 20242 18286 20244 18338
rect 18956 17276 19684 17332
rect 20188 17666 20244 18286
rect 20188 17614 20190 17666
rect 20242 17614 20244 17666
rect 20188 17332 20244 17614
rect 20300 17668 20356 19964
rect 20860 20020 20916 20030
rect 20860 19926 20916 19964
rect 20524 19122 20580 19134
rect 20524 19070 20526 19122
rect 20578 19070 20580 19122
rect 20524 18452 20580 19070
rect 20860 19012 20916 19022
rect 20860 18918 20916 18956
rect 20860 18676 20916 18686
rect 20748 18452 20804 18462
rect 20524 18386 20580 18396
rect 20636 18450 20804 18452
rect 20636 18398 20750 18450
rect 20802 18398 20804 18450
rect 20636 18396 20804 18398
rect 20300 17574 20356 17612
rect 20524 17668 20580 17678
rect 20636 17668 20692 18396
rect 20748 18386 20804 18396
rect 20748 17892 20804 17902
rect 20860 17892 20916 18620
rect 20972 18004 21028 20526
rect 21196 20244 21252 20282
rect 23100 20188 23156 21532
rect 23660 21588 23716 21598
rect 23660 21494 23716 21532
rect 23212 20804 23268 20814
rect 23212 20710 23268 20748
rect 23548 20580 23604 20590
rect 23548 20486 23604 20524
rect 23772 20188 23828 22094
rect 24220 22146 24388 22148
rect 24220 22094 24334 22146
rect 24386 22094 24388 22146
rect 24220 22092 24388 22094
rect 24220 21812 24276 22092
rect 24332 22082 24388 22092
rect 24444 21924 24500 24668
rect 24556 24658 24612 24668
rect 24892 24724 24948 24782
rect 24892 24658 24948 24668
rect 25900 24724 25956 25116
rect 26124 24836 26180 24846
rect 26124 24742 26180 24780
rect 25900 24722 26068 24724
rect 25900 24670 25902 24722
rect 25954 24670 26068 24722
rect 25900 24668 26068 24670
rect 25900 24658 25956 24668
rect 25340 23826 25396 23838
rect 25340 23774 25342 23826
rect 25394 23774 25396 23826
rect 24892 23716 24948 23726
rect 25340 23716 25396 23774
rect 24892 23714 25396 23716
rect 24892 23662 24894 23714
rect 24946 23662 25396 23714
rect 24892 23660 25396 23662
rect 25676 23716 25732 23726
rect 23996 21700 24052 21710
rect 23996 21606 24052 21644
rect 21196 20178 21252 20188
rect 22988 20132 23156 20188
rect 23436 20132 23828 20188
rect 23884 21588 23940 21598
rect 21644 20020 21700 20030
rect 21644 19926 21700 19964
rect 21644 19122 21700 19134
rect 21644 19070 21646 19122
rect 21698 19070 21700 19122
rect 21532 18676 21588 18686
rect 21644 18676 21700 19070
rect 21980 19124 22036 19134
rect 21980 19030 22036 19068
rect 21588 18620 21700 18676
rect 22428 19010 22484 19022
rect 22428 18958 22430 19010
rect 22482 18958 22484 19010
rect 21084 18562 21140 18574
rect 21084 18510 21086 18562
rect 21138 18510 21140 18562
rect 21532 18544 21588 18620
rect 21084 18452 21140 18510
rect 21084 18386 21140 18396
rect 20972 17948 21252 18004
rect 20748 17890 21140 17892
rect 20748 17838 20750 17890
rect 20802 17838 21140 17890
rect 20748 17836 21140 17838
rect 20748 17826 20804 17836
rect 20524 17666 20692 17668
rect 20524 17614 20526 17666
rect 20578 17614 20692 17666
rect 20524 17612 20692 17614
rect 18508 16996 18564 17006
rect 18508 16902 18564 16940
rect 18732 16884 18788 16894
rect 18732 16322 18788 16828
rect 18732 16270 18734 16322
rect 18786 16270 18788 16322
rect 18732 16258 18788 16270
rect 18284 16098 18452 16100
rect 18284 16046 18286 16098
rect 18338 16046 18452 16098
rect 18284 16044 18452 16046
rect 18508 16098 18564 16110
rect 18508 16046 18510 16098
rect 18562 16046 18564 16098
rect 18060 15428 18116 16044
rect 18172 15428 18228 15438
rect 17164 15426 18228 15428
rect 17164 15374 18174 15426
rect 18226 15374 18228 15426
rect 17164 15372 18228 15374
rect 17052 15316 17108 15326
rect 17052 15092 17108 15260
rect 16940 14308 16996 14318
rect 16268 8372 16772 8428
rect 16828 13748 16884 13758
rect 16268 6802 16324 8372
rect 16268 6750 16270 6802
rect 16322 6750 16324 6802
rect 16268 6738 16324 6750
rect 15932 6020 15988 6030
rect 15932 6018 16100 6020
rect 15932 5966 15934 6018
rect 15986 5966 16100 6018
rect 15932 5964 16100 5966
rect 15932 5954 15988 5964
rect 16044 5908 16100 5964
rect 14476 5796 14532 5806
rect 14028 4958 14030 5010
rect 14082 4958 14084 5010
rect 14028 4946 14084 4958
rect 14364 5794 14532 5796
rect 14364 5742 14478 5794
rect 14530 5742 14532 5794
rect 14364 5740 14532 5742
rect 14364 4452 14420 5740
rect 14476 5730 14532 5740
rect 14476 5122 14532 5134
rect 14476 5070 14478 5122
rect 14530 5070 14532 5122
rect 14476 4788 14532 5070
rect 15820 5012 15876 5022
rect 15820 4918 15876 4956
rect 14476 4722 14532 4732
rect 13356 3724 13748 3780
rect 14028 4450 14420 4452
rect 14028 4398 14366 4450
rect 14418 4398 14420 4450
rect 14028 4396 14420 4398
rect 13356 800 13412 3724
rect 13804 3444 13860 3454
rect 13804 3350 13860 3388
rect 14028 800 14084 4396
rect 14364 4386 14420 4396
rect 14700 3444 14756 3454
rect 14700 800 14756 3388
rect 15372 3444 15428 3454
rect 15372 800 15428 3388
rect 16044 800 16100 5852
rect 16716 5796 16772 5806
rect 16716 5702 16772 5740
rect 16604 5684 16660 5694
rect 16604 5012 16660 5628
rect 16716 5236 16772 5246
rect 16716 5142 16772 5180
rect 16604 4956 16772 5012
rect 16716 800 16772 4956
rect 16828 4562 16884 13692
rect 16828 4510 16830 4562
rect 16882 4510 16884 4562
rect 16828 4498 16884 4510
rect 16828 3780 16884 3790
rect 16940 3780 16996 14252
rect 17052 5796 17108 15036
rect 17052 5730 17108 5740
rect 17164 5236 17220 15372
rect 18172 15362 18228 15372
rect 18284 15428 18340 16044
rect 18284 15362 18340 15372
rect 18508 15876 18564 16046
rect 18844 16100 18900 16110
rect 18844 16006 18900 16044
rect 18956 15876 19012 17276
rect 19292 17108 19348 17118
rect 19628 17108 19684 17276
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20188 17266 20244 17276
rect 19836 17210 20100 17220
rect 19964 17108 20020 17118
rect 20524 17108 20580 17612
rect 20860 17554 20916 17566
rect 20860 17502 20862 17554
rect 20914 17502 20916 17554
rect 20860 17444 20916 17502
rect 20860 17378 20916 17388
rect 19628 17106 20580 17108
rect 19628 17054 19966 17106
rect 20018 17054 20580 17106
rect 19628 17052 20580 17054
rect 20860 17220 20916 17230
rect 19180 16884 19236 16894
rect 19180 16790 19236 16828
rect 18508 15316 18564 15820
rect 18508 15250 18564 15260
rect 18844 15820 19012 15876
rect 17724 15202 17780 15214
rect 17724 15150 17726 15202
rect 17778 15150 17780 15202
rect 17724 15092 17780 15150
rect 17724 15026 17780 15036
rect 18844 8428 18900 15820
rect 19292 15540 19348 17052
rect 19964 17042 20020 17052
rect 19516 16994 19572 17006
rect 19516 16942 19518 16994
rect 19570 16942 19572 16994
rect 19516 16212 19572 16942
rect 20412 16884 20468 16894
rect 20412 16790 20468 16828
rect 19516 16146 19572 16156
rect 20748 16772 20804 16782
rect 19404 15986 19460 15998
rect 19404 15934 19406 15986
rect 19458 15934 19460 15986
rect 19404 15876 19460 15934
rect 20188 15988 20244 15998
rect 19404 15810 19460 15820
rect 19740 15876 19796 15914
rect 20188 15894 20244 15932
rect 19740 15810 19796 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 18620 8372 18900 8428
rect 18956 15484 19348 15540
rect 18060 7362 18116 7374
rect 18060 7310 18062 7362
rect 18114 7310 18116 7362
rect 17276 6578 17332 6590
rect 17276 6526 17278 6578
rect 17330 6526 17332 6578
rect 17276 5684 17332 6526
rect 18060 6580 18116 7310
rect 18508 6580 18564 6590
rect 18060 6578 18564 6580
rect 18060 6526 18510 6578
rect 18562 6526 18564 6578
rect 18060 6524 18564 6526
rect 17276 5618 17332 5628
rect 17948 5794 18004 5806
rect 17948 5742 17950 5794
rect 18002 5742 18004 5794
rect 17948 5684 18004 5742
rect 17948 5618 18004 5628
rect 17164 5170 17220 5180
rect 16828 3778 16996 3780
rect 16828 3726 16830 3778
rect 16882 3726 16996 3778
rect 16828 3724 16996 3726
rect 17388 5012 17444 5022
rect 17388 4228 17444 4956
rect 17836 5012 17892 5022
rect 17836 4918 17892 4956
rect 17612 4228 17668 4238
rect 17388 4226 17668 4228
rect 17388 4174 17614 4226
rect 17666 4174 17668 4226
rect 17388 4172 17668 4174
rect 16828 3714 16884 3724
rect 17388 800 17444 4172
rect 17612 4162 17668 4172
rect 18060 4226 18116 4238
rect 18060 4174 18062 4226
rect 18114 4174 18116 4226
rect 17612 3444 17668 3454
rect 17612 3350 17668 3388
rect 18060 3444 18116 4174
rect 18060 3378 18116 3388
rect 18284 3220 18340 6524
rect 18508 6514 18564 6524
rect 18396 5908 18452 5918
rect 18396 5814 18452 5852
rect 18620 5234 18676 8372
rect 18956 5794 19012 15484
rect 19068 15316 19124 15326
rect 19068 15202 19124 15260
rect 19068 15150 19070 15202
rect 19122 15150 19124 15202
rect 19068 8428 19124 15150
rect 19628 15204 19684 15214
rect 19068 8372 19572 8428
rect 19516 6802 19572 8372
rect 19516 6750 19518 6802
rect 19570 6750 19572 6802
rect 19516 6738 19572 6750
rect 18956 5742 18958 5794
rect 19010 5742 19012 5794
rect 18956 5730 19012 5742
rect 19404 6020 19460 6030
rect 18620 5182 18622 5234
rect 18674 5182 18676 5234
rect 18620 5170 18676 5182
rect 18060 3164 18340 3220
rect 18732 5012 18788 5022
rect 18732 4228 18788 4956
rect 18844 4228 18900 4238
rect 18732 4226 18900 4228
rect 18732 4174 18846 4226
rect 18898 4174 18900 4226
rect 18732 4172 18900 4174
rect 18060 800 18116 3164
rect 18732 800 18788 4172
rect 18844 4162 18900 4172
rect 19404 800 19460 5964
rect 19516 5236 19572 5246
rect 19516 5010 19572 5180
rect 19516 4958 19518 5010
rect 19570 4958 19572 5010
rect 19516 2996 19572 4958
rect 19628 3668 19684 15148
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20636 6466 20692 6478
rect 20636 6414 20638 6466
rect 20690 6414 20692 6466
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20300 6020 20356 6030
rect 20636 6020 20692 6414
rect 20356 5964 20692 6020
rect 20300 5888 20356 5964
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19852 4452 19908 4462
rect 19852 4358 19908 4396
rect 20748 4226 20804 16716
rect 20860 5234 20916 17164
rect 21084 17108 21140 17836
rect 21084 16976 21140 17052
rect 21196 16772 21252 17948
rect 21196 16706 21252 16716
rect 21532 17668 21588 17678
rect 21532 17442 21588 17612
rect 21532 17390 21534 17442
rect 21586 17390 21588 17442
rect 21532 8428 21588 17390
rect 21980 17442 22036 17454
rect 21980 17390 21982 17442
rect 22034 17390 22036 17442
rect 21980 17220 22036 17390
rect 21980 17154 22036 17164
rect 22428 17220 22484 18958
rect 22428 17154 22484 17164
rect 22316 16772 22372 16782
rect 22316 16678 22372 16716
rect 22988 16770 23044 20132
rect 22988 16718 22990 16770
rect 23042 16718 23044 16770
rect 22988 16706 23044 16718
rect 23100 17220 23156 17230
rect 22876 16658 22932 16670
rect 22876 16606 22878 16658
rect 22930 16606 22932 16658
rect 22876 16322 22932 16606
rect 22876 16270 22878 16322
rect 22930 16270 22932 16322
rect 22876 16258 22932 16270
rect 22652 16100 22708 16110
rect 22652 16006 22708 16044
rect 20972 8372 21588 8428
rect 22652 15764 22708 15774
rect 20972 5794 21028 8372
rect 22428 6580 22484 6590
rect 22092 6578 22484 6580
rect 22092 6526 22430 6578
rect 22482 6526 22484 6578
rect 22092 6524 22484 6526
rect 21868 6468 21924 6478
rect 22092 6468 22148 6524
rect 22428 6514 22484 6524
rect 21868 6466 22148 6468
rect 21868 6414 21870 6466
rect 21922 6414 22148 6466
rect 21868 6412 22148 6414
rect 21868 6402 21924 6412
rect 21980 6020 22036 6030
rect 20972 5742 20974 5794
rect 21026 5742 21028 5794
rect 20972 5730 21028 5742
rect 21644 6018 22036 6020
rect 21644 5966 21982 6018
rect 22034 5966 22036 6018
rect 21644 5964 22036 5966
rect 20860 5182 20862 5234
rect 20914 5182 20916 5234
rect 20860 5170 20916 5182
rect 20748 4174 20750 4226
rect 20802 4174 20804 4226
rect 20748 4162 20804 4174
rect 20972 5124 21028 5134
rect 20972 4004 21028 5068
rect 21644 5124 21700 5964
rect 21980 5954 22036 5964
rect 21980 5236 22036 5246
rect 21980 5142 22036 5180
rect 21644 5030 21700 5068
rect 20748 3948 21028 4004
rect 21308 4452 21364 4462
rect 19740 3668 19796 3678
rect 19628 3666 19796 3668
rect 19628 3614 19742 3666
rect 19794 3614 19796 3666
rect 19628 3612 19796 3614
rect 19740 3602 19796 3612
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 19516 2940 20132 2996
rect 20076 800 20132 2940
rect 20748 800 20804 3948
rect 21308 3668 21364 4396
rect 21868 4450 21924 4462
rect 21868 4398 21870 4450
rect 21922 4398 21924 4450
rect 21308 3666 21476 3668
rect 21308 3614 21310 3666
rect 21362 3614 21476 3666
rect 21308 3612 21476 3614
rect 21308 3602 21364 3612
rect 21420 800 21476 3612
rect 21868 3556 21924 4398
rect 21868 3490 21924 3500
rect 22092 800 22148 6412
rect 22652 4226 22708 15708
rect 23100 8428 23156 17164
rect 23324 17108 23380 17118
rect 23212 16772 23268 16782
rect 23212 16678 23268 16716
rect 23212 16324 23268 16334
rect 23324 16324 23380 17052
rect 23212 16322 23380 16324
rect 23212 16270 23214 16322
rect 23266 16270 23380 16322
rect 23212 16268 23380 16270
rect 23436 16658 23492 20132
rect 23660 16884 23716 16894
rect 23660 16790 23716 16828
rect 23436 16606 23438 16658
rect 23490 16606 23492 16658
rect 23212 16258 23268 16268
rect 23436 15764 23492 16606
rect 23436 15698 23492 15708
rect 23884 15874 23940 21532
rect 24108 17444 24164 17454
rect 24220 17444 24276 21756
rect 24332 21868 24500 21924
rect 24556 22820 24612 22830
rect 24892 22820 24948 23660
rect 25676 23622 25732 23660
rect 26012 23716 26068 24668
rect 26572 24610 26628 25452
rect 27132 25396 27188 26236
rect 27020 25394 27188 25396
rect 27020 25342 27134 25394
rect 27186 25342 27188 25394
rect 27020 25340 27188 25342
rect 26684 25284 26740 25294
rect 26684 25190 26740 25228
rect 26572 24558 26574 24610
rect 26626 24558 26628 24610
rect 26124 23716 26180 23726
rect 26012 23714 26180 23716
rect 26012 23662 26126 23714
rect 26178 23662 26180 23714
rect 26012 23660 26180 23662
rect 24612 22764 24948 22820
rect 24332 20188 24388 21868
rect 24444 21588 24500 21598
rect 24444 21494 24500 21532
rect 24556 20188 24612 22764
rect 26012 20188 26068 23660
rect 26124 23650 26180 23660
rect 24332 20132 24500 20188
rect 24556 20132 24724 20188
rect 24108 17442 24276 17444
rect 24108 17390 24110 17442
rect 24162 17390 24276 17442
rect 24108 17388 24276 17390
rect 24108 17378 24164 17388
rect 23884 15822 23886 15874
rect 23938 15822 23940 15874
rect 23884 8428 23940 15822
rect 23100 8372 23380 8428
rect 23100 6020 23156 6030
rect 22652 4174 22654 4226
rect 22706 4174 22708 4226
rect 22652 4162 22708 4174
rect 22764 6018 23156 6020
rect 22764 5966 23102 6018
rect 23154 5966 23156 6018
rect 22764 5964 23156 5966
rect 22764 5122 22820 5964
rect 23100 5954 23156 5964
rect 22764 5070 22766 5122
rect 22818 5070 22820 5122
rect 22540 3556 22596 3566
rect 22540 3462 22596 3500
rect 22764 800 22820 5070
rect 23324 4228 23380 8372
rect 23660 8372 23940 8428
rect 24220 16884 24276 17388
rect 24444 17220 24500 20132
rect 24444 17106 24500 17164
rect 24444 17054 24446 17106
rect 24498 17054 24500 17106
rect 24444 17042 24500 17054
rect 23660 6802 23716 8372
rect 23660 6750 23662 6802
rect 23714 6750 23716 6802
rect 23660 6738 23716 6750
rect 24220 5794 24276 16828
rect 24668 16884 24724 20132
rect 25900 20132 26068 20188
rect 25900 17554 25956 20132
rect 25900 17502 25902 17554
rect 25954 17502 25956 17554
rect 25004 17444 25060 17454
rect 25340 17444 25396 17454
rect 25900 17444 25956 17502
rect 26236 17778 26292 17790
rect 26236 17726 26238 17778
rect 26290 17726 26292 17778
rect 25004 17442 25284 17444
rect 25004 17390 25006 17442
rect 25058 17390 25284 17442
rect 25004 17388 25284 17390
rect 25004 17378 25060 17388
rect 25228 17332 25284 17388
rect 24892 16884 24948 16894
rect 24668 16828 24892 16884
rect 24332 15874 24388 15886
rect 24332 15822 24334 15874
rect 24386 15822 24388 15874
rect 24332 15764 24388 15822
rect 24332 15698 24388 15708
rect 24220 5742 24222 5794
rect 24274 5742 24276 5794
rect 24220 5730 24276 5742
rect 24332 13412 24388 13422
rect 23772 5012 23828 5022
rect 23772 5010 24164 5012
rect 23772 4958 23774 5010
rect 23826 4958 24164 5010
rect 23772 4956 24164 4958
rect 23772 4946 23828 4956
rect 23436 4228 23492 4238
rect 23324 4226 23492 4228
rect 23324 4174 23438 4226
rect 23490 4174 23492 4226
rect 23324 4172 23492 4174
rect 23436 4162 23492 4172
rect 24108 4228 24164 4956
rect 23324 3556 23380 3566
rect 23324 2884 23380 3500
rect 23436 3444 23492 3454
rect 23436 3350 23492 3388
rect 23324 2828 23492 2884
rect 23436 800 23492 2828
rect 24108 800 24164 4172
rect 24332 3666 24388 13356
rect 24668 5234 24724 16828
rect 24892 16752 24948 16828
rect 25228 8428 25284 17276
rect 25340 17442 25956 17444
rect 25340 17390 25342 17442
rect 25394 17390 25956 17442
rect 25340 17388 25956 17390
rect 26012 17444 26068 17454
rect 25340 13412 25396 17388
rect 25676 17220 25732 17230
rect 25676 16882 25732 17164
rect 26012 16994 26068 17388
rect 26124 17442 26180 17454
rect 26124 17390 26126 17442
rect 26178 17390 26180 17442
rect 26124 17332 26180 17390
rect 26124 17266 26180 17276
rect 26012 16942 26014 16994
rect 26066 16942 26068 16994
rect 26012 16930 26068 16942
rect 25676 16830 25678 16882
rect 25730 16830 25732 16882
rect 25676 16818 25732 16830
rect 25900 16884 25956 16894
rect 25900 16790 25956 16828
rect 26236 16882 26292 17726
rect 26572 17332 26628 24558
rect 26572 17266 26628 17276
rect 26236 16830 26238 16882
rect 26290 16830 26292 16882
rect 26236 16818 26292 16830
rect 26684 16884 26740 16894
rect 26684 16790 26740 16828
rect 25340 13346 25396 13356
rect 25228 8372 25508 8428
rect 24668 5182 24670 5234
rect 24722 5182 24724 5234
rect 24668 5170 24724 5182
rect 25452 5234 25508 8372
rect 27020 6802 27076 25340
rect 27132 25330 27188 25340
rect 27020 6750 27022 6802
rect 27074 6750 27076 6802
rect 27020 6738 27076 6750
rect 25452 5182 25454 5234
rect 25506 5182 25508 5234
rect 25452 5170 25508 5182
rect 26572 6580 26628 6590
rect 26572 6466 26628 6524
rect 26572 6414 26574 6466
rect 26626 6414 26628 6466
rect 24332 3614 24334 3666
rect 24386 3614 24388 3666
rect 24332 3602 24388 3614
rect 24780 4450 24836 4462
rect 24780 4398 24782 4450
rect 24834 4398 24836 4450
rect 24780 4340 24836 4398
rect 24780 800 24836 4284
rect 26012 4340 26068 4350
rect 26012 4246 26068 4284
rect 25564 4228 25620 4238
rect 25564 4134 25620 4172
rect 26124 4228 26180 4238
rect 25340 3444 25396 3454
rect 25396 3388 25508 3444
rect 25340 3312 25396 3388
rect 25452 800 25508 3388
rect 26124 800 26180 4172
rect 26572 4004 26628 6414
rect 27244 5796 27300 26908
rect 27356 26292 27412 26302
rect 27356 26198 27412 26236
rect 27580 26068 27636 27468
rect 27916 26964 27972 26974
rect 27916 26870 27972 26908
rect 28252 26852 28308 26862
rect 28252 26758 28308 26796
rect 27692 26404 27748 26414
rect 27692 26310 27748 26348
rect 27580 26002 27636 26012
rect 27356 25956 27412 25966
rect 27356 8428 27412 25900
rect 27468 25844 27524 25854
rect 27468 20188 27524 25788
rect 27580 25508 27636 25518
rect 27580 25414 27636 25452
rect 27468 20132 27636 20188
rect 27356 8372 27524 8428
rect 27356 5796 27412 5806
rect 27244 5794 27412 5796
rect 27244 5742 27358 5794
rect 27410 5742 27412 5794
rect 27244 5740 27412 5742
rect 27356 5730 27412 5740
rect 26684 5012 26740 5022
rect 26684 5010 26852 5012
rect 26684 4958 26686 5010
rect 26738 4958 26852 5010
rect 26684 4956 26852 4958
rect 26684 4946 26740 4956
rect 26796 4228 26852 4956
rect 26796 4134 26852 4172
rect 27468 4226 27524 8372
rect 27580 5234 27636 20132
rect 28700 8428 28756 29932
rect 28812 29922 28868 29932
rect 30044 29988 30100 31054
rect 30380 30994 30436 31006
rect 30380 30942 30382 30994
rect 30434 30942 30436 30994
rect 30380 30436 30436 30942
rect 30716 30436 30772 31502
rect 31164 31554 31220 31612
rect 31164 31502 31166 31554
rect 31218 31502 31220 31554
rect 30940 31108 30996 31118
rect 30940 31014 30996 31052
rect 31164 30436 31220 31502
rect 31612 31556 31668 31566
rect 31612 31462 31668 31500
rect 31276 30996 31332 31006
rect 31276 30902 31332 30940
rect 30380 30380 30996 30436
rect 31164 30380 31332 30436
rect 30492 30100 30548 30110
rect 30492 30006 30548 30044
rect 30940 30100 30996 30380
rect 30044 29922 30100 29932
rect 30828 29988 30884 29998
rect 30828 29894 30884 29932
rect 28924 29538 28980 29550
rect 28924 29486 28926 29538
rect 28978 29486 28980 29538
rect 28924 29316 28980 29486
rect 30380 29540 30436 29550
rect 30380 29446 30436 29484
rect 28924 29250 28980 29260
rect 29260 29428 29316 29438
rect 28924 27972 28980 27982
rect 28924 27878 28980 27916
rect 28812 26964 28868 26974
rect 28812 26870 28868 26908
rect 29260 20188 29316 29372
rect 30044 29428 30100 29438
rect 30044 29334 30100 29372
rect 30940 29428 30996 30044
rect 31052 29428 31108 29438
rect 30940 29426 31108 29428
rect 30940 29374 31054 29426
rect 31106 29374 31108 29426
rect 30940 29372 31108 29374
rect 29372 28532 29428 28542
rect 29372 28082 29428 28476
rect 29596 28532 29652 28542
rect 29596 28438 29652 28476
rect 29932 28420 29988 28430
rect 29932 28326 29988 28364
rect 29372 28030 29374 28082
rect 29426 28030 29428 28082
rect 29372 28018 29428 28030
rect 29820 27860 29876 27870
rect 29820 27766 29876 27804
rect 29260 20132 29428 20188
rect 28588 8372 28756 8428
rect 28028 6580 28084 6590
rect 28028 6486 28084 6524
rect 27580 5182 27582 5234
rect 27634 5182 27636 5234
rect 27580 5170 27636 5182
rect 27692 6020 27748 6030
rect 27468 4174 27470 4226
rect 27522 4174 27524 4226
rect 27468 4162 27524 4174
rect 26572 3948 26852 4004
rect 26796 800 26852 3948
rect 27468 3444 27524 3454
rect 27468 3350 27524 3388
rect 27692 3220 27748 5964
rect 28364 5012 28420 5022
rect 27468 3164 27748 3220
rect 28140 4956 28364 5012
rect 27468 800 27524 3164
rect 28140 800 28196 4956
rect 28364 4880 28420 4956
rect 28476 3668 28532 3678
rect 28588 3668 28644 8372
rect 28700 6020 28756 6030
rect 28700 5926 28756 5964
rect 29372 5794 29428 20132
rect 30940 8428 30996 29372
rect 31052 29362 31108 29372
rect 30604 8372 30996 8428
rect 29596 6020 29652 6030
rect 29372 5742 29374 5794
rect 29426 5742 29428 5794
rect 29372 5730 29428 5742
rect 29484 5908 29540 5918
rect 29484 5234 29540 5852
rect 29484 5182 29486 5234
rect 29538 5182 29540 5234
rect 29484 5170 29540 5182
rect 29596 4676 29652 5964
rect 30380 6020 30436 6030
rect 30380 5926 30436 5964
rect 29932 5012 29988 5022
rect 29932 4918 29988 4956
rect 29484 4620 29652 4676
rect 28700 4452 28756 4462
rect 28700 4450 28868 4452
rect 28700 4398 28702 4450
rect 28754 4398 28868 4450
rect 28700 4396 28868 4398
rect 28700 4386 28756 4396
rect 28476 3666 28644 3668
rect 28476 3614 28478 3666
rect 28530 3614 28644 3666
rect 28476 3612 28644 3614
rect 28476 3602 28532 3612
rect 28812 2548 28868 4396
rect 29148 3442 29204 3454
rect 29148 3390 29150 3442
rect 29202 3390 29204 3442
rect 29148 2548 29204 3390
rect 28812 2492 29204 2548
rect 28812 800 28868 2492
rect 29484 800 29540 4620
rect 29820 4452 29876 4462
rect 29820 4358 29876 4396
rect 30604 4226 30660 8372
rect 31052 6466 31108 6478
rect 31052 6414 31054 6466
rect 31106 6414 31108 6466
rect 31052 6020 31108 6414
rect 31052 5954 31108 5964
rect 31276 5234 31332 30380
rect 31388 30100 31444 30110
rect 31388 30006 31444 30044
rect 31724 30100 31780 30110
rect 31724 30006 31780 30044
rect 31836 29540 31892 32398
rect 32284 32340 32340 32622
rect 32284 32274 32340 32284
rect 31948 31780 32004 31790
rect 31948 31686 32004 31724
rect 32284 31108 32340 31118
rect 32284 31014 32340 31052
rect 31388 29484 31892 29540
rect 32060 30996 32116 31006
rect 32060 30324 32116 30940
rect 32172 30324 32228 30334
rect 32060 30322 32228 30324
rect 32060 30270 32174 30322
rect 32226 30270 32228 30322
rect 32060 30268 32228 30270
rect 31388 20188 31444 29484
rect 31500 29316 31556 29326
rect 31500 29222 31556 29260
rect 32060 29204 32116 30268
rect 32172 30258 32228 30268
rect 31724 29148 32116 29204
rect 31388 20132 31556 20188
rect 31276 5182 31278 5234
rect 31330 5182 31332 5234
rect 31276 5170 31332 5182
rect 30604 4174 30606 4226
rect 30658 4174 30660 4226
rect 30604 4162 30660 4174
rect 30828 5122 30884 5134
rect 30828 5070 30830 5122
rect 30882 5070 30884 5122
rect 30828 4452 30884 5070
rect 29708 3444 29764 3454
rect 29708 2212 29764 3388
rect 29708 2156 30212 2212
rect 30156 800 30212 2156
rect 30828 800 30884 4396
rect 31500 4226 31556 20132
rect 31724 8428 31780 29148
rect 32396 8428 32452 33068
rect 32508 33058 32564 33068
rect 34300 32788 34356 33292
rect 34412 33124 34468 33134
rect 34412 33030 34468 33068
rect 34412 32788 34468 32798
rect 34300 32786 34468 32788
rect 34300 32734 34414 32786
rect 34466 32734 34468 32786
rect 34300 32732 34468 32734
rect 34412 32722 34468 32732
rect 33964 32676 34020 32686
rect 33964 32582 34020 32620
rect 32508 32564 32564 32574
rect 32508 32470 32564 32508
rect 33628 32564 33684 32574
rect 33628 31948 33684 32508
rect 33516 31892 33684 31948
rect 33516 31890 33572 31892
rect 33516 31838 33518 31890
rect 33570 31838 33572 31890
rect 33516 31826 33572 31838
rect 32844 31780 32900 31790
rect 32844 31686 32900 31724
rect 33964 31780 34020 31790
rect 33964 31686 34020 31724
rect 33068 31556 33124 31566
rect 33068 31462 33124 31500
rect 32732 30996 32788 31006
rect 32732 30902 32788 30940
rect 34860 8428 34916 33406
rect 31612 8372 31780 8428
rect 32172 8372 32452 8428
rect 34524 8372 34916 8428
rect 31612 5794 31668 8372
rect 31612 5742 31614 5794
rect 31666 5742 31668 5794
rect 31612 5730 31668 5742
rect 31500 4174 31502 4226
rect 31554 4174 31556 4226
rect 31500 4162 31556 4174
rect 31612 5460 31668 5470
rect 31388 3444 31444 3454
rect 31388 3350 31444 3388
rect 31612 1092 31668 5404
rect 32172 3666 32228 8372
rect 32396 6018 32452 6030
rect 32396 5966 32398 6018
rect 32450 5966 32452 6018
rect 32396 5460 32452 5966
rect 32396 5394 32452 5404
rect 33516 5794 33572 5806
rect 33516 5742 33518 5794
rect 33570 5742 33572 5794
rect 33516 5460 33572 5742
rect 33516 5394 33572 5404
rect 34524 5234 34580 8372
rect 34860 6020 34916 6030
rect 34636 5796 34692 5806
rect 34860 5796 34916 5964
rect 34636 5794 34916 5796
rect 34636 5742 34638 5794
rect 34690 5742 34916 5794
rect 34636 5740 34916 5742
rect 34636 5730 34692 5740
rect 34524 5182 34526 5234
rect 34578 5182 34580 5234
rect 34524 5170 34580 5182
rect 32172 3614 32174 3666
rect 32226 3614 32228 3666
rect 32172 3602 32228 3614
rect 32284 5010 32340 5022
rect 32284 4958 32286 5010
rect 32338 4958 32340 5010
rect 32284 4340 32340 4958
rect 33740 5012 33796 5022
rect 33740 5010 34244 5012
rect 33740 4958 33742 5010
rect 33794 4958 34244 5010
rect 33740 4956 34244 4958
rect 33740 4946 33796 4956
rect 32732 4452 32788 4462
rect 32732 4450 32900 4452
rect 32732 4398 32734 4450
rect 32786 4398 32900 4450
rect 32732 4396 32900 4398
rect 32732 4386 32788 4396
rect 32284 3108 32340 4284
rect 31500 1036 31668 1092
rect 32172 3052 32340 3108
rect 32844 4228 32900 4396
rect 33516 4340 33572 4350
rect 33516 4246 33572 4284
rect 31500 800 31556 1036
rect 32172 800 32228 3052
rect 32844 800 32900 4172
rect 33964 4228 34020 4238
rect 33964 4134 34020 4172
rect 34188 4228 34244 4956
rect 34524 4228 34580 4238
rect 34188 4226 34580 4228
rect 34188 4174 34526 4226
rect 34578 4174 34580 4226
rect 34188 4172 34580 4174
rect 33180 3444 33236 3454
rect 33180 3332 33236 3388
rect 33180 3276 33572 3332
rect 33516 800 33572 3276
rect 34188 800 34244 4172
rect 34524 4162 34580 4172
rect 34412 3444 34468 3454
rect 34412 3350 34468 3388
rect 34860 800 34916 5740
rect 34972 5236 35028 35644
rect 35420 35476 35476 35644
rect 35980 35700 36036 35710
rect 35980 35606 36036 35644
rect 36540 35588 36596 36316
rect 36988 35812 37044 35822
rect 36988 35718 37044 35756
rect 35420 35410 35476 35420
rect 36092 35476 36148 35486
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35308 34914 35364 34926
rect 35308 34862 35310 34914
rect 35362 34862 35364 34914
rect 35308 34804 35364 34862
rect 36092 34914 36148 35420
rect 36092 34862 36094 34914
rect 36146 34862 36148 34914
rect 36092 34850 36148 34862
rect 35084 34244 35140 34254
rect 35084 34150 35140 34188
rect 35308 34020 35364 34748
rect 36428 34804 36484 34814
rect 36428 34710 36484 34748
rect 35532 34692 35588 34702
rect 35532 34598 35588 34636
rect 36204 34132 36260 34142
rect 36204 34038 36260 34076
rect 35756 34020 35812 34030
rect 35308 34018 35812 34020
rect 35308 33966 35758 34018
rect 35810 33966 35812 34018
rect 35308 33964 35812 33966
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35756 31948 35812 33964
rect 35756 31892 36260 31948
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 36204 20188 36260 31892
rect 36204 20132 36372 20188
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 6020 35252 6030
rect 35196 5926 35252 5964
rect 36316 5794 36372 20132
rect 36540 8428 36596 35532
rect 36316 5742 36318 5794
rect 36370 5742 36372 5794
rect 36316 5730 36372 5742
rect 36428 8372 36596 8428
rect 36652 35700 36708 35710
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35308 5236 35364 5246
rect 34972 5234 35364 5236
rect 34972 5182 35310 5234
rect 35362 5182 35364 5234
rect 34972 5180 35364 5182
rect 35308 5170 35364 5180
rect 35644 5124 35700 5134
rect 35532 4450 35588 4462
rect 35532 4398 35534 4450
rect 35586 4398 35588 4450
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35532 3556 35588 4398
rect 35532 3490 35588 3500
rect 35196 3444 35252 3454
rect 35196 3350 35252 3388
rect 35644 3332 35700 5068
rect 36316 5124 36372 5134
rect 36316 5010 36372 5068
rect 36316 4958 36318 5010
rect 36370 4958 36372 5010
rect 36316 4946 36372 4958
rect 36316 3668 36372 3678
rect 36428 3668 36484 8372
rect 36540 4228 36596 4238
rect 36652 4228 36708 35644
rect 37324 31948 37380 37212
rect 38108 37268 38164 37278
rect 38108 37174 38164 37212
rect 38892 37154 38948 37884
rect 39116 37828 39172 37838
rect 39116 37734 39172 37772
rect 38892 37102 38894 37154
rect 38946 37102 38948 37154
rect 37548 36370 37604 36382
rect 37548 36318 37550 36370
rect 37602 36318 37604 36370
rect 37436 35588 37492 35598
rect 37548 35588 37604 36318
rect 37884 36260 37940 36270
rect 37884 36166 37940 36204
rect 37884 35700 37940 35710
rect 37884 35606 37940 35644
rect 38332 35700 38388 35710
rect 38332 35606 38388 35644
rect 37492 35532 37604 35588
rect 37436 35494 37492 35532
rect 37436 35364 37492 35374
rect 37436 35026 37492 35308
rect 37436 34974 37438 35026
rect 37490 34974 37492 35026
rect 37436 34962 37492 34974
rect 37324 31892 37604 31948
rect 37436 5124 37492 5134
rect 37436 5030 37492 5068
rect 36540 4226 36708 4228
rect 36540 4174 36542 4226
rect 36594 4174 36708 4226
rect 36540 4172 36708 4174
rect 37324 4228 37380 4238
rect 37548 4228 37604 31892
rect 38108 5796 38164 5806
rect 37996 4898 38052 4910
rect 37996 4846 37998 4898
rect 38050 4846 38052 4898
rect 37996 4788 38052 4846
rect 37996 4722 38052 4732
rect 37324 4226 37604 4228
rect 37324 4174 37326 4226
rect 37378 4174 37604 4226
rect 37324 4172 37604 4174
rect 38108 4450 38164 5740
rect 38780 5796 38836 5806
rect 38780 5702 38836 5740
rect 38892 5236 38948 37102
rect 38892 5170 38948 5180
rect 39116 37042 39172 37054
rect 39116 36990 39118 37042
rect 39170 36990 39172 37042
rect 38668 5010 38724 5022
rect 38668 4958 38670 5010
rect 38722 4958 38724 5010
rect 38108 4398 38110 4450
rect 38162 4398 38164 4450
rect 36540 4162 36596 4172
rect 37324 4162 37380 4172
rect 36316 3666 36484 3668
rect 36316 3614 36318 3666
rect 36370 3614 36484 3666
rect 36316 3612 36484 3614
rect 37884 3668 37940 3678
rect 36316 3602 36372 3612
rect 37884 3574 37940 3612
rect 35532 3276 35700 3332
rect 36204 3556 36260 3566
rect 35532 800 35588 3276
rect 36204 800 36260 3500
rect 36988 3556 37044 3566
rect 36988 3462 37044 3500
rect 36876 3444 36932 3454
rect 38108 3444 38164 4398
rect 36876 800 36932 3388
rect 37548 3388 38164 3444
rect 38220 4788 38276 4798
rect 37548 800 37604 3388
rect 38220 800 38276 4732
rect 38668 4788 38724 4958
rect 38668 4722 38724 4732
rect 39116 4226 39172 36990
rect 39116 4174 39118 4226
rect 39170 4174 39172 4226
rect 39116 4162 39172 4174
rect 38892 3668 38948 3678
rect 38332 3444 38388 3454
rect 38332 3350 38388 3388
rect 38892 800 38948 3612
rect 39004 3668 39060 3678
rect 39228 3668 39284 39452
rect 39788 39508 39844 39518
rect 39788 39414 39844 39452
rect 40684 39506 40740 39900
rect 40684 39454 40686 39506
rect 40738 39454 40740 39506
rect 40124 39396 40180 39406
rect 40124 39302 40180 39340
rect 39676 38948 39732 38958
rect 39676 38854 39732 38892
rect 39452 38836 39508 38846
rect 39452 37828 39508 38780
rect 40348 38724 40404 38734
rect 40684 38724 40740 39454
rect 41020 39620 41076 39630
rect 41020 39506 41076 39564
rect 41020 39454 41022 39506
rect 41074 39454 41076 39506
rect 41020 39442 41076 39454
rect 41468 39396 41524 39406
rect 41580 39396 41636 40348
rect 41468 39394 41636 39396
rect 41468 39342 41470 39394
rect 41522 39342 41636 39394
rect 41468 39340 41636 39342
rect 41468 39330 41524 39340
rect 40348 38722 40740 38724
rect 40348 38670 40350 38722
rect 40402 38670 40740 38722
rect 40348 38668 40740 38670
rect 40348 38658 40404 38668
rect 40012 37940 40068 37950
rect 40012 37846 40068 37884
rect 39564 37828 39620 37838
rect 39452 37826 39620 37828
rect 39452 37774 39566 37826
rect 39618 37774 39620 37826
rect 39452 37772 39620 37774
rect 39340 37268 39396 37278
rect 39340 37174 39396 37212
rect 39452 37042 39508 37772
rect 39564 37762 39620 37772
rect 39452 36990 39454 37042
rect 39506 36990 39508 37042
rect 39452 36978 39508 36990
rect 40236 5794 40292 5806
rect 40236 5742 40238 5794
rect 40290 5742 40292 5794
rect 39676 5236 39732 5246
rect 39676 5142 39732 5180
rect 40236 4788 40292 5742
rect 40460 5234 40516 38668
rect 40460 5182 40462 5234
rect 40514 5182 40516 5234
rect 40460 5170 40516 5182
rect 39004 3666 39284 3668
rect 39004 3614 39006 3666
rect 39058 3614 39284 3666
rect 39004 3612 39284 3614
rect 40124 4450 40180 4462
rect 40124 4398 40126 4450
rect 40178 4398 40180 4450
rect 40124 3668 40180 4398
rect 39004 3602 39060 3612
rect 40124 3602 40180 3612
rect 39564 3444 39620 3454
rect 39788 3444 39844 3454
rect 39620 3442 39844 3444
rect 39620 3390 39790 3442
rect 39842 3390 39844 3442
rect 39620 3388 39844 3390
rect 39564 800 39620 3388
rect 39788 3378 39844 3388
rect 40236 800 40292 4732
rect 41468 5010 41524 5022
rect 41468 4958 41470 5010
rect 41522 4958 41524 5010
rect 41468 4788 41524 4958
rect 41580 5012 41636 39340
rect 41580 4946 41636 4956
rect 41468 4722 41524 4732
rect 41692 4452 41748 4462
rect 41244 4450 41748 4452
rect 41244 4398 41694 4450
rect 41746 4398 41748 4450
rect 41244 4396 41748 4398
rect 41244 3442 41300 4396
rect 41692 4386 41748 4396
rect 41804 3666 41860 40572
rect 42140 40628 42196 41022
rect 42476 40964 42532 40974
rect 42476 40870 42532 40908
rect 42924 40962 42980 41804
rect 42924 40910 42926 40962
rect 42978 40910 42980 40962
rect 42140 40562 42196 40572
rect 42364 40628 42420 40638
rect 42364 40534 42420 40572
rect 41916 40516 41972 40526
rect 41916 40422 41972 40460
rect 42812 40404 42868 40414
rect 42812 40310 42868 40348
rect 41804 3614 41806 3666
rect 41858 3614 41860 3666
rect 41804 3602 41860 3614
rect 42252 5794 42308 5806
rect 42252 5742 42254 5794
rect 42306 5742 42308 5794
rect 42252 5012 42308 5742
rect 42924 5236 42980 40910
rect 43484 20188 43540 42588
rect 44268 42644 44324 42654
rect 44268 42550 44324 42588
rect 43708 42532 43764 42542
rect 43708 42438 43764 42476
rect 43596 41860 43652 41870
rect 43596 41766 43652 41804
rect 43484 20132 43652 20188
rect 42924 5170 42980 5180
rect 42588 5012 42644 5022
rect 42252 5010 42644 5012
rect 42252 4958 42590 5010
rect 42642 4958 42644 5010
rect 42252 4956 42644 4958
rect 41244 3390 41246 3442
rect 41298 3390 41300 3442
rect 41244 2660 41300 3390
rect 40908 2604 41300 2660
rect 41580 3444 41636 3454
rect 40908 800 40964 2604
rect 41580 800 41636 3388
rect 42252 800 42308 4956
rect 42588 4946 42644 4956
rect 42812 5012 42868 5022
rect 42812 4226 42868 4956
rect 42812 4174 42814 4226
rect 42866 4174 42868 4226
rect 42812 4162 42868 4174
rect 43596 4226 43652 20132
rect 43708 5236 43764 5246
rect 43708 5142 43764 5180
rect 44828 5122 44884 5134
rect 44828 5070 44830 5122
rect 44882 5070 44884 5122
rect 44828 5012 44884 5070
rect 44604 4452 44660 4462
rect 43596 4174 43598 4226
rect 43650 4174 43652 4226
rect 43596 4162 43652 4174
rect 44268 4450 44660 4452
rect 44268 4398 44606 4450
rect 44658 4398 44660 4450
rect 44268 4396 44660 4398
rect 43596 3668 43652 3678
rect 42924 3556 42980 3566
rect 42812 3444 42868 3454
rect 42812 3350 42868 3388
rect 42924 800 42980 3500
rect 43596 800 43652 3612
rect 44268 3666 44324 4396
rect 44604 4386 44660 4396
rect 44268 3614 44270 3666
rect 44322 3614 44324 3666
rect 44268 3556 44324 3614
rect 44268 3490 44324 3500
rect 44380 4228 44436 4238
rect 43708 3444 43764 3454
rect 43708 3350 43764 3388
rect 44380 3332 44436 4172
rect 44268 3276 44436 3332
rect 44828 3332 44884 4956
rect 44940 3666 44996 43374
rect 46396 8428 46452 44156
rect 46732 44100 46788 44492
rect 46732 44098 46900 44100
rect 46732 44046 46734 44098
rect 46786 44046 46900 44098
rect 46732 44044 46900 44046
rect 46732 44034 46788 44044
rect 46844 20188 46900 44044
rect 46844 20132 47012 20188
rect 46396 8372 46900 8428
rect 46732 6020 46788 6030
rect 45388 5794 45444 5806
rect 45388 5742 45390 5794
rect 45442 5742 45444 5794
rect 45388 4228 45444 5742
rect 46732 5794 46788 5964
rect 46732 5742 46734 5794
rect 46786 5742 46788 5794
rect 45612 5012 45668 5022
rect 45612 4918 45668 4956
rect 45388 4162 45444 4172
rect 45724 4450 45780 4462
rect 45724 4398 45726 4450
rect 45778 4398 45780 4450
rect 45724 4228 45780 4398
rect 45724 4162 45780 4172
rect 46284 4228 46340 4238
rect 44940 3614 44942 3666
rect 44994 3614 44996 3666
rect 44940 3602 44996 3614
rect 45948 3668 46004 3678
rect 45612 3444 45668 3454
rect 44828 3276 44996 3332
rect 44268 800 44324 3276
rect 44940 800 44996 3276
rect 45612 800 45668 3388
rect 45948 3442 46004 3612
rect 45948 3390 45950 3442
rect 46002 3390 46004 3442
rect 45948 3378 46004 3390
rect 46284 800 46340 4172
rect 46732 4004 46788 5742
rect 46844 4226 46900 8372
rect 46956 5234 47012 20132
rect 47292 6020 47348 6030
rect 47292 5926 47348 5964
rect 46956 5182 46958 5234
rect 47010 5182 47012 5234
rect 46956 5170 47012 5182
rect 47740 5236 47796 45612
rect 48188 45602 48244 45612
rect 47740 5170 47796 5180
rect 47852 45108 47908 45118
rect 47852 44996 47908 45052
rect 48300 44996 48356 45006
rect 47852 44994 48356 44996
rect 47852 44942 47854 44994
rect 47906 44942 48302 44994
rect 48354 44942 48356 44994
rect 47852 44940 48356 44942
rect 47628 5012 47684 5022
rect 46844 4174 46846 4226
rect 46898 4174 46900 4226
rect 46844 4162 46900 4174
rect 47516 5010 47684 5012
rect 47516 4958 47630 5010
rect 47682 4958 47684 5010
rect 47516 4956 47684 4958
rect 47516 4228 47572 4956
rect 47628 4946 47684 4956
rect 47516 4134 47572 4172
rect 47628 4116 47684 4126
rect 46732 3948 47012 4004
rect 46844 3668 46900 3678
rect 46844 3574 46900 3612
rect 46956 800 47012 3948
rect 47628 800 47684 4060
rect 47852 3668 47908 44940
rect 48300 44930 48356 44940
rect 48412 31948 48468 46508
rect 48860 43708 48916 47182
rect 48860 43652 49252 43708
rect 48188 31892 48468 31948
rect 48188 20188 48244 31892
rect 49196 20188 49252 43652
rect 49756 20188 49812 48078
rect 48188 20132 48468 20188
rect 49196 20132 49588 20188
rect 49756 20132 49924 20188
rect 48412 5794 48468 20132
rect 48412 5742 48414 5794
rect 48466 5742 48468 5794
rect 48412 5730 48468 5742
rect 48972 5796 49028 5806
rect 48748 5236 48804 5246
rect 48748 5142 48804 5180
rect 47852 3602 47908 3612
rect 48300 5124 48356 5134
rect 48188 3444 48244 3454
rect 48188 3350 48244 3388
rect 48300 800 48356 5068
rect 48748 4226 48804 4238
rect 48748 4174 48750 4226
rect 48802 4174 48804 4226
rect 48748 4116 48804 4174
rect 48748 4050 48804 4060
rect 48860 3668 48916 3678
rect 48860 3574 48916 3612
rect 48972 800 49028 5740
rect 49532 4226 49588 20132
rect 49644 5796 49700 5806
rect 49644 5702 49700 5740
rect 49644 5124 49700 5134
rect 49644 5030 49700 5068
rect 49868 4340 49924 20132
rect 49980 5908 50036 48412
rect 50092 48242 50148 49756
rect 50652 49812 50708 49822
rect 50876 49812 50932 50316
rect 50652 49718 50708 49756
rect 50764 49756 50932 49812
rect 50988 49812 51044 50652
rect 51100 50596 51156 50606
rect 51660 50596 51716 50606
rect 51100 50594 51716 50596
rect 51100 50542 51102 50594
rect 51154 50542 51662 50594
rect 51714 50542 51716 50594
rect 51100 50540 51716 50542
rect 51100 50530 51156 50540
rect 51660 50530 51716 50540
rect 51772 50596 51828 50606
rect 51772 50502 51828 50540
rect 51996 49924 52052 51214
rect 52332 50596 52388 50606
rect 52332 50502 52388 50540
rect 50316 49698 50372 49710
rect 50316 49646 50318 49698
rect 50370 49646 50372 49698
rect 50316 48916 50372 49646
rect 50652 49252 50708 49262
rect 50652 49138 50708 49196
rect 50652 49086 50654 49138
rect 50706 49086 50708 49138
rect 50652 49074 50708 49086
rect 50092 48190 50094 48242
rect 50146 48190 50148 48242
rect 50092 48178 50148 48190
rect 50204 48860 50372 48916
rect 50204 47572 50260 48860
rect 50540 48804 50596 48814
rect 50316 48802 50596 48804
rect 50316 48750 50542 48802
rect 50594 48750 50596 48802
rect 50316 48748 50596 48750
rect 50764 48804 50820 49756
rect 50988 49746 51044 49756
rect 51884 49868 52052 49924
rect 51548 49700 51604 49710
rect 51548 49606 51604 49644
rect 50876 49588 50932 49598
rect 51436 49588 51492 49598
rect 50876 49586 51492 49588
rect 50876 49534 50878 49586
rect 50930 49534 51438 49586
rect 51490 49534 51492 49586
rect 50876 49532 51492 49534
rect 50876 49522 50932 49532
rect 51436 49522 51492 49532
rect 51212 49252 51268 49262
rect 51212 49138 51268 49196
rect 51212 49086 51214 49138
rect 51266 49086 51268 49138
rect 51212 49074 51268 49086
rect 50764 48748 51380 48804
rect 50316 48242 50372 48748
rect 50540 48738 50596 48748
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50316 48190 50318 48242
rect 50370 48190 50372 48242
rect 50316 48178 50372 48190
rect 50092 47516 50260 47572
rect 50092 43708 50148 47516
rect 50204 47348 50260 47358
rect 50204 47254 50260 47292
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50092 43652 50260 43708
rect 49980 5842 50036 5852
rect 49868 4274 49924 4284
rect 49532 4174 49534 4226
rect 49586 4174 49588 4226
rect 49532 4162 49588 4174
rect 49644 4228 49700 4238
rect 49644 800 49700 4172
rect 50204 3780 50260 43652
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50540 5908 50596 5918
rect 50540 5814 50596 5852
rect 51212 5908 51268 5918
rect 51212 5814 51268 5852
rect 50764 5348 50820 5358
rect 50764 5122 50820 5292
rect 50764 5070 50766 5122
rect 50818 5070 50820 5122
rect 50764 5058 50820 5070
rect 50988 5236 51044 5246
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 50540 4450 50596 4462
rect 50540 4398 50542 4450
rect 50594 4398 50596 4450
rect 50540 4116 50596 4398
rect 50540 4050 50596 4060
rect 50204 3714 50260 3724
rect 50316 3668 50372 3678
rect 49868 3444 49924 3454
rect 49868 3350 49924 3388
rect 50316 800 50372 3612
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 50988 800 51044 5180
rect 51324 5122 51380 48748
rect 51884 43708 51940 49868
rect 51996 49700 52052 49710
rect 51996 49606 52052 49644
rect 51884 43652 52052 43708
rect 51996 6244 52052 43652
rect 52444 6580 52500 51772
rect 52556 51378 52612 52108
rect 52556 51326 52558 51378
rect 52610 51326 52612 51378
rect 52556 51314 52612 51326
rect 52780 51940 52836 51950
rect 52444 6514 52500 6524
rect 52780 6356 52836 51884
rect 52892 51604 52948 52894
rect 53116 52948 53172 52958
rect 53452 52948 53508 53454
rect 53564 52948 53620 52958
rect 53452 52946 53620 52948
rect 53452 52894 53566 52946
rect 53618 52894 53620 52946
rect 53452 52892 53620 52894
rect 53116 52854 53172 52892
rect 53564 52882 53620 52892
rect 52892 51538 52948 51548
rect 53004 52834 53060 52846
rect 53004 52782 53006 52834
rect 53058 52782 53060 52834
rect 53004 6468 53060 52782
rect 53340 52836 53396 52846
rect 53340 52742 53396 52780
rect 53676 52836 53732 53564
rect 54796 53508 54852 53518
rect 53676 52770 53732 52780
rect 53900 53506 54852 53508
rect 53900 53454 54798 53506
rect 54850 53454 54852 53506
rect 53900 53452 54852 53454
rect 53564 51938 53620 51950
rect 53564 51886 53566 51938
rect 53618 51886 53620 51938
rect 53340 51604 53396 51614
rect 53564 51604 53620 51886
rect 53676 51940 53732 51950
rect 53676 51846 53732 51884
rect 53788 51938 53844 51950
rect 53788 51886 53790 51938
rect 53842 51886 53844 51938
rect 53396 51548 53620 51604
rect 53676 51604 53732 51614
rect 53340 51510 53396 51548
rect 53676 51490 53732 51548
rect 53676 51438 53678 51490
rect 53730 51438 53732 51490
rect 53676 50594 53732 51438
rect 53788 51492 53844 51886
rect 53788 51426 53844 51436
rect 53676 50542 53678 50594
rect 53730 50542 53732 50594
rect 53676 50530 53732 50542
rect 53452 50372 53508 50382
rect 53452 50278 53508 50316
rect 53676 17442 53732 17454
rect 53676 17390 53678 17442
rect 53730 17390 53732 17442
rect 53676 17108 53732 17390
rect 53676 17042 53732 17052
rect 53676 14308 53732 14318
rect 53676 14214 53732 14252
rect 53004 6402 53060 6412
rect 52780 6290 52836 6300
rect 51996 6178 52052 6188
rect 53004 6244 53060 6254
rect 53004 6130 53060 6188
rect 53004 6078 53006 6130
rect 53058 6078 53060 6130
rect 53004 6066 53060 6078
rect 53340 6244 53396 6254
rect 51660 5794 51716 5806
rect 51660 5742 51662 5794
rect 51714 5742 51716 5794
rect 51660 5348 51716 5742
rect 51660 5282 51716 5292
rect 51996 5236 52052 5246
rect 51996 5142 52052 5180
rect 51324 5070 51326 5122
rect 51378 5070 51380 5122
rect 51100 3668 51156 3678
rect 51324 3668 51380 5070
rect 53004 5012 53060 5022
rect 51100 3666 51380 3668
rect 51100 3614 51102 3666
rect 51154 3614 51380 3666
rect 51100 3612 51380 3614
rect 51548 4340 51604 4350
rect 51548 3666 51604 4284
rect 52220 4228 52276 4238
rect 52220 4134 52276 4172
rect 51548 3614 51550 3666
rect 51602 3614 51604 3666
rect 51100 3602 51156 3612
rect 51548 3602 51604 3614
rect 52108 3780 52164 3790
rect 52108 3666 52164 3724
rect 52108 3614 52110 3666
rect 52162 3614 52164 3666
rect 52108 3602 52164 3614
rect 52780 3780 52836 3790
rect 51660 3556 51716 3566
rect 51660 800 51716 3500
rect 52780 3554 52836 3724
rect 52780 3502 52782 3554
rect 52834 3502 52836 3554
rect 52780 3490 52836 3502
rect 52332 3444 52388 3454
rect 52332 800 52388 3388
rect 53004 800 53060 4956
rect 53340 4338 53396 6188
rect 53900 6020 53956 53452
rect 54796 53442 54852 53452
rect 54908 53508 54964 53518
rect 54908 53414 54964 53452
rect 54124 52836 54180 52846
rect 54124 52742 54180 52780
rect 54012 52724 54068 52734
rect 54012 52274 54068 52668
rect 54236 52388 54292 52398
rect 54236 52294 54292 52332
rect 54012 52222 54014 52274
rect 54066 52222 54068 52274
rect 54012 52210 54068 52222
rect 55132 31948 55188 55020
rect 55356 55010 55412 55020
rect 55580 54964 55636 55412
rect 55692 55412 55748 56030
rect 55692 55280 55748 55356
rect 55468 54908 55636 54964
rect 54348 31892 55188 31948
rect 55244 54404 55300 54414
rect 54124 17668 54180 17678
rect 54124 17574 54180 17612
rect 54124 15204 54180 15214
rect 54124 14642 54180 15148
rect 54124 14590 54126 14642
rect 54178 14590 54180 14642
rect 54124 14578 54180 14590
rect 53900 5954 53956 5964
rect 54236 6580 54292 6590
rect 54236 6130 54292 6524
rect 54348 6244 54404 31892
rect 54908 18564 54964 18574
rect 54572 18338 54628 18350
rect 54572 18286 54574 18338
rect 54626 18286 54628 18338
rect 54572 16884 54628 18286
rect 54908 17668 54964 18508
rect 55020 18340 55076 18350
rect 55132 18340 55188 18350
rect 55020 18338 55132 18340
rect 55020 18286 55022 18338
rect 55074 18286 55132 18338
rect 55020 18284 55132 18286
rect 55020 18274 55076 18284
rect 55020 17668 55076 17678
rect 54908 17666 55076 17668
rect 54908 17614 55022 17666
rect 55074 17614 55076 17666
rect 54908 17612 55076 17614
rect 54572 16790 54628 16828
rect 54908 14530 54964 14542
rect 54908 14478 54910 14530
rect 54962 14478 54964 14530
rect 54572 13748 54628 13758
rect 54908 13748 54964 14478
rect 55020 14306 55076 17612
rect 55132 17442 55188 18284
rect 55132 17390 55134 17442
rect 55186 17390 55188 17442
rect 55132 17108 55188 17390
rect 55132 17042 55188 17052
rect 55020 14254 55022 14306
rect 55074 14254 55076 14306
rect 55020 14242 55076 14254
rect 55132 14530 55188 14542
rect 55132 14478 55134 14530
rect 55186 14478 55188 14530
rect 55132 14308 55188 14478
rect 55132 14242 55188 14252
rect 55020 13748 55076 13758
rect 54908 13692 55020 13748
rect 54572 13654 54628 13692
rect 55020 13074 55076 13692
rect 55020 13022 55022 13074
rect 55074 13022 55076 13074
rect 55020 13010 55076 13022
rect 54348 6178 54404 6188
rect 54460 6356 54516 6366
rect 54236 6078 54238 6130
rect 54290 6078 54292 6130
rect 53564 5012 53620 5022
rect 53564 4918 53620 4956
rect 54236 4900 54292 6078
rect 54460 5122 54516 6300
rect 55020 6132 55076 6142
rect 55244 6132 55300 54348
rect 55356 54292 55412 54302
rect 55356 54198 55412 54236
rect 55468 49588 55524 54908
rect 55580 53508 55636 53518
rect 55580 53414 55636 53452
rect 55580 51940 55636 51950
rect 55804 51940 55860 59612
rect 57820 59442 57876 59948
rect 58044 60004 58100 60014
rect 58044 59910 58100 59948
rect 59948 60002 60004 60060
rect 59948 59950 59950 60002
rect 60002 59950 60004 60002
rect 58156 59892 58212 59902
rect 58156 59798 58212 59836
rect 58940 59780 58996 59790
rect 58940 59778 59892 59780
rect 58940 59726 58942 59778
rect 58994 59726 59892 59778
rect 58940 59724 59892 59726
rect 58940 59714 58996 59724
rect 57820 59390 57822 59442
rect 57874 59390 57876 59442
rect 57820 59378 57876 59390
rect 59612 59556 59668 59566
rect 59612 59442 59668 59500
rect 59612 59390 59614 59442
rect 59666 59390 59668 59442
rect 59612 59378 59668 59390
rect 59836 59442 59892 59724
rect 59948 59556 60004 59950
rect 60396 60114 60452 60620
rect 60396 60062 60398 60114
rect 60450 60062 60452 60114
rect 60172 59892 60228 59902
rect 60172 59798 60228 59836
rect 59948 59490 60004 59500
rect 60060 59778 60116 59790
rect 60060 59726 60062 59778
rect 60114 59726 60116 59778
rect 59836 59390 59838 59442
rect 59890 59390 59892 59442
rect 59836 59378 59892 59390
rect 60060 59332 60116 59726
rect 59948 59276 60116 59332
rect 60284 59780 60340 59790
rect 58380 59220 58436 59230
rect 58380 59126 58436 59164
rect 58940 59220 58996 59230
rect 58940 59126 58996 59164
rect 57372 59108 57428 59118
rect 57260 58436 57316 58446
rect 57260 58342 57316 58380
rect 57148 58322 57204 58334
rect 57148 58270 57150 58322
rect 57202 58270 57204 58322
rect 56700 58212 56756 58222
rect 56700 58118 56756 58156
rect 57148 58212 57204 58270
rect 57372 58212 57428 59052
rect 59724 59106 59780 59118
rect 59724 59054 59726 59106
rect 59778 59054 59780 59106
rect 58492 58994 58548 59006
rect 58492 58942 58494 58994
rect 58546 58942 58548 58994
rect 58492 58660 58548 58942
rect 58604 58660 58660 58670
rect 58492 58658 58660 58660
rect 58492 58606 58606 58658
rect 58658 58606 58660 58658
rect 58492 58604 58660 58606
rect 58604 58594 58660 58604
rect 58156 58436 58212 58446
rect 58156 58342 58212 58380
rect 58268 58434 58324 58446
rect 58268 58382 58270 58434
rect 58322 58382 58324 58434
rect 57148 58146 57204 58156
rect 57260 58156 57428 58212
rect 57932 58210 57988 58222
rect 57932 58158 57934 58210
rect 57986 58158 57988 58210
rect 56140 57652 56196 57662
rect 56140 57558 56196 57596
rect 56028 57540 56084 57550
rect 56028 57446 56084 57484
rect 56588 57540 56644 57550
rect 56588 57446 56644 57484
rect 55916 57092 55972 57102
rect 55916 55468 55972 57036
rect 56140 56756 56196 56766
rect 56140 56662 56196 56700
rect 56588 56756 56644 56766
rect 56588 56662 56644 56700
rect 56700 56642 56756 56654
rect 56700 56590 56702 56642
rect 56754 56590 56756 56642
rect 56700 56308 56756 56590
rect 56700 56242 56756 56252
rect 56700 56084 56756 56094
rect 56700 55990 56756 56028
rect 56028 55860 56084 55870
rect 56588 55860 56644 55870
rect 56028 55858 56644 55860
rect 56028 55806 56030 55858
rect 56082 55806 56590 55858
rect 56642 55806 56644 55858
rect 56028 55804 56644 55806
rect 56028 55794 56084 55804
rect 56588 55794 56644 55804
rect 57260 55468 57316 58156
rect 57820 57876 57876 57886
rect 57932 57876 57988 58158
rect 58044 58212 58100 58222
rect 58044 58210 58212 58212
rect 58044 58158 58046 58210
rect 58098 58158 58212 58210
rect 58044 58156 58212 58158
rect 58044 58146 58100 58156
rect 57708 57874 57988 57876
rect 57708 57822 57822 57874
rect 57874 57822 57988 57874
rect 57708 57820 57988 57822
rect 57596 56868 57652 56878
rect 57596 56774 57652 56812
rect 55916 55412 56084 55468
rect 55916 55300 55972 55310
rect 55916 55206 55972 55244
rect 56028 54628 56084 55412
rect 57148 55412 57316 55468
rect 57372 56642 57428 56654
rect 57372 56590 57374 56642
rect 57426 56590 57428 56642
rect 56588 55300 56644 55310
rect 56364 55188 56420 55198
rect 56364 55074 56420 55132
rect 56364 55022 56366 55074
rect 56418 55022 56420 55074
rect 56028 54626 56196 54628
rect 56028 54574 56030 54626
rect 56082 54574 56196 54626
rect 56028 54572 56196 54574
rect 56028 54562 56084 54572
rect 55916 54292 55972 54302
rect 55916 54198 55972 54236
rect 56140 53954 56196 54572
rect 56140 53902 56142 53954
rect 56194 53902 56196 53954
rect 56140 53890 56196 53902
rect 55916 53618 55972 53630
rect 55916 53566 55918 53618
rect 55970 53566 55972 53618
rect 55916 52500 55972 53566
rect 55916 52444 56308 52500
rect 56140 52162 56196 52174
rect 56140 52110 56142 52162
rect 56194 52110 56196 52162
rect 56140 51940 56196 52110
rect 55580 51938 56196 51940
rect 55580 51886 55582 51938
rect 55634 51886 56196 51938
rect 55580 51884 56196 51886
rect 55580 51874 55636 51884
rect 55468 49522 55524 49532
rect 55692 51380 55748 51390
rect 55692 51266 55748 51324
rect 55692 51214 55694 51266
rect 55746 51214 55748 51266
rect 55580 18564 55636 18574
rect 55580 18470 55636 18508
rect 55692 17778 55748 51214
rect 56140 43708 56196 51884
rect 56252 51604 56308 52444
rect 56364 52050 56420 55022
rect 56588 54738 56644 55244
rect 56924 55188 56980 55198
rect 56924 55094 56980 55132
rect 56588 54686 56590 54738
rect 56642 54686 56644 54738
rect 56588 54674 56644 54686
rect 56700 54628 56756 54638
rect 56700 54534 56756 54572
rect 56476 53954 56532 53966
rect 56476 53902 56478 53954
rect 56530 53902 56532 53954
rect 56476 53842 56532 53902
rect 56476 53790 56478 53842
rect 56530 53790 56532 53842
rect 56476 53778 56532 53790
rect 57036 53618 57092 53630
rect 57036 53566 57038 53618
rect 57090 53566 57092 53618
rect 56700 52836 56756 52846
rect 56700 52834 56980 52836
rect 56700 52782 56702 52834
rect 56754 52782 56980 52834
rect 56700 52780 56980 52782
rect 56700 52770 56756 52780
rect 56364 51998 56366 52050
rect 56418 51998 56420 52050
rect 56364 51986 56420 51998
rect 56924 52050 56980 52780
rect 56924 51998 56926 52050
rect 56978 51998 56980 52050
rect 56252 51538 56308 51548
rect 56588 51492 56644 51502
rect 56252 51380 56308 51418
rect 56588 51398 56644 51436
rect 56252 51314 56308 51324
rect 56924 51380 56980 51998
rect 57036 51604 57092 53566
rect 57148 52052 57204 55412
rect 57372 55300 57428 56590
rect 57484 56642 57540 56654
rect 57484 56590 57486 56642
rect 57538 56590 57540 56642
rect 57484 55522 57540 56590
rect 57484 55470 57486 55522
rect 57538 55470 57540 55522
rect 57484 55458 57540 55470
rect 57596 56308 57652 56318
rect 57708 56308 57764 57820
rect 57820 57810 57876 57820
rect 58044 57652 58100 57690
rect 58044 57586 58100 57596
rect 57932 57538 57988 57550
rect 57932 57486 57934 57538
rect 57986 57486 57988 57538
rect 57820 56980 57876 56990
rect 57820 56886 57876 56924
rect 57596 56306 57764 56308
rect 57596 56254 57598 56306
rect 57650 56254 57764 56306
rect 57596 56252 57764 56254
rect 57820 56308 57876 56318
rect 57596 55300 57652 56252
rect 57820 56214 57876 56252
rect 57820 56084 57876 56094
rect 57708 55972 57764 55982
rect 57708 55878 57764 55916
rect 57372 55244 57652 55300
rect 57708 55522 57764 55534
rect 57708 55470 57710 55522
rect 57762 55470 57764 55522
rect 57260 55188 57316 55198
rect 57260 55094 57316 55132
rect 57372 54852 57428 55244
rect 57260 54796 57428 54852
rect 57260 53620 57316 54796
rect 57372 54628 57428 54638
rect 57372 54534 57428 54572
rect 57596 53956 57652 53966
rect 57372 53620 57428 53630
rect 57260 53618 57428 53620
rect 57260 53566 57374 53618
rect 57426 53566 57428 53618
rect 57260 53564 57428 53566
rect 57372 53554 57428 53564
rect 57596 53058 57652 53900
rect 57596 53006 57598 53058
rect 57650 53006 57652 53058
rect 57596 52994 57652 53006
rect 57484 52722 57540 52734
rect 57484 52670 57486 52722
rect 57538 52670 57540 52722
rect 57484 52612 57540 52670
rect 57484 52546 57540 52556
rect 57260 52052 57316 52062
rect 57148 52050 57316 52052
rect 57148 51998 57262 52050
rect 57314 51998 57316 52050
rect 57148 51996 57316 51998
rect 57260 51986 57316 51996
rect 57036 51538 57092 51548
rect 56924 51314 56980 51324
rect 56924 49588 56980 49598
rect 56140 43652 56308 43708
rect 56252 18674 56308 43652
rect 56252 18622 56254 18674
rect 56306 18622 56308 18674
rect 56252 18610 56308 18622
rect 55804 18450 55860 18462
rect 55804 18398 55806 18450
rect 55858 18398 55860 18450
rect 55804 18340 55860 18398
rect 55804 18274 55860 18284
rect 56028 18450 56084 18462
rect 56028 18398 56030 18450
rect 56082 18398 56084 18450
rect 55692 17726 55694 17778
rect 55746 17726 55748 17778
rect 55692 17714 55748 17726
rect 55580 17668 55636 17678
rect 55580 17574 55636 17612
rect 55356 17444 55412 17454
rect 55356 16884 55412 17388
rect 56028 17444 56084 18398
rect 56252 18450 56308 18462
rect 56252 18398 56254 18450
rect 56306 18398 56308 18450
rect 56252 17890 56308 18398
rect 56252 17838 56254 17890
rect 56306 17838 56308 17890
rect 56252 17826 56308 17838
rect 56140 17668 56196 17678
rect 56140 17574 56196 17612
rect 56700 17668 56756 17678
rect 56028 17378 56084 17388
rect 56700 17442 56756 17612
rect 56700 17390 56702 17442
rect 56754 17390 56756 17442
rect 55356 16818 55412 16828
rect 56364 15428 56420 15438
rect 56364 15334 56420 15372
rect 56028 15316 56084 15326
rect 56028 15222 56084 15260
rect 55356 15204 55412 15214
rect 55468 15204 55524 15214
rect 55412 15202 55524 15204
rect 55412 15150 55470 15202
rect 55522 15150 55524 15202
rect 55412 15148 55524 15150
rect 55356 14754 55412 15148
rect 55468 15138 55524 15148
rect 55356 14702 55358 14754
rect 55410 14702 55412 14754
rect 55356 14690 55412 14702
rect 56140 14532 56196 14542
rect 56140 14438 56196 14476
rect 56364 14308 56420 14318
rect 56364 14214 56420 14252
rect 55692 13860 55748 13870
rect 55692 13766 55748 13804
rect 55356 13748 55412 13758
rect 55356 13654 55412 13692
rect 56700 13634 56756 17390
rect 56812 14532 56868 14542
rect 56812 14438 56868 14476
rect 56700 13582 56702 13634
rect 56754 13582 56756 13634
rect 56700 13524 56756 13582
rect 56700 13458 56756 13468
rect 55804 6468 55860 6478
rect 55020 6130 55300 6132
rect 55020 6078 55022 6130
rect 55074 6078 55300 6130
rect 55020 6076 55300 6078
rect 55020 6066 55076 6076
rect 54460 5070 54462 5122
rect 54514 5070 54516 5122
rect 54460 5058 54516 5070
rect 55020 5236 55076 5246
rect 54236 4844 54628 4900
rect 53340 4286 53342 4338
rect 53394 4286 53396 4338
rect 53340 4274 53396 4286
rect 53676 4228 53732 4238
rect 53564 3668 53620 3678
rect 53564 3574 53620 3612
rect 53676 800 53732 4172
rect 54012 4226 54068 4238
rect 54012 4174 54014 4226
rect 54066 4174 54068 4226
rect 54012 3556 54068 4174
rect 54012 3490 54068 3500
rect 54348 3668 54404 3678
rect 54348 800 54404 3612
rect 54572 3554 54628 4844
rect 54572 3502 54574 3554
rect 54626 3502 54628 3554
rect 54572 3490 54628 3502
rect 55020 800 55076 5180
rect 55244 5122 55300 6076
rect 55356 6356 55412 6366
rect 55356 6130 55412 6300
rect 55356 6078 55358 6130
rect 55410 6078 55412 6130
rect 55356 6066 55412 6078
rect 55244 5070 55246 5122
rect 55298 5070 55300 5122
rect 55244 5058 55300 5070
rect 55804 5794 55860 6412
rect 56924 6244 56980 49532
rect 57484 13746 57540 13758
rect 57484 13694 57486 13746
rect 57538 13694 57540 13746
rect 57484 13524 57540 13694
rect 57484 13458 57540 13468
rect 56924 6178 56980 6188
rect 57372 6356 57428 6366
rect 57372 6132 57428 6300
rect 57708 6356 57764 55470
rect 57820 55410 57876 56028
rect 57820 55358 57822 55410
rect 57874 55358 57876 55410
rect 57820 55346 57876 55358
rect 57820 13858 57876 13870
rect 57820 13806 57822 13858
rect 57874 13806 57876 13858
rect 57820 13748 57876 13806
rect 57820 13682 57876 13692
rect 57932 6692 57988 57486
rect 58044 57428 58100 57438
rect 58044 57090 58100 57372
rect 58044 57038 58046 57090
rect 58098 57038 58100 57090
rect 58044 57026 58100 57038
rect 58044 56868 58100 56878
rect 58044 56082 58100 56812
rect 58044 56030 58046 56082
rect 58098 56030 58100 56082
rect 58044 55188 58100 56030
rect 58044 55122 58100 55132
rect 58044 53956 58100 53966
rect 58044 53170 58100 53900
rect 58044 53118 58046 53170
rect 58098 53118 58100 53170
rect 58044 53106 58100 53118
rect 58156 8428 58212 58156
rect 58268 57650 58324 58382
rect 59276 58322 59332 58334
rect 59276 58270 59278 58322
rect 59330 58270 59332 58322
rect 59164 58210 59220 58222
rect 59164 58158 59166 58210
rect 59218 58158 59220 58210
rect 58268 57598 58270 57650
rect 58322 57598 58324 57650
rect 58268 56980 58324 57598
rect 58492 57652 58548 57662
rect 58492 57558 58548 57596
rect 59164 57652 59220 58158
rect 59276 58212 59332 58270
rect 59276 58146 59332 58156
rect 59164 57586 59220 57596
rect 58268 56914 58324 56924
rect 58940 56756 58996 56766
rect 58940 56662 58996 56700
rect 59500 56756 59556 56766
rect 59500 56662 59556 56700
rect 58828 56642 58884 56654
rect 58828 56590 58830 56642
rect 58882 56590 58884 56642
rect 58268 56084 58324 56094
rect 58268 55990 58324 56028
rect 58828 56084 58884 56590
rect 58828 56018 58884 56028
rect 57932 6626 57988 6636
rect 58044 8372 58212 8428
rect 58604 55972 58660 55982
rect 58044 6468 58100 8372
rect 58044 6402 58100 6412
rect 57708 6290 57764 6300
rect 58156 6244 58212 6254
rect 58156 6132 58212 6188
rect 58604 6132 58660 55916
rect 59276 52276 59332 52286
rect 59276 52182 59332 52220
rect 59388 52164 59444 52174
rect 59388 52070 59444 52108
rect 59164 6468 59220 6478
rect 58716 6132 58772 6142
rect 57372 6130 57540 6132
rect 57372 6078 57374 6130
rect 57426 6078 57540 6130
rect 57372 6076 57540 6078
rect 57372 6066 57428 6076
rect 55804 5742 55806 5794
rect 55858 5742 55860 5794
rect 55804 4340 55860 5742
rect 56364 6020 56420 6030
rect 56364 5796 56420 5964
rect 56364 5794 56532 5796
rect 56364 5742 56366 5794
rect 56418 5742 56532 5794
rect 56364 5740 56532 5742
rect 56364 5730 56420 5740
rect 55916 5236 55972 5246
rect 55916 5142 55972 5180
rect 56140 4340 56196 4350
rect 55804 4338 56196 4340
rect 55804 4286 56142 4338
rect 56194 4286 56196 4338
rect 55804 4284 56196 4286
rect 56140 4274 56196 4284
rect 55468 4228 55524 4238
rect 55468 4134 55524 4172
rect 55804 3556 55860 3566
rect 56476 3556 56532 5740
rect 57372 5124 57428 5134
rect 57036 5122 57428 5124
rect 57036 5070 57374 5122
rect 57426 5070 57428 5122
rect 57036 5068 57428 5070
rect 56700 3556 56756 3566
rect 56476 3554 56756 3556
rect 56476 3502 56702 3554
rect 56754 3502 56756 3554
rect 56476 3500 56756 3502
rect 55692 3444 55748 3454
rect 55692 3350 55748 3388
rect 55804 2100 55860 3500
rect 56700 3490 56756 3500
rect 55692 2044 55860 2100
rect 56364 3444 56420 3454
rect 55692 800 55748 2044
rect 56364 800 56420 3388
rect 57036 800 57092 5068
rect 57372 5058 57428 5068
rect 57484 4338 57540 6076
rect 58156 6130 58436 6132
rect 58156 6078 58158 6130
rect 58210 6078 58436 6130
rect 58156 6076 58436 6078
rect 58156 6066 58212 6076
rect 58380 4900 58436 6076
rect 58604 6130 58772 6132
rect 58604 6078 58718 6130
rect 58770 6078 58772 6130
rect 58604 6076 58772 6078
rect 58492 5124 58548 5134
rect 58604 5124 58660 6076
rect 58716 6066 58772 6076
rect 59164 6130 59220 6412
rect 59612 6356 59668 6366
rect 59612 6132 59668 6300
rect 59724 6244 59780 59054
rect 59836 58212 59892 58222
rect 59836 58118 59892 58156
rect 59948 55468 60004 59276
rect 60284 59218 60340 59724
rect 60284 59166 60286 59218
rect 60338 59166 60340 59218
rect 60284 59154 60340 59166
rect 60060 59106 60116 59118
rect 60060 59054 60062 59106
rect 60114 59054 60116 59106
rect 60060 58996 60116 59054
rect 60396 58996 60452 60062
rect 60844 60674 60900 60686
rect 60844 60622 60846 60674
rect 60898 60622 60900 60674
rect 60620 60004 60676 60014
rect 60620 59910 60676 59948
rect 60060 58940 60452 58996
rect 60844 55468 60900 60622
rect 61068 60116 61124 60844
rect 61964 60786 62020 61292
rect 62188 61254 62244 61292
rect 62748 61346 62804 61358
rect 62748 61294 62750 61346
rect 62802 61294 62804 61346
rect 62412 61012 62468 61022
rect 62412 60918 62468 60956
rect 62636 60900 62692 60910
rect 62636 60806 62692 60844
rect 61964 60734 61966 60786
rect 62018 60734 62020 60786
rect 61964 60722 62020 60734
rect 61180 60676 61236 60686
rect 61180 60582 61236 60620
rect 62188 60676 62244 60686
rect 62188 60582 62244 60620
rect 62524 60676 62580 60686
rect 62524 60582 62580 60620
rect 61404 60564 61460 60574
rect 61404 60470 61460 60508
rect 61068 59442 61124 60060
rect 62748 60452 62804 61294
rect 61516 59892 61572 59902
rect 61516 59798 61572 59836
rect 62076 59892 62132 59902
rect 62076 59798 62132 59836
rect 61404 59780 61460 59790
rect 61404 59686 61460 59724
rect 61068 59390 61070 59442
rect 61122 59390 61124 59442
rect 61068 59378 61124 59390
rect 61292 59218 61348 59230
rect 61292 59166 61294 59218
rect 61346 59166 61348 59218
rect 61292 59108 61348 59166
rect 61292 59042 61348 59052
rect 61852 59108 61908 59118
rect 61852 59014 61908 59052
rect 62748 59108 62804 60396
rect 62748 59042 62804 59052
rect 62860 58100 62916 62190
rect 63196 61348 63252 62524
rect 63308 62914 63364 62926
rect 63308 62862 63310 62914
rect 63362 62862 63364 62914
rect 63308 61572 63364 62862
rect 63420 62916 63476 62926
rect 63420 62822 63476 62860
rect 63532 61796 63588 63084
rect 63532 61730 63588 61740
rect 63644 62916 63700 62926
rect 63308 61516 63588 61572
rect 63308 61348 63364 61358
rect 63196 61346 63364 61348
rect 63196 61294 63310 61346
rect 63362 61294 63364 61346
rect 63196 61292 63364 61294
rect 63308 61282 63364 61292
rect 63196 60676 63252 60686
rect 62860 58044 63028 58100
rect 62860 57764 62916 57774
rect 62860 57670 62916 57708
rect 62748 57428 62804 57438
rect 62748 57334 62804 57372
rect 59948 55412 60116 55468
rect 60844 55412 61684 55468
rect 59948 52164 60004 52174
rect 59948 52070 60004 52108
rect 60060 6356 60116 55412
rect 61404 53844 61460 53854
rect 60508 52500 60564 52510
rect 60508 52386 60564 52444
rect 60508 52334 60510 52386
rect 60562 52334 60564 52386
rect 60508 52322 60564 52334
rect 60620 52276 60676 52286
rect 61404 52276 61460 53788
rect 60620 52274 61460 52276
rect 60620 52222 60622 52274
rect 60674 52222 61406 52274
rect 61458 52222 61460 52274
rect 60620 52220 61460 52222
rect 60620 52210 60676 52220
rect 61404 52210 61460 52220
rect 61628 8428 61684 55412
rect 62972 31948 63028 58044
rect 61180 8372 61684 8428
rect 62860 31892 63028 31948
rect 60060 6290 60116 6300
rect 60284 6692 60340 6702
rect 59724 6178 59780 6188
rect 59164 6078 59166 6130
rect 59218 6078 59220 6130
rect 58492 5122 58660 5124
rect 58492 5070 58494 5122
rect 58546 5070 58660 5122
rect 58492 5068 58660 5070
rect 59164 5124 59220 6078
rect 59388 6130 59668 6132
rect 59388 6078 59614 6130
rect 59666 6078 59668 6130
rect 59388 6076 59668 6078
rect 59276 5124 59332 5134
rect 59164 5122 59332 5124
rect 59164 5070 59278 5122
rect 59330 5070 59332 5122
rect 59164 5068 59332 5070
rect 58492 5058 58548 5068
rect 59276 5058 59332 5068
rect 58380 4844 58548 4900
rect 57484 4286 57486 4338
rect 57538 4286 57540 4338
rect 57484 4274 57540 4286
rect 57708 4228 57764 4238
rect 57372 3668 57428 3678
rect 57372 3574 57428 3612
rect 57708 800 57764 4172
rect 58156 4226 58212 4238
rect 58156 4174 58158 4226
rect 58210 4174 58212 4226
rect 58156 3556 58212 4174
rect 58156 3490 58212 3500
rect 58380 3556 58436 3566
rect 58380 800 58436 3500
rect 58492 3554 58548 4844
rect 59388 4338 59444 6076
rect 59612 6066 59668 6076
rect 60284 6132 60340 6636
rect 61068 6244 61124 6254
rect 60284 6130 60676 6132
rect 60284 6078 60286 6130
rect 60338 6078 60676 6130
rect 60284 6076 60676 6078
rect 60284 6066 60340 6076
rect 59948 5236 60004 5246
rect 59388 4286 59390 4338
rect 59442 4286 59444 4338
rect 59388 4274 59444 4286
rect 59500 5234 60004 5236
rect 59500 5182 59950 5234
rect 60002 5182 60004 5234
rect 59500 5180 60004 5182
rect 58492 3502 58494 3554
rect 58546 3502 58548 3554
rect 58492 3490 58548 3502
rect 59164 3666 59220 3678
rect 59164 3614 59166 3666
rect 59218 3614 59220 3666
rect 59164 3444 59220 3614
rect 59164 3378 59220 3388
rect 59500 980 59556 5180
rect 59948 5170 60004 5180
rect 59948 4228 60004 4238
rect 59948 4134 60004 4172
rect 59052 924 59556 980
rect 59724 3780 59780 3790
rect 59052 800 59108 924
rect 59724 800 59780 3724
rect 60396 3668 60452 3678
rect 60396 800 60452 3612
rect 60620 3554 60676 6076
rect 60620 3502 60622 3554
rect 60674 3502 60676 3554
rect 60620 3490 60676 3502
rect 60956 5236 61012 5246
rect 60956 2548 61012 5180
rect 61068 4338 61124 6188
rect 61180 6130 61236 8372
rect 62076 6356 62132 6366
rect 61180 6078 61182 6130
rect 61234 6078 61236 6130
rect 61180 5124 61236 6078
rect 61516 6244 61572 6254
rect 61516 6130 61572 6188
rect 61516 6078 61518 6130
rect 61570 6078 61572 6130
rect 61516 6066 61572 6078
rect 62076 6132 62132 6300
rect 62860 6244 62916 31892
rect 62860 6178 62916 6188
rect 62076 6130 62468 6132
rect 62076 6078 62078 6130
rect 62130 6078 62468 6130
rect 62076 6076 62468 6078
rect 62076 6066 62132 6076
rect 62076 5236 62132 5246
rect 62076 5142 62132 5180
rect 61404 5124 61460 5134
rect 61180 5122 61460 5124
rect 61180 5070 61406 5122
rect 61458 5070 61460 5122
rect 61180 5068 61460 5070
rect 61404 5058 61460 5068
rect 61068 4286 61070 4338
rect 61122 4286 61124 4338
rect 61068 4274 61124 4286
rect 61740 4226 61796 4238
rect 61740 4174 61742 4226
rect 61794 4174 61796 4226
rect 61740 3780 61796 4174
rect 61740 3714 61796 3724
rect 61852 4228 61908 4238
rect 61292 3666 61348 3678
rect 61292 3614 61294 3666
rect 61346 3614 61348 3666
rect 61292 3556 61348 3614
rect 61292 3490 61348 3500
rect 60956 2492 61124 2548
rect 61068 800 61124 2492
rect 61852 2100 61908 4172
rect 62412 3554 62468 6076
rect 63196 4340 63252 60620
rect 63308 60116 63364 60126
rect 63308 57874 63364 60060
rect 63308 57822 63310 57874
rect 63362 57822 63364 57874
rect 63308 57764 63364 57822
rect 63308 57698 63364 57708
rect 63532 6356 63588 61516
rect 63644 61458 63700 62860
rect 63756 62580 63812 62590
rect 63756 62486 63812 62524
rect 63980 62356 64036 62366
rect 63980 62262 64036 62300
rect 64092 62354 64148 63084
rect 64092 62302 64094 62354
rect 64146 62302 64148 62354
rect 64092 62290 64148 62302
rect 63868 62242 63924 62254
rect 63868 62190 63870 62242
rect 63922 62190 63924 62242
rect 63644 61406 63646 61458
rect 63698 61406 63700 61458
rect 63644 60452 63700 61406
rect 63644 60386 63700 60396
rect 63756 61684 63812 61694
rect 63532 6290 63588 6300
rect 63420 5012 63476 5022
rect 63196 4274 63252 4284
rect 63308 5010 63476 5012
rect 63308 4958 63422 5010
rect 63474 4958 63476 5010
rect 63308 4956 63476 4958
rect 62972 4228 63028 4238
rect 62972 4134 63028 4172
rect 63084 3668 63140 3678
rect 63084 3574 63140 3612
rect 62412 3502 62414 3554
rect 62466 3502 62468 3554
rect 62412 3490 62468 3502
rect 62524 3556 62580 3566
rect 61740 2044 61908 2100
rect 61740 800 61796 2044
rect 62524 1764 62580 3500
rect 62412 1708 62580 1764
rect 62412 800 62468 1708
rect 63308 980 63364 4956
rect 63420 4946 63476 4956
rect 63756 4452 63812 61628
rect 63868 55468 63924 62190
rect 64428 62244 64484 62282
rect 64428 62178 64484 62188
rect 64540 60676 64596 60686
rect 64540 60582 64596 60620
rect 64428 60564 64484 60574
rect 64428 60470 64484 60508
rect 65212 55468 65268 64430
rect 65324 64484 65380 64494
rect 65324 64390 65380 64428
rect 65436 64148 65492 64654
rect 65436 64082 65492 64092
rect 65548 64596 65604 64606
rect 65324 63924 65380 63934
rect 65548 63924 65604 64540
rect 65380 63922 65604 63924
rect 65380 63870 65550 63922
rect 65602 63870 65604 63922
rect 65380 63868 65604 63870
rect 65324 63250 65380 63868
rect 65548 63858 65604 63868
rect 65324 63198 65326 63250
rect 65378 63198 65380 63250
rect 65324 63186 65380 63198
rect 65660 62188 65716 64876
rect 65772 64866 65828 64876
rect 66444 64818 66500 64988
rect 66444 64766 66446 64818
rect 66498 64766 66500 64818
rect 66444 64754 66500 64766
rect 65772 64708 65828 64718
rect 66332 64708 66388 64718
rect 65772 64706 66388 64708
rect 65772 64654 65774 64706
rect 65826 64654 66334 64706
rect 66386 64654 66388 64706
rect 65772 64652 66388 64654
rect 65772 64642 65828 64652
rect 66332 64642 66388 64652
rect 66332 64260 66388 64270
rect 65772 64148 65828 64158
rect 65772 64054 65828 64092
rect 66332 64146 66388 64204
rect 66332 64094 66334 64146
rect 66386 64094 66388 64146
rect 66332 64082 66388 64094
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 65996 62916 66052 62926
rect 65996 62822 66052 62860
rect 66556 62188 66612 65212
rect 66668 64260 66724 65436
rect 66780 65380 66836 65390
rect 66780 65378 66948 65380
rect 66780 65326 66782 65378
rect 66834 65326 66948 65378
rect 66780 65324 66948 65326
rect 66780 65314 66836 65324
rect 66892 64596 66948 65324
rect 67004 64820 67060 66220
rect 67116 65378 67172 65390
rect 67116 65326 67118 65378
rect 67170 65326 67172 65378
rect 67116 65156 67172 65326
rect 67116 65090 67172 65100
rect 67004 64764 67172 64820
rect 67004 64596 67060 64606
rect 66948 64594 67060 64596
rect 66948 64542 67006 64594
rect 67058 64542 67060 64594
rect 66948 64540 67060 64542
rect 66892 64464 66948 64540
rect 67004 64530 67060 64540
rect 66668 64194 66724 64204
rect 66668 63924 66724 63934
rect 66668 62916 66724 63868
rect 66668 62850 66724 62860
rect 67004 62916 67060 62926
rect 67004 62822 67060 62860
rect 65660 62132 66388 62188
rect 66556 62132 66948 62188
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 65324 60676 65380 60686
rect 65324 60582 65380 60620
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 66332 55468 66388 62132
rect 66556 60228 66612 60238
rect 66556 60114 66612 60172
rect 66556 60062 66558 60114
rect 66610 60062 66612 60114
rect 66556 60050 66612 60062
rect 66444 60004 66500 60014
rect 66444 59910 66500 59948
rect 63868 55412 64708 55468
rect 65212 55412 65492 55468
rect 66332 55412 66612 55468
rect 64652 20188 64708 55412
rect 64652 20132 65380 20188
rect 64204 6244 64260 6254
rect 64204 6132 64260 6188
rect 64204 6130 64484 6132
rect 64204 6078 64206 6130
rect 64258 6078 64484 6130
rect 64204 6076 64484 6078
rect 64204 6066 64260 6076
rect 63756 4386 63812 4396
rect 63868 4340 63924 4350
rect 63868 4246 63924 4284
rect 63084 924 63364 980
rect 63756 4116 63812 4126
rect 64428 4116 64484 6076
rect 65324 6130 65380 20132
rect 65436 6244 65492 55412
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 66556 43708 66612 55412
rect 66668 49140 66724 49150
rect 66668 49046 66724 49084
rect 66556 43652 66724 43708
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 66668 6580 66724 43652
rect 66780 6580 66836 6590
rect 66668 6578 66836 6580
rect 66668 6526 66782 6578
rect 66834 6526 66836 6578
rect 66668 6524 66836 6526
rect 66780 6468 66836 6524
rect 66780 6402 66836 6412
rect 65436 6178 65492 6188
rect 65772 6356 65828 6366
rect 65772 6132 65828 6300
rect 65324 6078 65326 6130
rect 65378 6078 65380 6130
rect 64540 5124 64596 5134
rect 65324 5124 65380 6078
rect 64540 5122 65380 5124
rect 64540 5070 64542 5122
rect 64594 5070 65380 5122
rect 64540 5068 65380 5070
rect 65660 6130 65828 6132
rect 65660 6078 65774 6130
rect 65826 6078 65828 6130
rect 65660 6076 65828 6078
rect 64540 5058 64596 5068
rect 65436 5012 65492 5022
rect 65100 5010 65492 5012
rect 65100 4958 65438 5010
rect 65490 4958 65492 5010
rect 65100 4956 65492 4958
rect 64540 4340 64596 4350
rect 64540 4246 64596 4284
rect 64428 4060 64596 4116
rect 63084 800 63140 924
rect 63756 800 63812 4060
rect 64540 3554 64596 4060
rect 64540 3502 64542 3554
rect 64594 3502 64596 3554
rect 64540 3490 64596 3502
rect 64428 3444 64484 3454
rect 64428 800 64484 3388
rect 65100 800 65156 4956
rect 65436 4946 65492 4956
rect 65660 4338 65716 6076
rect 65772 6066 65828 6076
rect 66332 6244 66388 6254
rect 66332 6130 66388 6188
rect 66332 6078 66334 6130
rect 66386 6078 66388 6130
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 66332 5122 66388 6078
rect 66780 6244 66836 6254
rect 66780 6130 66836 6188
rect 66780 6078 66782 6130
rect 66834 6078 66836 6130
rect 66780 6066 66836 6078
rect 66332 5070 66334 5122
rect 66386 5070 66388 5122
rect 66332 5058 66388 5070
rect 66556 5236 66612 5246
rect 65660 4286 65662 4338
rect 65714 4286 65716 4338
rect 65660 4274 65716 4286
rect 65772 4228 65828 4238
rect 65212 3666 65268 3678
rect 65212 3614 65214 3666
rect 65266 3614 65268 3666
rect 65212 3556 65268 3614
rect 65212 3490 65268 3500
rect 65772 800 65828 4172
rect 66108 4226 66164 4238
rect 66108 4174 66110 4226
rect 66162 4174 66164 4226
rect 66108 4116 66164 4174
rect 66108 4050 66164 4060
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 66444 3444 66500 3454
rect 66444 3350 66500 3388
rect 66556 2660 66612 5180
rect 66892 4340 66948 62132
rect 67116 61236 67172 64764
rect 67340 64596 67396 64606
rect 67340 64502 67396 64540
rect 67340 63924 67396 63934
rect 67340 63830 67396 63868
rect 67004 61180 67172 61236
rect 67004 6244 67060 61180
rect 67116 60228 67172 60238
rect 67116 60114 67172 60172
rect 67116 60062 67118 60114
rect 67170 60062 67172 60114
rect 67116 60050 67172 60062
rect 67564 55468 67620 66892
rect 67676 66050 67732 67004
rect 67788 66276 67844 67564
rect 68012 67554 68068 67564
rect 68348 67282 68404 68348
rect 68460 68180 68516 68190
rect 68460 67954 68516 68124
rect 68460 67902 68462 67954
rect 68514 67902 68516 67954
rect 68460 67890 68516 67902
rect 68348 67230 68350 67282
rect 68402 67230 68404 67282
rect 68348 67218 68404 67230
rect 68124 67060 68180 67070
rect 68124 66966 68180 67004
rect 68460 67058 68516 67070
rect 68460 67006 68462 67058
rect 68514 67006 68516 67058
rect 68236 66948 68292 66958
rect 68236 66854 68292 66892
rect 67788 66210 67844 66220
rect 67900 66834 67956 66846
rect 67900 66782 67902 66834
rect 67954 66782 67956 66834
rect 67900 66274 67956 66782
rect 68460 66724 68516 67006
rect 68124 66668 68516 66724
rect 68124 66386 68180 66668
rect 68348 66500 68404 66510
rect 68348 66406 68404 66444
rect 68124 66334 68126 66386
rect 68178 66334 68180 66386
rect 68124 66322 68180 66334
rect 67900 66222 67902 66274
rect 67954 66222 67956 66274
rect 67900 66210 67956 66222
rect 68236 66276 68292 66286
rect 67676 65998 67678 66050
rect 67730 65998 67732 66050
rect 67676 65492 67732 65998
rect 67676 65426 67732 65436
rect 67788 66050 67844 66062
rect 67788 65998 67790 66050
rect 67842 65998 67844 66050
rect 67676 64148 67732 64158
rect 67676 64054 67732 64092
rect 67564 55412 67732 55468
rect 67116 49140 67172 49150
rect 67116 49046 67172 49084
rect 67228 48804 67284 48814
rect 67228 48710 67284 48748
rect 67676 6692 67732 55412
rect 67676 6626 67732 6636
rect 67004 6178 67060 6188
rect 67116 6468 67172 6478
rect 67116 5122 67172 6412
rect 67340 6244 67396 6254
rect 67340 5906 67396 6188
rect 67340 5854 67342 5906
rect 67394 5854 67396 5906
rect 67340 5842 67396 5854
rect 67116 5070 67118 5122
rect 67170 5070 67172 5122
rect 67116 5058 67172 5070
rect 67228 5796 67284 5806
rect 67228 4900 67284 5740
rect 67788 5572 67844 65998
rect 68236 65714 68292 66220
rect 68236 65662 68238 65714
rect 68290 65662 68292 65714
rect 68236 65650 68292 65662
rect 68012 65492 68068 65502
rect 68012 64148 68068 65436
rect 68460 65490 68516 66668
rect 68460 65438 68462 65490
rect 68514 65438 68516 65490
rect 68124 65380 68180 65390
rect 68124 65286 68180 65324
rect 68012 64082 68068 64092
rect 68124 65044 68180 65054
rect 68124 62468 68180 64988
rect 68236 64708 68292 64718
rect 68460 64708 68516 65438
rect 68236 64706 68516 64708
rect 68236 64654 68238 64706
rect 68290 64654 68516 64706
rect 68236 64652 68516 64654
rect 68236 64596 68292 64652
rect 68236 64530 68292 64540
rect 68572 64482 68628 68348
rect 68684 68402 68740 68414
rect 68684 68350 68686 68402
rect 68738 68350 68740 68402
rect 68684 67060 68740 68350
rect 68796 67060 68852 67070
rect 68684 67058 68852 67060
rect 68684 67006 68798 67058
rect 68850 67006 68852 67058
rect 68684 67004 68852 67006
rect 68796 66994 68852 67004
rect 68684 65604 68740 65614
rect 68684 65490 68740 65548
rect 68684 65438 68686 65490
rect 68738 65438 68740 65490
rect 68684 65426 68740 65438
rect 68572 64430 68574 64482
rect 68626 64430 68628 64482
rect 68572 64372 68628 64430
rect 68348 64316 68628 64372
rect 68796 65380 68852 65390
rect 69132 65380 69188 72380
rect 69356 72304 69412 72380
rect 69692 72436 69748 73166
rect 71820 73220 71876 73230
rect 69692 72370 69748 72380
rect 70140 72436 70196 72446
rect 70140 72342 70196 72380
rect 71820 72434 71876 73164
rect 72380 73218 72436 73230
rect 72380 73166 72382 73218
rect 72434 73166 72436 73218
rect 72156 72548 72212 72558
rect 72156 72454 72212 72492
rect 72380 72548 72436 73166
rect 72380 72482 72436 72492
rect 71820 72382 71822 72434
rect 71874 72382 71876 72434
rect 71820 72370 71876 72382
rect 69468 72324 69524 72334
rect 69468 72230 69524 72268
rect 69580 72322 69636 72334
rect 69580 72270 69582 72322
rect 69634 72270 69636 72322
rect 69580 71988 69636 72270
rect 69580 71922 69636 71932
rect 72492 71986 72548 73276
rect 73052 72548 73108 72558
rect 73500 72548 73556 73836
rect 73612 73826 73668 73836
rect 73724 73554 73780 75068
rect 74956 75124 75012 75630
rect 74956 75058 75012 75068
rect 74956 74900 75012 74910
rect 74732 74898 75012 74900
rect 74732 74846 74958 74898
rect 75010 74846 75012 74898
rect 74732 74844 75012 74846
rect 73724 73502 73726 73554
rect 73778 73502 73780 73554
rect 73724 73490 73780 73502
rect 74060 73890 74116 73902
rect 74060 73838 74062 73890
rect 74114 73838 74116 73890
rect 73836 73444 73892 73454
rect 73612 73108 73668 73118
rect 73612 72660 73668 73052
rect 73612 72594 73668 72604
rect 73108 72492 73220 72548
rect 73052 72416 73108 72492
rect 72492 71934 72494 71986
rect 72546 71934 72548 71986
rect 72492 71922 72548 71934
rect 71260 71876 71316 71886
rect 71260 71782 71316 71820
rect 71596 71876 71652 71886
rect 71596 71782 71652 71820
rect 72268 71876 72324 71886
rect 70812 71764 70868 71774
rect 70812 71670 70868 71708
rect 71932 71764 71988 71774
rect 70588 71652 70644 71662
rect 70140 70868 70196 70878
rect 70140 70774 70196 70812
rect 70588 70866 70644 71596
rect 70588 70814 70590 70866
rect 70642 70814 70644 70866
rect 70588 70802 70644 70814
rect 70700 71316 70756 71326
rect 69916 70308 69972 70318
rect 69916 70214 69972 70252
rect 69468 70196 69524 70206
rect 69468 70102 69524 70140
rect 70252 70196 70308 70206
rect 70252 70102 70308 70140
rect 69580 70084 69636 70094
rect 69356 69188 69412 69198
rect 69356 69094 69412 69132
rect 69580 68852 69636 70028
rect 69468 68796 69636 68852
rect 69692 69300 69748 69310
rect 69468 67954 69524 68796
rect 69692 68516 69748 69244
rect 70252 69300 70308 69310
rect 70252 69206 70308 69244
rect 70588 69300 70644 69310
rect 70700 69300 70756 71260
rect 70924 70868 70980 70878
rect 70924 70774 70980 70812
rect 71596 70868 71652 70878
rect 71596 70774 71652 70812
rect 71932 70866 71988 71708
rect 71932 70814 71934 70866
rect 71986 70814 71988 70866
rect 71932 70802 71988 70814
rect 72268 71762 72324 71820
rect 72268 71710 72270 71762
rect 72322 71710 72324 71762
rect 72268 70756 72324 71710
rect 72268 70690 72324 70700
rect 72380 70868 72436 70878
rect 72380 70756 72436 70812
rect 72492 70756 72548 70766
rect 72380 70754 72548 70756
rect 72380 70702 72494 70754
rect 72546 70702 72548 70754
rect 72380 70700 72548 70702
rect 71260 70644 71316 70654
rect 71260 70418 71316 70588
rect 71260 70366 71262 70418
rect 71314 70366 71316 70418
rect 71260 70354 71316 70366
rect 70588 69298 70756 69300
rect 70588 69246 70590 69298
rect 70642 69246 70756 69298
rect 70588 69244 70756 69246
rect 70924 70196 70980 70206
rect 70588 69234 70644 69244
rect 69916 68516 69972 68526
rect 69692 68514 69972 68516
rect 69692 68462 69918 68514
rect 69970 68462 69972 68514
rect 69692 68460 69972 68462
rect 69468 67902 69470 67954
rect 69522 67902 69524 67954
rect 69468 67890 69524 67902
rect 69580 68292 69636 68302
rect 69356 67620 69412 67630
rect 69244 67618 69412 67620
rect 69244 67566 69358 67618
rect 69410 67566 69412 67618
rect 69244 67564 69412 67566
rect 69244 65604 69300 67564
rect 69356 67554 69412 67564
rect 69468 67172 69524 67182
rect 69580 67172 69636 68236
rect 69468 67170 69636 67172
rect 69468 67118 69470 67170
rect 69522 67118 69636 67170
rect 69468 67116 69636 67118
rect 69468 67106 69524 67116
rect 69356 66834 69412 66846
rect 69356 66782 69358 66834
rect 69410 66782 69412 66834
rect 69356 66500 69412 66782
rect 69356 66434 69412 66444
rect 69244 65538 69300 65548
rect 69132 65324 69524 65380
rect 68236 62468 68292 62478
rect 68124 62412 68236 62468
rect 68236 62336 68292 62412
rect 68124 62244 68180 62282
rect 68124 62178 68180 62188
rect 68348 62188 68404 64316
rect 68684 62468 68740 62478
rect 68684 62374 68740 62412
rect 68348 62132 68628 62188
rect 68572 55468 68628 62132
rect 68348 55412 68628 55468
rect 68348 49138 68404 55412
rect 68348 49086 68350 49138
rect 68402 49086 68404 49138
rect 68348 48916 68404 49086
rect 68572 49028 68628 49038
rect 68572 48934 68628 48972
rect 68348 48850 68404 48860
rect 67900 48802 67956 48814
rect 67900 48750 67902 48802
rect 67954 48750 67956 48802
rect 67900 48692 67956 48750
rect 67900 48626 67956 48636
rect 68012 48802 68068 48814
rect 68012 48750 68014 48802
rect 68066 48750 68068 48802
rect 68012 43708 68068 48750
rect 68124 48804 68180 48814
rect 68124 48710 68180 48748
rect 68012 43652 68180 43708
rect 68012 5796 68068 5806
rect 68012 5702 68068 5740
rect 67788 5506 67844 5516
rect 68124 5460 68180 43652
rect 68684 6692 68740 6702
rect 68684 6598 68740 6636
rect 68796 5908 68852 65324
rect 69356 64594 69412 64606
rect 69356 64542 69358 64594
rect 69410 64542 69412 64594
rect 69356 64148 69412 64542
rect 69468 64484 69524 65324
rect 69692 64484 69748 64494
rect 69468 64482 69748 64484
rect 69468 64430 69694 64482
rect 69746 64430 69748 64482
rect 69468 64428 69748 64430
rect 69356 64082 69412 64092
rect 69692 55468 69748 64428
rect 68908 55412 69748 55468
rect 68908 48692 68964 55412
rect 69468 49140 69524 49150
rect 69468 49046 69524 49084
rect 69356 49028 69412 49038
rect 69356 48934 69412 48972
rect 68908 48466 68964 48636
rect 68908 48414 68910 48466
rect 68962 48414 68964 48466
rect 68908 48402 68964 48414
rect 69356 6692 69412 6702
rect 69356 6598 69412 6636
rect 68796 5842 68852 5852
rect 68124 5394 68180 5404
rect 69244 5794 69300 5806
rect 69244 5742 69246 5794
rect 69298 5742 69300 5794
rect 67788 5236 67844 5246
rect 67788 5142 67844 5180
rect 68012 5236 68068 5246
rect 66892 4274 66948 4284
rect 67116 4844 67284 4900
rect 66444 2604 66612 2660
rect 66444 800 66500 2604
rect 67116 800 67172 4844
rect 67452 4452 67508 4462
rect 67340 4228 67396 4238
rect 67340 4134 67396 4172
rect 67452 3668 67508 4396
rect 67452 3554 67508 3612
rect 67452 3502 67454 3554
rect 67506 3502 67508 3554
rect 67452 3490 67508 3502
rect 68012 980 68068 5180
rect 68460 5124 68516 5134
rect 68236 4340 68292 4350
rect 68236 4246 68292 4284
rect 68348 3668 68404 3678
rect 68348 3574 68404 3612
rect 67788 924 68068 980
rect 67788 800 67844 924
rect 68460 800 68516 5068
rect 69244 5124 69300 5742
rect 69244 5058 69300 5068
rect 69356 5572 69412 5582
rect 69356 5122 69412 5516
rect 69356 5070 69358 5122
rect 69410 5070 69412 5122
rect 69356 4564 69412 5070
rect 69468 4564 69524 4574
rect 69356 4562 69524 4564
rect 69356 4510 69470 4562
rect 69522 4510 69524 4562
rect 69356 4508 69524 4510
rect 69468 4498 69524 4508
rect 68908 4340 68964 4350
rect 68908 4246 68964 4284
rect 69132 3780 69188 3790
rect 69132 800 69188 3724
rect 69916 3668 69972 68460
rect 70028 48916 70084 48926
rect 70028 48822 70084 48860
rect 70028 6802 70084 6814
rect 70028 6750 70030 6802
rect 70082 6750 70084 6802
rect 70028 3780 70084 6750
rect 70140 5908 70196 5918
rect 70140 5814 70196 5852
rect 70812 5908 70868 5918
rect 70812 5814 70868 5852
rect 70140 5236 70196 5246
rect 70140 5142 70196 5180
rect 70812 4452 70868 4462
rect 70476 4450 70868 4452
rect 70476 4398 70814 4450
rect 70866 4398 70868 4450
rect 70476 4396 70868 4398
rect 70252 4228 70308 4238
rect 70476 4228 70532 4396
rect 70812 4386 70868 4396
rect 70252 4226 70532 4228
rect 70252 4174 70254 4226
rect 70306 4174 70532 4226
rect 70252 4172 70532 4174
rect 70252 4162 70308 4172
rect 70028 3714 70084 3724
rect 69916 3602 69972 3612
rect 69580 3444 69636 3454
rect 70140 3444 70196 3454
rect 69580 3442 70196 3444
rect 69580 3390 69582 3442
rect 69634 3390 70142 3442
rect 70194 3390 70196 3442
rect 69580 3388 70196 3390
rect 69580 3378 69636 3388
rect 69804 800 69860 3388
rect 70140 3378 70196 3388
rect 70476 800 70532 4172
rect 70924 4228 70980 70140
rect 71708 70196 71764 70206
rect 71708 70102 71764 70140
rect 71148 69300 71204 69310
rect 71148 69206 71204 69244
rect 72156 50708 72212 50718
rect 72156 50614 72212 50652
rect 71596 5124 71652 5134
rect 71596 5122 71876 5124
rect 71596 5070 71598 5122
rect 71650 5070 71876 5122
rect 71596 5068 71876 5070
rect 71596 5058 71652 5068
rect 70924 4162 70980 4172
rect 71820 5012 71876 5068
rect 72268 5012 72324 5022
rect 71820 5010 72324 5012
rect 71820 4958 72270 5010
rect 72322 4958 72324 5010
rect 71820 4956 72324 4958
rect 71260 3668 71316 3678
rect 71260 3574 71316 3612
rect 71148 3444 71204 3454
rect 71148 800 71204 3388
rect 71820 800 71876 4956
rect 72268 4946 72324 4956
rect 71932 4228 71988 4238
rect 71932 4134 71988 4172
rect 72380 3666 72436 70700
rect 72492 70690 72548 70700
rect 72828 70756 72884 70766
rect 72828 70662 72884 70700
rect 72940 69524 72996 69534
rect 72940 69430 72996 69468
rect 72940 64820 72996 64830
rect 72940 64726 72996 64764
rect 72940 60114 72996 60126
rect 72940 60062 72942 60114
rect 72994 60062 72996 60114
rect 72940 59892 72996 60062
rect 72940 59826 72996 59836
rect 72604 50708 72660 50718
rect 72604 50614 72660 50652
rect 72716 50370 72772 50382
rect 72716 50318 72718 50370
rect 72770 50318 72772 50370
rect 72716 50036 72772 50318
rect 72716 49970 72772 49980
rect 72604 49812 72660 49822
rect 72604 49698 72660 49756
rect 72604 49646 72606 49698
rect 72658 49646 72660 49698
rect 72604 48916 72660 49646
rect 72604 48850 72660 48860
rect 73052 48802 73108 48814
rect 73052 48750 73054 48802
rect 73106 48750 73108 48802
rect 73052 48692 73108 48750
rect 73052 48626 73108 48636
rect 72380 3614 72382 3666
rect 72434 3614 72436 3666
rect 72380 3602 72436 3614
rect 72492 4452 72548 4462
rect 72492 800 72548 4396
rect 72716 4226 72772 4238
rect 72716 4174 72718 4226
rect 72770 4174 72772 4226
rect 72716 3444 72772 4174
rect 73164 4228 73220 72492
rect 73500 72482 73556 72492
rect 73276 72436 73332 72446
rect 73276 72342 73332 72380
rect 73836 72324 73892 73388
rect 74060 73332 74116 73838
rect 74060 73276 74340 73332
rect 74284 73220 74340 73276
rect 74396 73220 74452 73230
rect 74284 73218 74452 73220
rect 74284 73166 74398 73218
rect 74450 73166 74452 73218
rect 74284 73164 74452 73166
rect 74172 73108 74228 73118
rect 74060 73106 74228 73108
rect 74060 73054 74174 73106
rect 74226 73054 74228 73106
rect 74060 73052 74228 73054
rect 74060 72658 74116 73052
rect 74172 73042 74228 73052
rect 74060 72606 74062 72658
rect 74114 72606 74116 72658
rect 74060 72594 74116 72606
rect 74172 72660 74228 72670
rect 74396 72660 74452 73164
rect 74732 73106 74788 74844
rect 74956 74834 75012 74844
rect 75516 74564 75572 75740
rect 75628 75730 75684 75740
rect 75516 74498 75572 74508
rect 75628 74786 75684 74798
rect 75628 74734 75630 74786
rect 75682 74734 75684 74786
rect 74956 74228 75012 74238
rect 74732 73054 74734 73106
rect 74786 73054 74788 73106
rect 74732 73042 74788 73054
rect 74844 74226 75012 74228
rect 74844 74174 74958 74226
rect 75010 74174 75012 74226
rect 74844 74172 75012 74174
rect 74228 72604 74452 72660
rect 74172 72566 74228 72604
rect 73836 72258 73892 72268
rect 73948 72322 74004 72334
rect 73948 72270 73950 72322
rect 74002 72270 74004 72322
rect 73388 71988 73444 71998
rect 73388 71894 73444 71932
rect 73948 71988 74004 72270
rect 73948 71922 74004 71932
rect 74060 72324 74116 72334
rect 74060 71986 74116 72268
rect 74060 71934 74062 71986
rect 74114 71934 74116 71986
rect 74060 71922 74116 71934
rect 73500 71650 73556 71662
rect 73500 71598 73502 71650
rect 73554 71598 73556 71650
rect 73276 70756 73332 70766
rect 73500 70756 73556 71598
rect 74172 71650 74228 71662
rect 74172 71598 74174 71650
rect 74226 71598 74228 71650
rect 73724 70756 73780 70766
rect 73500 70754 73780 70756
rect 73500 70702 73726 70754
rect 73778 70702 73780 70754
rect 73500 70700 73780 70702
rect 74172 70756 74228 71598
rect 74396 70756 74452 70766
rect 74172 70700 74396 70756
rect 73276 5234 73332 70700
rect 73500 50708 73556 50718
rect 73500 50614 73556 50652
rect 73388 50370 73444 50382
rect 73388 50318 73390 50370
rect 73442 50318 73444 50370
rect 73388 49810 73444 50318
rect 73388 49758 73390 49810
rect 73442 49758 73444 49810
rect 73388 49746 73444 49758
rect 73612 49812 73668 49822
rect 73612 49718 73668 49756
rect 73276 5182 73278 5234
rect 73330 5182 73332 5234
rect 73276 5170 73332 5182
rect 73388 5794 73444 5806
rect 73388 5742 73390 5794
rect 73442 5742 73444 5794
rect 73388 4452 73444 5742
rect 73388 4386 73444 4396
rect 73500 5682 73556 5694
rect 73500 5630 73502 5682
rect 73554 5630 73556 5682
rect 73500 5012 73556 5630
rect 73724 5236 73780 70700
rect 74396 70662 74452 70700
rect 74172 70532 74228 70542
rect 74060 50708 74116 50718
rect 74172 50708 74228 70476
rect 74844 70532 74900 74172
rect 74956 74162 75012 74172
rect 75628 74004 75684 74734
rect 75516 73948 75684 74004
rect 76300 74004 76356 74014
rect 74956 73332 75012 73342
rect 74956 73238 75012 73276
rect 75516 73220 75572 73948
rect 76300 73910 76356 73948
rect 77308 74004 77364 74014
rect 77308 73910 77364 73948
rect 76748 73330 76804 73342
rect 76748 73278 76750 73330
rect 76802 73278 76804 73330
rect 75516 73154 75572 73164
rect 75964 73218 76020 73230
rect 75964 73166 75966 73218
rect 76018 73166 76020 73218
rect 75068 72546 75124 72558
rect 75068 72494 75070 72546
rect 75122 72494 75124 72546
rect 74956 71762 75012 71774
rect 74956 71710 74958 71762
rect 75010 71710 75012 71762
rect 74956 71316 75012 71710
rect 74956 71250 75012 71260
rect 74844 70466 74900 70476
rect 74956 71090 75012 71102
rect 74956 71038 74958 71090
rect 75010 71038 75012 71090
rect 74956 70084 75012 71038
rect 75068 70644 75124 72494
rect 75964 71876 76020 73166
rect 75964 71810 76020 71820
rect 76076 72434 76132 72446
rect 76076 72382 76078 72434
rect 76130 72382 76132 72434
rect 75628 71652 75684 71662
rect 75516 71650 75684 71652
rect 75516 71598 75630 71650
rect 75682 71598 75684 71650
rect 75516 71596 75684 71598
rect 75068 70578 75124 70588
rect 75404 70756 75460 70766
rect 74956 70018 75012 70028
rect 75068 70082 75124 70094
rect 75068 70030 75070 70082
rect 75122 70030 75124 70082
rect 74956 69522 75012 69534
rect 74956 69470 74958 69522
rect 75010 69470 75012 69522
rect 74956 69412 75012 69470
rect 74956 69346 75012 69356
rect 74284 69298 74340 69310
rect 74284 69246 74286 69298
rect 74338 69246 74340 69298
rect 74284 69188 74340 69246
rect 74284 69122 74340 69132
rect 74508 69188 74564 69198
rect 74508 68850 74564 69132
rect 74508 68798 74510 68850
rect 74562 68798 74564 68850
rect 74508 68786 74564 68798
rect 75068 68292 75124 70030
rect 75068 68226 75124 68236
rect 75180 68514 75236 68526
rect 75180 68462 75182 68514
rect 75234 68462 75236 68514
rect 74956 67956 75012 67966
rect 74956 67862 75012 67900
rect 75180 67172 75236 68462
rect 75180 67106 75236 67116
rect 75180 66946 75236 66958
rect 75180 66894 75182 66946
rect 75234 66894 75236 66946
rect 75068 66386 75124 66398
rect 75068 66334 75070 66386
rect 75122 66334 75124 66386
rect 74956 65378 75012 65390
rect 74956 65326 74958 65378
rect 75010 65326 75012 65378
rect 74956 65044 75012 65326
rect 74956 64978 75012 64988
rect 74956 64818 75012 64830
rect 74956 64766 74958 64818
rect 75010 64766 75012 64818
rect 74284 64594 74340 64606
rect 74284 64542 74286 64594
rect 74338 64542 74340 64594
rect 74284 64484 74340 64542
rect 74284 64418 74340 64428
rect 74508 64484 74564 64494
rect 74508 64146 74564 64428
rect 74956 64372 75012 64766
rect 75068 64708 75124 66334
rect 75180 65156 75236 66894
rect 75180 65090 75236 65100
rect 75068 64642 75124 64652
rect 74956 64306 75012 64316
rect 74508 64094 74510 64146
rect 74562 64094 74564 64146
rect 74508 64082 74564 64094
rect 75180 63810 75236 63822
rect 75180 63758 75182 63810
rect 75234 63758 75236 63810
rect 74956 63252 75012 63262
rect 74620 63250 75012 63252
rect 74620 63198 74958 63250
rect 75010 63198 75012 63250
rect 74620 63196 75012 63198
rect 74620 60676 74676 63196
rect 74956 63186 75012 63196
rect 75068 62242 75124 62254
rect 75068 62190 75070 62242
rect 75122 62190 75124 62242
rect 74956 61684 75012 61694
rect 74620 60610 74676 60620
rect 74732 61682 75012 61684
rect 74732 61630 74958 61682
rect 75010 61630 75012 61682
rect 74732 61628 75012 61630
rect 74284 59890 74340 59902
rect 74284 59838 74286 59890
rect 74338 59838 74340 59890
rect 74284 59780 74340 59838
rect 74284 59714 74340 59724
rect 74508 59780 74564 59790
rect 74508 59442 74564 59724
rect 74508 59390 74510 59442
rect 74562 59390 74564 59442
rect 74508 59378 74564 59390
rect 74732 59220 74788 61628
rect 74956 61618 75012 61628
rect 74956 60674 75012 60686
rect 74956 60622 74958 60674
rect 75010 60622 75012 60674
rect 74956 60340 75012 60622
rect 74732 59154 74788 59164
rect 74844 60284 75012 60340
rect 74844 58212 74900 60284
rect 75068 60228 75124 62190
rect 75180 61348 75236 63758
rect 75180 61282 75236 61292
rect 75068 60162 75124 60172
rect 74956 60116 75012 60126
rect 74956 60022 75012 60060
rect 75180 59106 75236 59118
rect 75180 59054 75182 59106
rect 75234 59054 75236 59106
rect 74844 58146 74900 58156
rect 75068 58546 75124 58558
rect 75068 58494 75070 58546
rect 75122 58494 75124 58546
rect 74956 57540 75012 57550
rect 74844 57538 75012 57540
rect 74844 57486 74958 57538
rect 75010 57486 75012 57538
rect 74844 57484 75012 57486
rect 74844 54628 74900 57484
rect 74956 57474 75012 57484
rect 74956 56980 75012 56990
rect 74956 56886 75012 56924
rect 75068 56308 75124 58494
rect 75180 56756 75236 59054
rect 75180 56690 75236 56700
rect 75068 56242 75124 56252
rect 75068 55970 75124 55982
rect 75068 55918 75070 55970
rect 75122 55918 75124 55970
rect 75068 54740 75124 55918
rect 75068 54674 75124 54684
rect 75180 55410 75236 55422
rect 75180 55358 75182 55410
rect 75234 55358 75236 55410
rect 74844 54562 74900 54572
rect 75068 54402 75124 54414
rect 75068 54350 75070 54402
rect 75122 54350 75124 54402
rect 75068 53956 75124 54350
rect 75068 53890 75124 53900
rect 74956 53844 75012 53854
rect 74956 53750 75012 53788
rect 75068 52834 75124 52846
rect 75068 52782 75070 52834
rect 75122 52782 75124 52834
rect 75068 52164 75124 52782
rect 75180 52836 75236 55358
rect 75180 52770 75236 52780
rect 75068 52098 75124 52108
rect 75180 52274 75236 52286
rect 75180 52222 75182 52274
rect 75234 52222 75236 52274
rect 75068 51266 75124 51278
rect 75068 51214 75070 51266
rect 75122 51214 75124 51266
rect 74956 50708 75012 50718
rect 74116 50652 74228 50708
rect 74844 50706 75012 50708
rect 74844 50654 74958 50706
rect 75010 50654 75012 50706
rect 74844 50652 75012 50654
rect 74060 50576 74116 50652
rect 73836 50036 73892 50046
rect 73836 49942 73892 49980
rect 74060 49810 74116 49822
rect 74060 49758 74062 49810
rect 74114 49758 74116 49810
rect 73948 49698 74004 49710
rect 73948 49646 73950 49698
rect 74002 49646 74004 49698
rect 73948 20188 74004 49646
rect 74060 48692 74116 49758
rect 74844 49252 74900 50652
rect 74956 50642 75012 50652
rect 75068 49700 75124 51214
rect 75180 50596 75236 52222
rect 75180 50530 75236 50540
rect 75068 49634 75124 49644
rect 75180 49698 75236 49710
rect 75180 49646 75182 49698
rect 75234 49646 75236 49698
rect 74844 49186 74900 49196
rect 74956 49140 75012 49150
rect 74956 49046 75012 49084
rect 74060 48626 74116 48636
rect 74956 48244 75012 48254
rect 74508 48242 75012 48244
rect 74508 48190 74958 48242
rect 75010 48190 75012 48242
rect 74508 48188 75012 48190
rect 74508 48130 74564 48188
rect 74956 48178 75012 48188
rect 74508 48078 74510 48130
rect 74562 48078 74564 48130
rect 74396 47236 74452 47246
rect 74284 47234 74452 47236
rect 74284 47182 74398 47234
rect 74450 47182 74452 47234
rect 74284 47180 74452 47182
rect 74284 47012 74340 47180
rect 74396 47170 74452 47180
rect 74284 45780 74340 46956
rect 74508 46900 74564 48078
rect 74956 47458 75012 47470
rect 74956 47406 74958 47458
rect 75010 47406 75012 47458
rect 74956 47012 75012 47406
rect 75180 47348 75236 49646
rect 75180 47282 75236 47292
rect 74956 46946 75012 46956
rect 74508 46834 74564 46844
rect 74956 46676 75012 46686
rect 74284 45714 74340 45724
rect 74508 46674 75012 46676
rect 74508 46622 74958 46674
rect 75010 46622 75012 46674
rect 74508 46620 75012 46622
rect 74508 46562 74564 46620
rect 74956 46610 75012 46620
rect 74508 46510 74510 46562
rect 74562 46510 74564 46562
rect 74396 45668 74452 45678
rect 74396 45574 74452 45612
rect 74508 45332 74564 46510
rect 74956 45890 75012 45902
rect 74956 45838 74958 45890
rect 75010 45838 75012 45890
rect 74956 45668 75012 45838
rect 74956 45602 75012 45612
rect 74508 45266 74564 45276
rect 74956 45108 75012 45118
rect 74508 45106 75012 45108
rect 74508 45054 74958 45106
rect 75010 45054 75012 45106
rect 74508 45052 75012 45054
rect 74508 44994 74564 45052
rect 74956 45042 75012 45052
rect 74508 44942 74510 44994
rect 74562 44942 74564 44994
rect 74396 44098 74452 44110
rect 74396 44046 74398 44098
rect 74450 44046 74452 44098
rect 74396 43764 74452 44046
rect 74508 44100 74564 44942
rect 74508 44034 74564 44044
rect 74956 44322 75012 44334
rect 74956 44270 74958 44322
rect 75010 44270 75012 44322
rect 74396 43698 74452 43708
rect 74956 43764 75012 44270
rect 74956 43698 75012 43708
rect 74956 43540 75012 43550
rect 74508 43538 75012 43540
rect 74508 43486 74958 43538
rect 75010 43486 75012 43538
rect 74508 43484 75012 43486
rect 74508 43426 74564 43484
rect 74956 43474 75012 43484
rect 74508 43374 74510 43426
rect 74562 43374 74564 43426
rect 74396 42756 74452 42766
rect 74396 42530 74452 42700
rect 74396 42478 74398 42530
rect 74450 42478 74452 42530
rect 74396 42084 74452 42478
rect 74508 42532 74564 43374
rect 74956 42756 75012 42766
rect 74956 42662 75012 42700
rect 74508 42466 74564 42476
rect 74396 42018 74452 42028
rect 74956 41972 75012 41982
rect 74508 41970 75012 41972
rect 74508 41918 74958 41970
rect 75010 41918 75012 41970
rect 74508 41916 75012 41918
rect 74508 41858 74564 41916
rect 74956 41906 75012 41916
rect 74508 41806 74510 41858
rect 74562 41806 74564 41858
rect 74396 41188 74452 41198
rect 74396 40962 74452 41132
rect 74396 40910 74398 40962
rect 74450 40910 74452 40962
rect 74396 40516 74452 40910
rect 74508 40964 74564 41806
rect 74956 41188 75012 41198
rect 74956 41094 75012 41132
rect 74508 40898 74564 40908
rect 74396 40450 74452 40460
rect 74508 40404 74564 40414
rect 74956 40404 75012 40414
rect 74508 40402 75012 40404
rect 74508 40350 74510 40402
rect 74562 40350 74958 40402
rect 75010 40350 75012 40402
rect 74508 40348 75012 40350
rect 74508 39620 74564 40348
rect 74956 40338 75012 40348
rect 74508 39554 74564 39564
rect 74956 39618 75012 39630
rect 74956 39566 74958 39618
rect 75010 39566 75012 39618
rect 74508 39396 74564 39406
rect 74508 39302 74564 39340
rect 74956 39396 75012 39566
rect 74956 39330 75012 39340
rect 74508 38948 74564 38958
rect 74508 38854 74564 38892
rect 74956 38948 75012 38958
rect 74956 38834 75012 38892
rect 74956 38782 74958 38834
rect 75010 38782 75012 38834
rect 74956 38770 75012 38782
rect 74956 38050 75012 38062
rect 74956 37998 74958 38050
rect 75010 37998 75012 38050
rect 74508 37828 74564 37838
rect 74508 37734 74564 37772
rect 74956 37828 75012 37998
rect 74956 37762 75012 37772
rect 74508 37380 74564 37390
rect 74508 37286 74564 37324
rect 74956 37380 75012 37390
rect 74956 37266 75012 37324
rect 74956 37214 74958 37266
rect 75010 37214 75012 37266
rect 74956 37202 75012 37214
rect 74956 36482 75012 36494
rect 74956 36430 74958 36482
rect 75010 36430 75012 36482
rect 74508 36260 74564 36270
rect 74508 36166 74564 36204
rect 74956 36260 75012 36430
rect 74956 36194 75012 36204
rect 74508 35812 74564 35822
rect 74508 35718 74564 35756
rect 74956 35812 75012 35822
rect 74956 35698 75012 35756
rect 74956 35646 74958 35698
rect 75010 35646 75012 35698
rect 74956 35634 75012 35646
rect 74956 34914 75012 34926
rect 74956 34862 74958 34914
rect 75010 34862 75012 34914
rect 74508 34804 74564 34814
rect 74508 34710 74564 34748
rect 74956 34804 75012 34862
rect 74956 34738 75012 34748
rect 74508 34244 74564 34254
rect 74508 34150 74564 34188
rect 74956 34244 75012 34254
rect 74956 34130 75012 34188
rect 74956 34078 74958 34130
rect 75010 34078 75012 34130
rect 74956 34066 75012 34078
rect 74956 33346 75012 33358
rect 74956 33294 74958 33346
rect 75010 33294 75012 33346
rect 74508 33124 74564 33134
rect 74508 33030 74564 33068
rect 74956 33124 75012 33294
rect 74956 33058 75012 33068
rect 74508 32676 74564 32686
rect 74508 32582 74564 32620
rect 74956 32676 75012 32686
rect 74956 32562 75012 32620
rect 74956 32510 74958 32562
rect 75010 32510 75012 32562
rect 74956 32498 75012 32510
rect 74956 31778 75012 31790
rect 74956 31726 74958 31778
rect 75010 31726 75012 31778
rect 74508 31556 74564 31566
rect 74508 31462 74564 31500
rect 74956 31556 75012 31726
rect 74956 31490 75012 31500
rect 74508 31108 74564 31118
rect 74508 31014 74564 31052
rect 74956 31108 75012 31118
rect 74956 30994 75012 31052
rect 74956 30942 74958 30994
rect 75010 30942 75012 30994
rect 74956 30930 75012 30942
rect 74956 30210 75012 30222
rect 74956 30158 74958 30210
rect 75010 30158 75012 30210
rect 74508 30100 74564 30110
rect 74508 30006 74564 30044
rect 74956 30100 75012 30158
rect 74956 30034 75012 30044
rect 74508 29540 74564 29550
rect 74508 29446 74564 29484
rect 74956 29540 75012 29550
rect 74956 29426 75012 29484
rect 74956 29374 74958 29426
rect 75010 29374 75012 29426
rect 74956 29362 75012 29374
rect 74508 28642 74564 28654
rect 74508 28590 74510 28642
rect 74562 28590 74564 28642
rect 74508 28420 74564 28590
rect 74508 28354 74564 28364
rect 74956 28642 75012 28654
rect 74956 28590 74958 28642
rect 75010 28590 75012 28642
rect 74956 28420 75012 28590
rect 74956 28354 75012 28364
rect 74508 27972 74564 27982
rect 74508 27878 74564 27916
rect 74956 27972 75012 27982
rect 74956 27858 75012 27916
rect 74956 27806 74958 27858
rect 75010 27806 75012 27858
rect 74956 27794 75012 27806
rect 74956 27074 75012 27086
rect 74956 27022 74958 27074
rect 75010 27022 75012 27074
rect 74508 26962 74564 26974
rect 74508 26910 74510 26962
rect 74562 26910 74564 26962
rect 74508 26852 74564 26910
rect 74508 26786 74564 26796
rect 74956 26852 75012 27022
rect 74956 26786 75012 26796
rect 74508 26404 74564 26414
rect 74508 26310 74564 26348
rect 74956 26404 75012 26414
rect 74956 26290 75012 26348
rect 74956 26238 74958 26290
rect 75010 26238 75012 26290
rect 74956 26226 75012 26238
rect 74956 25506 75012 25518
rect 74956 25454 74958 25506
rect 75010 25454 75012 25506
rect 74508 25284 74564 25294
rect 74508 25190 74564 25228
rect 74956 25284 75012 25454
rect 74956 25218 75012 25228
rect 74508 24724 74564 24734
rect 74508 24630 74564 24668
rect 74956 24724 75012 24734
rect 74956 24630 75012 24668
rect 74956 23938 75012 23950
rect 74956 23886 74958 23938
rect 75010 23886 75012 23938
rect 74508 23716 74564 23726
rect 74508 23622 74564 23660
rect 74956 23716 75012 23886
rect 74956 23650 75012 23660
rect 74508 23268 74564 23278
rect 74508 23174 74564 23212
rect 74956 23268 75012 23278
rect 74956 23154 75012 23212
rect 74956 23102 74958 23154
rect 75010 23102 75012 23154
rect 74956 23090 75012 23102
rect 74956 22370 75012 22382
rect 74956 22318 74958 22370
rect 75010 22318 75012 22370
rect 74508 22148 74564 22158
rect 74508 22054 74564 22092
rect 74956 22148 75012 22318
rect 74956 22082 75012 22092
rect 74508 21700 74564 21710
rect 74508 21606 74564 21644
rect 74956 21700 75012 21710
rect 74956 21586 75012 21644
rect 74956 21534 74958 21586
rect 75010 21534 75012 21586
rect 74956 21522 75012 21534
rect 74956 20802 75012 20814
rect 74956 20750 74958 20802
rect 75010 20750 75012 20802
rect 74508 20580 74564 20590
rect 74508 20486 74564 20524
rect 74956 20580 75012 20750
rect 74956 20514 75012 20524
rect 73948 20132 74228 20188
rect 73836 5794 73892 5806
rect 73836 5742 73838 5794
rect 73890 5742 73892 5794
rect 73836 5682 73892 5742
rect 73836 5630 73838 5682
rect 73890 5630 73892 5682
rect 73836 5618 73892 5630
rect 74060 5236 74116 5246
rect 73724 5234 74116 5236
rect 73724 5182 74062 5234
rect 74114 5182 74116 5234
rect 73724 5180 74116 5182
rect 74060 5170 74116 5180
rect 73388 4228 73444 4238
rect 73164 4226 73444 4228
rect 73164 4174 73390 4226
rect 73442 4174 73444 4226
rect 73164 4172 73444 4174
rect 73388 4162 73444 4172
rect 73500 3668 73556 4956
rect 74172 3780 74228 20132
rect 74956 20020 75012 20030
rect 74508 20018 75012 20020
rect 74508 19966 74958 20018
rect 75010 19966 75012 20018
rect 74508 19964 75012 19966
rect 74508 19908 74564 19964
rect 74956 19954 75012 19964
rect 74396 19906 74564 19908
rect 74396 19854 74510 19906
rect 74562 19854 74564 19906
rect 74396 19852 74564 19854
rect 74396 19012 74452 19852
rect 74508 19842 74564 19852
rect 74956 19234 75012 19246
rect 74956 19182 74958 19234
rect 75010 19182 75012 19234
rect 74508 19124 74564 19134
rect 74508 19030 74564 19068
rect 74956 19124 75012 19182
rect 74956 19058 75012 19068
rect 74396 18946 74452 18956
rect 74508 18452 74564 18462
rect 74508 18358 74564 18396
rect 74956 18452 75012 18462
rect 74956 18358 75012 18396
rect 74956 17666 75012 17678
rect 74956 17614 74958 17666
rect 75010 17614 75012 17666
rect 74508 17556 74564 17566
rect 74508 17462 74564 17500
rect 74956 17556 75012 17614
rect 74956 17490 75012 17500
rect 74508 16996 74564 17006
rect 74508 16902 74564 16940
rect 74956 16996 75012 17006
rect 74956 16882 75012 16940
rect 74956 16830 74958 16882
rect 75010 16830 75012 16882
rect 74956 16818 75012 16830
rect 74508 16100 74564 16110
rect 74508 16006 74564 16044
rect 74956 16100 75012 16110
rect 74956 16006 75012 16044
rect 74508 15428 74564 15438
rect 74508 15334 74564 15372
rect 74956 15428 75012 15438
rect 74956 15314 75012 15372
rect 74956 15262 74958 15314
rect 75010 15262 75012 15314
rect 74956 15250 75012 15262
rect 74956 14530 75012 14542
rect 74956 14478 74958 14530
rect 75010 14478 75012 14530
rect 74508 14308 74564 14318
rect 74508 14214 74564 14252
rect 74956 14308 75012 14478
rect 74956 14242 75012 14252
rect 74508 13860 74564 13870
rect 74508 13766 74564 13804
rect 74956 13860 75012 13870
rect 74396 13748 74452 13758
rect 74396 13076 74452 13692
rect 74956 13746 75012 13804
rect 74956 13694 74958 13746
rect 75010 13694 75012 13746
rect 74956 13682 75012 13694
rect 74508 13076 74564 13086
rect 74396 13074 74564 13076
rect 74396 13022 74510 13074
rect 74562 13022 74564 13074
rect 74396 13020 74564 13022
rect 74508 12964 74564 13020
rect 74956 12964 75012 12974
rect 74508 12962 75012 12964
rect 74508 12910 74958 12962
rect 75010 12910 75012 12962
rect 74508 12908 75012 12910
rect 74956 12898 75012 12908
rect 74508 12292 74564 12302
rect 74508 12198 74564 12236
rect 74956 12292 75012 12302
rect 74956 12178 75012 12236
rect 74956 12126 74958 12178
rect 75010 12126 75012 12178
rect 74956 12114 75012 12126
rect 74956 11394 75012 11406
rect 74956 11342 74958 11394
rect 75010 11342 75012 11394
rect 74508 11284 74564 11294
rect 74508 11190 74564 11228
rect 74956 11284 75012 11342
rect 74956 11218 75012 11228
rect 74508 10724 74564 10734
rect 74508 10630 74564 10668
rect 74956 10724 75012 10734
rect 74956 10610 75012 10668
rect 74956 10558 74958 10610
rect 75010 10558 75012 10610
rect 74956 10546 75012 10558
rect 74956 9826 75012 9838
rect 74956 9774 74958 9826
rect 75010 9774 75012 9826
rect 74508 9604 74564 9614
rect 74508 9510 74564 9548
rect 74956 9604 75012 9774
rect 74956 9538 75012 9548
rect 74508 9156 74564 9166
rect 74508 9062 74564 9100
rect 74956 9156 75012 9166
rect 74956 9042 75012 9100
rect 74956 8990 74958 9042
rect 75010 8990 75012 9042
rect 74956 8978 75012 8990
rect 74956 8258 75012 8270
rect 74956 8206 74958 8258
rect 75010 8206 75012 8258
rect 74508 8036 74564 8046
rect 74508 7942 74564 7980
rect 74956 8036 75012 8206
rect 74956 7970 75012 7980
rect 74508 7588 74564 7598
rect 74508 7494 74564 7532
rect 74956 7588 75012 7598
rect 74956 7474 75012 7532
rect 74956 7422 74958 7474
rect 75010 7422 75012 7474
rect 74956 7410 75012 7422
rect 74956 6690 75012 6702
rect 74956 6638 74958 6690
rect 75010 6638 75012 6690
rect 74508 6466 74564 6478
rect 74508 6414 74510 6466
rect 74562 6414 74564 6466
rect 74508 6132 74564 6414
rect 74508 6066 74564 6076
rect 74956 6132 75012 6638
rect 74956 6066 75012 6076
rect 74956 5908 75012 5918
rect 74508 5906 75012 5908
rect 74508 5854 74958 5906
rect 75010 5854 75012 5906
rect 74508 5852 75012 5854
rect 74508 5794 74564 5852
rect 74956 5842 75012 5852
rect 74508 5742 74510 5794
rect 74562 5742 74564 5794
rect 74508 4564 74564 5742
rect 75068 5012 75124 5022
rect 75068 4918 75124 4956
rect 74508 4498 74564 4508
rect 74396 4452 74452 4462
rect 74396 4358 74452 4396
rect 75404 4226 75460 70700
rect 75516 69860 75572 71596
rect 75628 71586 75684 71596
rect 76076 70644 76132 72382
rect 76748 72436 76804 73278
rect 77868 73218 77924 73230
rect 77868 73166 77870 73218
rect 77922 73166 77924 73218
rect 77868 72548 77924 73166
rect 77868 72482 77924 72492
rect 76748 72370 76804 72380
rect 76748 71764 76804 71774
rect 76748 71670 76804 71708
rect 77868 71650 77924 71662
rect 77868 71598 77870 71650
rect 77922 71598 77924 71650
rect 77868 71204 77924 71598
rect 77868 71138 77924 71148
rect 76300 70868 76356 70878
rect 76300 70774 76356 70812
rect 77308 70868 77364 70878
rect 77308 70754 77364 70812
rect 77308 70702 77310 70754
rect 77362 70702 77364 70754
rect 77308 70644 77364 70702
rect 77308 70588 77588 70644
rect 76076 70578 76132 70588
rect 76300 70306 76356 70318
rect 76300 70254 76302 70306
rect 76354 70254 76356 70306
rect 76300 70084 76356 70254
rect 76860 70084 76916 70094
rect 76300 70082 76916 70084
rect 76300 70030 76862 70082
rect 76914 70030 76916 70082
rect 76300 70028 76916 70030
rect 75516 69794 75572 69804
rect 76300 69300 76356 69310
rect 76300 69206 76356 69244
rect 76300 68740 76356 68750
rect 76300 68646 76356 68684
rect 76748 67844 76804 70028
rect 76860 70018 76916 70028
rect 77308 69300 77364 69310
rect 77308 69188 77364 69244
rect 77308 69186 77476 69188
rect 77308 69134 77310 69186
rect 77362 69134 77476 69186
rect 77308 69132 77476 69134
rect 77308 69122 77364 69132
rect 76860 68740 76916 68750
rect 76860 68516 76916 68684
rect 76860 68514 77028 68516
rect 76860 68462 76862 68514
rect 76914 68462 77028 68514
rect 76860 68460 77028 68462
rect 76860 68450 76916 68460
rect 76748 67778 76804 67788
rect 76300 67732 76356 67742
rect 76300 67638 76356 67676
rect 76300 67172 76356 67182
rect 76300 67078 76356 67116
rect 76860 67172 76916 67182
rect 76860 66946 76916 67116
rect 76860 66894 76862 66946
rect 76914 66894 76916 66946
rect 76300 66162 76356 66174
rect 76300 66110 76302 66162
rect 76354 66110 76356 66162
rect 76300 66052 76356 66110
rect 76300 65986 76356 65996
rect 76300 65604 76356 65614
rect 76860 65604 76916 66894
rect 76972 66500 77028 68460
rect 77308 67732 77364 67742
rect 77308 66948 77364 67676
rect 77420 67172 77476 69132
rect 77532 68516 77588 70588
rect 77532 68450 77588 68460
rect 77420 67106 77476 67116
rect 77308 66892 77476 66948
rect 76972 66434 77028 66444
rect 76300 65602 76804 65604
rect 76300 65550 76302 65602
rect 76354 65550 76804 65602
rect 76300 65548 76804 65550
rect 76300 65538 76356 65548
rect 76748 65380 76804 65548
rect 77308 66052 77364 66062
rect 77308 65604 77364 65996
rect 77420 65828 77476 66892
rect 77420 65762 77476 65772
rect 77308 65548 77588 65604
rect 76860 65538 76916 65548
rect 76860 65380 76916 65390
rect 76748 65378 76916 65380
rect 76748 65326 76862 65378
rect 76914 65326 76916 65378
rect 76748 65324 76916 65326
rect 76300 64596 76356 64606
rect 76300 64502 76356 64540
rect 76300 64034 76356 64046
rect 76300 63982 76302 64034
rect 76354 63982 76356 64034
rect 76300 63812 76356 63982
rect 76300 63746 76356 63756
rect 76748 63140 76804 65324
rect 76860 65314 76916 65324
rect 77308 64596 77364 64606
rect 77308 64484 77364 64540
rect 77308 64482 77476 64484
rect 77308 64430 77310 64482
rect 77362 64430 77476 64482
rect 77308 64428 77476 64430
rect 77308 64418 77364 64428
rect 76860 63922 76916 63934
rect 76860 63870 76862 63922
rect 76914 63870 76916 63922
rect 76860 63812 76916 63870
rect 76860 63252 76916 63756
rect 76860 63196 77140 63252
rect 76748 63074 76804 63084
rect 76300 63028 76356 63038
rect 76300 62934 76356 62972
rect 76300 62468 76356 62478
rect 76300 62466 76916 62468
rect 76300 62414 76302 62466
rect 76354 62414 76916 62466
rect 76300 62412 76916 62414
rect 76300 62402 76356 62412
rect 76860 62244 76916 62412
rect 76860 62242 77028 62244
rect 76860 62190 76862 62242
rect 76914 62190 77028 62242
rect 76860 62188 77028 62190
rect 76860 62178 76916 62188
rect 76300 61460 76356 61470
rect 76300 61366 76356 61404
rect 76300 60900 76356 60910
rect 76300 60898 76916 60900
rect 76300 60846 76302 60898
rect 76354 60846 76916 60898
rect 76300 60844 76916 60846
rect 76300 60834 76356 60844
rect 76860 60674 76916 60844
rect 76860 60622 76862 60674
rect 76914 60622 76916 60674
rect 76860 60004 76916 60622
rect 76972 60564 77028 62188
rect 77084 61796 77140 63196
rect 77308 63028 77364 63038
rect 77308 62914 77364 62972
rect 77308 62862 77310 62914
rect 77362 62862 77364 62914
rect 77308 62244 77364 62862
rect 77420 62468 77476 64428
rect 77532 63924 77588 65548
rect 77532 63858 77588 63868
rect 77420 62402 77476 62412
rect 77308 62188 77476 62244
rect 77084 61730 77140 61740
rect 76972 60498 77028 60508
rect 77196 61460 77252 61470
rect 77196 61348 77252 61404
rect 77308 61348 77364 61358
rect 77196 61346 77364 61348
rect 77196 61294 77310 61346
rect 77362 61294 77364 61346
rect 77196 61292 77364 61294
rect 76860 59948 77028 60004
rect 76300 59892 76356 59902
rect 76300 59798 76356 59836
rect 76300 59332 76356 59342
rect 76300 59330 76804 59332
rect 76300 59278 76302 59330
rect 76354 59278 76804 59330
rect 76300 59276 76804 59278
rect 76300 59266 76356 59276
rect 76748 59108 76804 59276
rect 76860 59108 76916 59118
rect 76748 59106 76916 59108
rect 76748 59054 76862 59106
rect 76914 59054 76916 59106
rect 76748 59052 76916 59054
rect 76300 58324 76356 58334
rect 76300 58230 76356 58268
rect 76300 57764 76356 57774
rect 76300 57670 76356 57708
rect 76748 57316 76804 59052
rect 76860 59042 76916 59052
rect 76972 58436 77028 59948
rect 77196 59108 77252 61292
rect 77308 61282 77364 61292
rect 77420 61124 77476 62188
rect 77420 61058 77476 61068
rect 77308 59892 77364 59902
rect 77308 59780 77364 59836
rect 77308 59778 77476 59780
rect 77308 59726 77310 59778
rect 77362 59726 77476 59778
rect 77308 59724 77476 59726
rect 77308 59714 77364 59724
rect 77196 59042 77252 59052
rect 76972 58370 77028 58380
rect 77308 58324 77364 58334
rect 77308 58210 77364 58268
rect 77308 58158 77310 58210
rect 77362 58158 77364 58210
rect 76860 57764 76916 57774
rect 76860 57540 76916 57708
rect 77308 57540 77364 58158
rect 77420 57764 77476 59724
rect 77420 57698 77476 57708
rect 76860 57538 77028 57540
rect 76860 57486 76862 57538
rect 76914 57486 77028 57538
rect 76860 57484 77028 57486
rect 77308 57484 77476 57540
rect 76860 57474 76916 57484
rect 76748 57250 76804 57260
rect 76300 56756 76356 56766
rect 76300 56662 76356 56700
rect 76300 56196 76356 56206
rect 76300 56102 76356 56140
rect 76860 56196 76916 56206
rect 76860 55468 76916 56140
rect 76972 55748 77028 57484
rect 76972 55682 77028 55692
rect 77308 56756 77364 56766
rect 77308 56642 77364 56700
rect 77308 56590 77310 56642
rect 77362 56590 77364 56642
rect 77308 55524 77364 56590
rect 77420 56420 77476 57484
rect 77420 56354 77476 56364
rect 76860 55412 77028 55468
rect 77308 55458 77364 55468
rect 76300 55188 76356 55198
rect 76300 55094 76356 55132
rect 76300 54628 76356 54638
rect 76300 54534 76356 54572
rect 76860 54628 76916 54638
rect 76860 54402 76916 54572
rect 76860 54350 76862 54402
rect 76914 54350 76916 54402
rect 76300 53620 76356 53630
rect 76300 53526 76356 53564
rect 76860 53284 76916 54350
rect 76972 54404 77028 55412
rect 76972 54338 77028 54348
rect 77308 55188 77364 55198
rect 77308 55074 77364 55132
rect 77308 55022 77310 55074
rect 77362 55022 77364 55074
rect 77308 53844 77364 55022
rect 77308 53778 77364 53788
rect 76860 53218 76916 53228
rect 77308 53620 77364 53630
rect 77308 53506 77364 53564
rect 77308 53454 77310 53506
rect 77362 53454 77364 53506
rect 76300 53060 76356 53070
rect 76300 52966 76356 53004
rect 76860 53060 76916 53070
rect 76860 52834 76916 53004
rect 76860 52782 76862 52834
rect 76914 52782 76916 52834
rect 76300 52052 76356 52062
rect 76300 51958 76356 51996
rect 76860 51716 76916 52782
rect 77308 52388 77364 53454
rect 77308 52322 77364 52332
rect 76860 51650 76916 51660
rect 77308 52162 77364 52174
rect 77308 52110 77310 52162
rect 77362 52110 77364 52162
rect 77308 52052 77364 52110
rect 76300 51492 76356 51502
rect 76300 51398 76356 51436
rect 76860 51492 76916 51502
rect 76860 51266 76916 51436
rect 76860 51214 76862 51266
rect 76914 51214 76916 51266
rect 76300 50484 76356 50494
rect 76300 50390 76356 50428
rect 76860 50372 76916 51214
rect 77308 51044 77364 51996
rect 77308 50978 77364 50988
rect 76860 50306 76916 50316
rect 77308 50484 77364 50494
rect 76300 49924 76356 49934
rect 76300 49830 76356 49868
rect 76860 49924 76916 49934
rect 76860 49698 76916 49868
rect 76860 49646 76862 49698
rect 76914 49646 76916 49698
rect 76860 49028 76916 49646
rect 77308 49700 77364 50428
rect 77308 49634 77364 49644
rect 76860 48962 76916 48972
rect 76300 48916 76356 48926
rect 76300 48822 76356 48860
rect 77308 48916 77364 48926
rect 77308 48802 77364 48860
rect 77308 48750 77310 48802
rect 77362 48750 77364 48802
rect 77308 48356 77364 48750
rect 77308 48290 77364 48300
rect 76748 48242 76804 48254
rect 76748 48190 76750 48242
rect 76802 48190 76804 48242
rect 75964 48130 76020 48142
rect 75964 48078 75966 48130
rect 76018 48078 76020 48130
rect 75964 47124 76020 48078
rect 75964 47058 76020 47068
rect 76076 47346 76132 47358
rect 76076 47294 76078 47346
rect 76130 47294 76132 47346
rect 75964 46562 76020 46574
rect 75964 46510 75966 46562
rect 76018 46510 76020 46562
rect 75964 45668 76020 46510
rect 76076 46340 76132 47294
rect 76748 47236 76804 48190
rect 77868 48130 77924 48142
rect 77868 48078 77870 48130
rect 77922 48078 77924 48130
rect 77868 47684 77924 48078
rect 77868 47618 77924 47628
rect 76748 47170 76804 47180
rect 77196 47236 77252 47246
rect 77196 47142 77252 47180
rect 76076 46274 76132 46284
rect 75964 45602 76020 45612
rect 76076 45778 76132 45790
rect 76076 45726 76078 45778
rect 76130 45726 76132 45778
rect 75964 44994 76020 45006
rect 75964 44942 75966 44994
rect 76018 44942 76020 44994
rect 75964 44324 76020 44942
rect 76076 44996 76132 45726
rect 76076 44930 76132 44940
rect 75964 44258 76020 44268
rect 76076 44210 76132 44222
rect 76076 44158 76078 44210
rect 76130 44158 76132 44210
rect 76076 43764 76132 44158
rect 76076 43698 76132 43708
rect 76076 43426 76132 43438
rect 76076 43374 76078 43426
rect 76130 43374 76132 43426
rect 76076 42980 76132 43374
rect 76076 42914 76132 42924
rect 76076 42642 76132 42654
rect 76076 42590 76078 42642
rect 76130 42590 76132 42642
rect 76076 42308 76132 42590
rect 76076 42242 76132 42252
rect 76076 41858 76132 41870
rect 76076 41806 76078 41858
rect 76130 41806 76132 41858
rect 76076 41636 76132 41806
rect 76076 41570 76132 41580
rect 76076 41074 76132 41086
rect 76076 41022 76078 41074
rect 76130 41022 76132 41074
rect 76076 40964 76132 41022
rect 76076 40898 76132 40908
rect 76076 40404 76132 40414
rect 76076 40310 76132 40348
rect 76076 39620 76132 39630
rect 76076 39526 76132 39564
rect 76076 38948 76132 38958
rect 76076 38854 76132 38892
rect 76076 38276 76132 38286
rect 76076 38162 76132 38220
rect 76076 38110 76078 38162
rect 76130 38110 76132 38162
rect 76076 38098 76132 38110
rect 76076 37604 76132 37614
rect 76076 37378 76132 37548
rect 76076 37326 76078 37378
rect 76130 37326 76132 37378
rect 76076 37314 76132 37326
rect 76076 36932 76132 36942
rect 76076 36594 76132 36876
rect 76076 36542 76078 36594
rect 76130 36542 76132 36594
rect 76076 36530 76132 36542
rect 76076 36260 76132 36270
rect 76076 35810 76132 36204
rect 76076 35758 76078 35810
rect 76130 35758 76132 35810
rect 76076 35746 76132 35758
rect 76748 35698 76804 35710
rect 76748 35646 76750 35698
rect 76802 35646 76804 35698
rect 76076 35588 76132 35598
rect 76076 35026 76132 35532
rect 76076 34974 76078 35026
rect 76130 34974 76132 35026
rect 76076 34962 76132 34974
rect 76748 34692 76804 35646
rect 77868 35586 77924 35598
rect 77868 35534 77870 35586
rect 77922 35534 77924 35586
rect 77868 34916 77924 35534
rect 77868 34850 77924 34860
rect 76748 34626 76804 34636
rect 77196 34692 77252 34702
rect 77196 34598 77252 34636
rect 76076 34244 76132 34254
rect 76076 34150 76132 34188
rect 76076 33572 76132 33582
rect 76076 33458 76132 33516
rect 76076 33406 76078 33458
rect 76130 33406 76132 33458
rect 76076 33394 76132 33406
rect 76076 32900 76132 32910
rect 76076 32674 76132 32844
rect 76076 32622 76078 32674
rect 76130 32622 76132 32674
rect 76076 32610 76132 32622
rect 76076 31892 76132 31902
rect 76076 31798 76132 31836
rect 76076 31556 76132 31566
rect 76076 31106 76132 31500
rect 76076 31054 76078 31106
rect 76130 31054 76132 31106
rect 76076 31042 76132 31054
rect 76748 30994 76804 31006
rect 76748 30942 76750 30994
rect 76802 30942 76804 30994
rect 76076 30884 76132 30894
rect 76076 30210 76132 30828
rect 76076 30158 76078 30210
rect 76130 30158 76132 30210
rect 76076 30146 76132 30158
rect 76748 29988 76804 30942
rect 77868 30882 77924 30894
rect 77868 30830 77870 30882
rect 77922 30830 77924 30882
rect 77868 30324 77924 30830
rect 77868 30258 77924 30268
rect 76748 29922 76804 29932
rect 77196 29988 77252 29998
rect 77196 29894 77252 29932
rect 76076 29540 76132 29550
rect 76076 29446 76132 29484
rect 76076 28868 76132 28878
rect 76076 28754 76132 28812
rect 76076 28702 76078 28754
rect 76130 28702 76132 28754
rect 76076 28690 76132 28702
rect 76076 28196 76132 28206
rect 76076 27970 76132 28140
rect 76076 27918 76078 27970
rect 76130 27918 76132 27970
rect 76076 27906 76132 27918
rect 76076 27524 76132 27534
rect 76076 27186 76132 27468
rect 76076 27134 76078 27186
rect 76130 27134 76132 27186
rect 76076 27122 76132 27134
rect 76076 26852 76132 26862
rect 76076 26402 76132 26796
rect 76076 26350 76078 26402
rect 76130 26350 76132 26402
rect 76076 26338 76132 26350
rect 76972 26292 77028 26302
rect 76972 26290 77252 26292
rect 76972 26238 76974 26290
rect 77026 26238 77252 26290
rect 76972 26236 77252 26238
rect 76972 26226 77028 26236
rect 76076 26180 76132 26190
rect 76076 25618 76132 26124
rect 76076 25566 76078 25618
rect 76130 25566 76132 25618
rect 76076 25554 76132 25566
rect 77196 25282 77252 26236
rect 77868 26178 77924 26190
rect 77868 26126 77870 26178
rect 77922 26126 77924 26178
rect 77868 25508 77924 26126
rect 77868 25442 77924 25452
rect 77196 25230 77198 25282
rect 77250 25230 77252 25282
rect 77196 24948 77252 25230
rect 77196 24882 77252 24892
rect 76076 24836 76132 24846
rect 76076 24742 76132 24780
rect 76076 24164 76132 24174
rect 76076 24050 76132 24108
rect 76076 23998 76078 24050
rect 76130 23998 76132 24050
rect 76076 23986 76132 23998
rect 76076 23492 76132 23502
rect 76076 23266 76132 23436
rect 76076 23214 76078 23266
rect 76130 23214 76132 23266
rect 76076 23202 76132 23214
rect 76076 22820 76132 22830
rect 76076 22482 76132 22764
rect 76076 22430 76078 22482
rect 76130 22430 76132 22482
rect 76076 22418 76132 22430
rect 76076 22148 76132 22158
rect 76076 21698 76132 22092
rect 76076 21646 76078 21698
rect 76130 21646 76132 21698
rect 76076 21634 76132 21646
rect 76972 21588 77028 21598
rect 76972 21586 77252 21588
rect 76972 21534 76974 21586
rect 77026 21534 77252 21586
rect 76972 21532 77252 21534
rect 76972 21522 77028 21532
rect 76076 21476 76132 21486
rect 76076 20914 76132 21420
rect 76076 20862 76078 20914
rect 76130 20862 76132 20914
rect 76076 20850 76132 20862
rect 77196 20578 77252 21532
rect 77868 21474 77924 21486
rect 77868 21422 77870 21474
rect 77922 21422 77924 21474
rect 77868 20804 77924 21422
rect 77868 20738 77924 20748
rect 77196 20526 77198 20578
rect 77250 20526 77252 20578
rect 77196 20244 77252 20526
rect 77196 20178 77252 20188
rect 76076 20132 76132 20142
rect 76076 20038 76132 20076
rect 76076 19460 76132 19470
rect 76076 19346 76132 19404
rect 76076 19294 76078 19346
rect 76130 19294 76132 19346
rect 76076 19282 76132 19294
rect 76076 18788 76132 18798
rect 76076 18450 76132 18732
rect 76076 18398 76078 18450
rect 76130 18398 76132 18450
rect 76076 18386 76132 18398
rect 76076 18116 76132 18126
rect 76076 17778 76132 18060
rect 76076 17726 76078 17778
rect 76130 17726 76132 17778
rect 76076 17714 76132 17726
rect 76076 17444 76132 17454
rect 76076 16994 76132 17388
rect 76076 16942 76078 16994
rect 76130 16942 76132 16994
rect 76076 16930 76132 16942
rect 76748 16882 76804 16894
rect 76748 16830 76750 16882
rect 76802 16830 76804 16882
rect 76076 16772 76132 16782
rect 76076 16210 76132 16716
rect 76076 16158 76078 16210
rect 76130 16158 76132 16210
rect 76076 16146 76132 16158
rect 76748 15876 76804 16830
rect 77868 16882 77924 16894
rect 77868 16830 77870 16882
rect 77922 16830 77924 16882
rect 77868 16100 77924 16830
rect 77868 16034 77924 16044
rect 76748 15810 76804 15820
rect 77196 15876 77252 15886
rect 77196 15782 77252 15820
rect 76076 15428 76132 15438
rect 76076 15334 76132 15372
rect 76076 14756 76132 14766
rect 76076 14642 76132 14700
rect 76076 14590 76078 14642
rect 76130 14590 76132 14642
rect 76076 14578 76132 14590
rect 76076 14084 76132 14094
rect 76076 13858 76132 14028
rect 76076 13806 76078 13858
rect 76130 13806 76132 13858
rect 76076 13794 76132 13806
rect 76076 13412 76132 13422
rect 76076 13074 76132 13356
rect 76076 13022 76078 13074
rect 76130 13022 76132 13074
rect 76076 13010 76132 13022
rect 76076 12740 76132 12750
rect 76076 12290 76132 12684
rect 76076 12238 76078 12290
rect 76130 12238 76132 12290
rect 76076 12226 76132 12238
rect 76748 12178 76804 12190
rect 76748 12126 76750 12178
rect 76802 12126 76804 12178
rect 76076 12068 76132 12078
rect 76076 11506 76132 12012
rect 76076 11454 76078 11506
rect 76130 11454 76132 11506
rect 76076 11442 76132 11454
rect 76748 11172 76804 12126
rect 77868 12066 77924 12078
rect 77868 12014 77870 12066
rect 77922 12014 77924 12066
rect 77868 11396 77924 12014
rect 77868 11330 77924 11340
rect 76748 11106 76804 11116
rect 77196 11172 77252 11182
rect 77196 11078 77252 11116
rect 76076 10724 76132 10734
rect 76076 10630 76132 10668
rect 76076 10052 76132 10062
rect 76076 9938 76132 9996
rect 76076 9886 76078 9938
rect 76130 9886 76132 9938
rect 76076 9874 76132 9886
rect 76076 9380 76132 9390
rect 76076 9154 76132 9324
rect 76076 9102 76078 9154
rect 76130 9102 76132 9154
rect 76076 9090 76132 9102
rect 76076 8372 76132 8382
rect 76076 8278 76132 8316
rect 76076 8036 76132 8046
rect 76076 7586 76132 7980
rect 76076 7534 76078 7586
rect 76130 7534 76132 7586
rect 76076 7522 76132 7534
rect 76748 7474 76804 7486
rect 76748 7422 76750 7474
rect 76802 7422 76804 7474
rect 76076 7364 76132 7374
rect 76076 6690 76132 7308
rect 76076 6638 76078 6690
rect 76130 6638 76132 6690
rect 76076 6626 76132 6638
rect 76748 6580 76804 7422
rect 77868 7362 77924 7374
rect 77868 7310 77870 7362
rect 77922 7310 77924 7362
rect 77868 6804 77924 7310
rect 77868 6738 77924 6748
rect 76748 6514 76804 6524
rect 77196 6580 77252 6590
rect 77196 6486 77252 6524
rect 76076 6020 76132 6030
rect 76076 5926 76132 5964
rect 76748 5908 76804 5918
rect 76524 5906 76804 5908
rect 76524 5854 76750 5906
rect 76802 5854 76804 5906
rect 76524 5852 76804 5854
rect 76524 5122 76580 5852
rect 76748 5842 76804 5852
rect 77868 5794 77924 5806
rect 77868 5742 77870 5794
rect 77922 5742 77924 5794
rect 77868 5348 77924 5742
rect 77868 5282 77924 5292
rect 76524 5070 76526 5122
rect 76578 5070 76580 5122
rect 76524 4900 76580 5070
rect 76524 4834 76580 4844
rect 75404 4174 75406 4226
rect 75458 4174 75460 4226
rect 75404 4162 75460 4174
rect 76412 4450 76468 4462
rect 76412 4398 76414 4450
rect 76466 4398 76468 4450
rect 74172 3714 74228 3724
rect 75628 3780 75684 3790
rect 72716 3378 72772 3388
rect 73164 3612 73556 3668
rect 73836 3668 73892 3678
rect 73164 800 73220 3612
rect 73388 3444 73444 3454
rect 73388 3350 73444 3388
rect 73836 800 73892 3612
rect 75628 3666 75684 3724
rect 75628 3614 75630 3666
rect 75682 3614 75684 3666
rect 75628 3602 75684 3614
rect 76300 3780 76356 3790
rect 76300 3554 76356 3724
rect 76300 3502 76302 3554
rect 76354 3502 76356 3554
rect 76300 3490 76356 3502
rect 74508 3444 74564 3454
rect 74508 800 74564 3388
rect 75068 3444 75124 3454
rect 75068 3350 75124 3388
rect 76412 3444 76468 4398
rect 76972 3668 77028 3678
rect 76972 3574 77028 3612
rect 76412 3378 76468 3388
rect 5264 0 5376 800
rect 5936 0 6048 800
rect 6608 0 6720 800
rect 7280 0 7392 800
rect 7952 0 8064 800
rect 8624 0 8736 800
rect 9296 0 9408 800
rect 9968 0 10080 800
rect 10640 0 10752 800
rect 11312 0 11424 800
rect 11984 0 12096 800
rect 12656 0 12768 800
rect 13328 0 13440 800
rect 14000 0 14112 800
rect 14672 0 14784 800
rect 15344 0 15456 800
rect 16016 0 16128 800
rect 16688 0 16800 800
rect 17360 0 17472 800
rect 18032 0 18144 800
rect 18704 0 18816 800
rect 19376 0 19488 800
rect 20048 0 20160 800
rect 20720 0 20832 800
rect 21392 0 21504 800
rect 22064 0 22176 800
rect 22736 0 22848 800
rect 23408 0 23520 800
rect 24080 0 24192 800
rect 24752 0 24864 800
rect 25424 0 25536 800
rect 26096 0 26208 800
rect 26768 0 26880 800
rect 27440 0 27552 800
rect 28112 0 28224 800
rect 28784 0 28896 800
rect 29456 0 29568 800
rect 30128 0 30240 800
rect 30800 0 30912 800
rect 31472 0 31584 800
rect 32144 0 32256 800
rect 32816 0 32928 800
rect 33488 0 33600 800
rect 34160 0 34272 800
rect 34832 0 34944 800
rect 35504 0 35616 800
rect 36176 0 36288 800
rect 36848 0 36960 800
rect 37520 0 37632 800
rect 38192 0 38304 800
rect 38864 0 38976 800
rect 39536 0 39648 800
rect 40208 0 40320 800
rect 40880 0 40992 800
rect 41552 0 41664 800
rect 42224 0 42336 800
rect 42896 0 43008 800
rect 43568 0 43680 800
rect 44240 0 44352 800
rect 44912 0 45024 800
rect 45584 0 45696 800
rect 46256 0 46368 800
rect 46928 0 47040 800
rect 47600 0 47712 800
rect 48272 0 48384 800
rect 48944 0 49056 800
rect 49616 0 49728 800
rect 50288 0 50400 800
rect 50960 0 51072 800
rect 51632 0 51744 800
rect 52304 0 52416 800
rect 52976 0 53088 800
rect 53648 0 53760 800
rect 54320 0 54432 800
rect 54992 0 55104 800
rect 55664 0 55776 800
rect 56336 0 56448 800
rect 57008 0 57120 800
rect 57680 0 57792 800
rect 58352 0 58464 800
rect 59024 0 59136 800
rect 59696 0 59808 800
rect 60368 0 60480 800
rect 61040 0 61152 800
rect 61712 0 61824 800
rect 62384 0 62496 800
rect 63056 0 63168 800
rect 63728 0 63840 800
rect 64400 0 64512 800
rect 65072 0 65184 800
rect 65744 0 65856 800
rect 66416 0 66528 800
rect 67088 0 67200 800
rect 67760 0 67872 800
rect 68432 0 68544 800
rect 69104 0 69216 800
rect 69776 0 69888 800
rect 70448 0 70560 800
rect 71120 0 71232 800
rect 71792 0 71904 800
rect 72464 0 72576 800
rect 73136 0 73248 800
rect 73808 0 73920 800
rect 74480 0 74592 800
<< via2 >>
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 3052 74898 3108 74900
rect 3052 74846 3054 74898
rect 3054 74846 3106 74898
rect 3106 74846 3108 74898
rect 3052 74844 3108 74846
rect 2044 74508 2100 74564
rect 2268 74002 2324 74004
rect 2268 73950 2270 74002
rect 2270 73950 2322 74002
rect 2322 73950 2324 74002
rect 2268 73948 2324 73950
rect 3052 73330 3108 73332
rect 3052 73278 3054 73330
rect 3054 73278 3106 73330
rect 3106 73278 3108 73330
rect 3052 73276 3108 73278
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 73724 75068 73780 75124
rect 3500 73500 3556 73556
rect 3612 74844 3668 74900
rect 1932 73164 1988 73220
rect 3052 72268 3108 72324
rect 2044 71820 2100 71876
rect 3052 71762 3108 71764
rect 3052 71710 3054 71762
rect 3054 71710 3106 71762
rect 3106 71710 3108 71762
rect 3052 71708 3108 71710
rect 1820 70476 1876 70532
rect 1932 70306 1988 70308
rect 1932 70254 1934 70306
rect 1934 70254 1986 70306
rect 1986 70254 1988 70306
rect 1932 70252 1988 70254
rect 1708 69244 1764 69300
rect 2044 69804 2100 69860
rect 2156 70700 2212 70756
rect 2268 69298 2324 69300
rect 2268 69246 2270 69298
rect 2270 69246 2322 69298
rect 2322 69246 2324 69298
rect 2268 69244 2324 69246
rect 2156 69132 2212 69188
rect 3388 70924 3444 70980
rect 3388 69916 3444 69972
rect 3052 69132 3108 69188
rect 1820 67788 1876 67844
rect 2268 68738 2324 68740
rect 2268 68686 2270 68738
rect 2270 68686 2322 68738
rect 2322 68686 2324 68738
rect 2268 68684 2324 68686
rect 2156 67340 2212 67396
rect 2268 67730 2324 67732
rect 2268 67678 2270 67730
rect 2270 67678 2322 67730
rect 2322 67678 2324 67730
rect 2268 67676 2324 67678
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 4172 74002 4228 74004
rect 4172 73950 4174 74002
rect 4174 73950 4226 74002
rect 4226 73950 4228 74002
rect 4172 73948 4228 73950
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 68908 73554 68964 73556
rect 68908 73502 68910 73554
rect 68910 73502 68962 73554
rect 68962 73502 68964 73554
rect 68908 73500 68964 73502
rect 69020 73442 69076 73444
rect 69020 73390 69022 73442
rect 69022 73390 69074 73442
rect 69074 73390 69076 73442
rect 69020 73388 69076 73390
rect 3836 73276 3892 73332
rect 3612 72604 3668 72660
rect 3724 72492 3780 72548
rect 72492 73276 72548 73332
rect 4844 73164 4900 73220
rect 5404 73218 5460 73220
rect 5404 73166 5406 73218
rect 5406 73166 5458 73218
rect 5458 73166 5460 73218
rect 5404 73164 5460 73166
rect 68460 73052 68516 73108
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 3836 72156 3892 72212
rect 3948 72322 4004 72324
rect 3948 72270 3950 72322
rect 3950 72270 4002 72322
rect 4002 72270 4004 72322
rect 3948 72268 4004 72270
rect 3612 71708 3668 71764
rect 3724 71148 3780 71204
rect 3836 70924 3892 70980
rect 3724 70754 3780 70756
rect 3724 70702 3726 70754
rect 3726 70702 3778 70754
rect 3778 70702 3780 70754
rect 3724 70700 3780 70702
rect 3724 70306 3780 70308
rect 3724 70254 3726 70306
rect 3726 70254 3778 70306
rect 3778 70254 3780 70306
rect 3724 70252 3780 70254
rect 3724 68684 3780 68740
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 4844 71596 4900 71652
rect 5404 71650 5460 71652
rect 5404 71598 5406 71650
rect 5406 71598 5458 71650
rect 5458 71598 5460 71650
rect 5404 71596 5460 71598
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 3948 70252 4004 70308
rect 4060 69916 4116 69972
rect 3836 68572 3892 68628
rect 1708 67004 1764 67060
rect 2156 67004 2212 67060
rect 2044 65996 2100 66052
rect 1820 65324 1876 65380
rect 1820 63084 1876 63140
rect 1932 64652 1988 64708
rect 3948 68460 4004 68516
rect 2268 65772 2324 65828
rect 3388 65436 3444 65492
rect 2156 65100 2212 65156
rect 3388 65100 3444 65156
rect 2044 64428 2100 64484
rect 3724 67058 3780 67060
rect 3724 67006 3726 67058
rect 3726 67006 3778 67058
rect 3778 67006 3780 67058
rect 3724 67004 3780 67006
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 66780 69356 66836 69412
rect 4172 69298 4228 69300
rect 4172 69246 4174 69298
rect 4174 69246 4226 69298
rect 4226 69246 4228 69298
rect 4172 69244 4228 69246
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 5292 68348 5348 68404
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 4172 67730 4228 67732
rect 4172 67678 4174 67730
rect 4174 67678 4226 67730
rect 4226 67678 4228 67730
rect 4172 67676 4228 67678
rect 4060 67564 4116 67620
rect 3836 66892 3892 66948
rect 3612 66108 3668 66164
rect 3724 66050 3780 66052
rect 3724 65998 3726 66050
rect 3726 65998 3778 66050
rect 3778 65998 3780 66050
rect 3724 65996 3780 65998
rect 3724 65378 3780 65380
rect 3724 65326 3726 65378
rect 3726 65326 3778 65378
rect 3778 65326 3780 65378
rect 3724 65324 3780 65326
rect 3500 64540 3556 64596
rect 1932 62636 1988 62692
rect 2044 64204 2100 64260
rect 1932 62466 1988 62468
rect 1932 62414 1934 62466
rect 1934 62414 1986 62466
rect 1986 62414 1988 62466
rect 1932 62412 1988 62414
rect 3724 64204 3780 64260
rect 2044 61740 2100 61796
rect 2156 62860 2212 62916
rect 1820 60396 1876 60452
rect 2044 61292 2100 61348
rect 3276 61682 3332 61684
rect 3276 61630 3278 61682
rect 3278 61630 3330 61682
rect 3330 61630 3332 61682
rect 3276 61628 3332 61630
rect 2156 61068 2212 61124
rect 3500 62076 3556 62132
rect 3948 63756 4004 63812
rect 3724 62972 3780 63028
rect 3724 62466 3780 62468
rect 3724 62414 3726 62466
rect 3726 62414 3778 62466
rect 3778 62414 3780 62466
rect 3724 62412 3780 62414
rect 3612 61404 3668 61460
rect 3724 61346 3780 61348
rect 3724 61294 3726 61346
rect 3726 61294 3778 61346
rect 3778 61294 3780 61346
rect 3724 61292 3780 61294
rect 2044 59724 2100 59780
rect 2156 60620 2212 60676
rect 1932 59330 1988 59332
rect 1932 59278 1934 59330
rect 1934 59278 1986 59330
rect 1986 59278 1988 59330
rect 1932 59276 1988 59278
rect 2156 58380 2212 58436
rect 2268 59724 2324 59780
rect 2044 58156 2100 58212
rect 1820 57036 1876 57092
rect 1932 57484 1988 57540
rect 1820 56140 1876 56196
rect 3500 58716 3556 58772
rect 3724 60674 3780 60676
rect 3724 60622 3726 60674
rect 3726 60622 3778 60674
rect 3778 60622 3780 60674
rect 3724 60620 3780 60622
rect 3836 59948 3892 60004
rect 3724 59276 3780 59332
rect 3612 58604 3668 58660
rect 3948 59052 4004 59108
rect 2268 57708 2324 57764
rect 2044 56364 2100 56420
rect 2268 56754 2324 56756
rect 2268 56702 2270 56754
rect 2270 56702 2322 56754
rect 2322 56702 2324 56754
rect 2268 56700 2324 56702
rect 1932 55692 1988 55748
rect 3724 57538 3780 57540
rect 3724 57486 3726 57538
rect 3726 57486 3778 57538
rect 3778 57486 3780 57538
rect 3724 57484 3780 57486
rect 3724 57036 3780 57092
rect 3836 56812 3892 56868
rect 2268 56194 2324 56196
rect 2268 56142 2270 56194
rect 2270 56142 2322 56194
rect 2322 56142 2324 56194
rect 2268 56140 2324 56142
rect 2156 55468 2212 55524
rect 3276 55410 3332 55412
rect 3276 55358 3278 55410
rect 3278 55358 3330 55410
rect 3330 55358 3332 55410
rect 3276 55356 3332 55358
rect 1820 54348 1876 54404
rect 2044 55020 2100 55076
rect 2044 53788 2100 53844
rect 2156 54684 2212 54740
rect 2044 53452 2100 53508
rect 1932 52780 1988 52836
rect 3500 55132 3556 55188
rect 3388 54572 3444 54628
rect 3724 56754 3780 56756
rect 3724 56702 3726 56754
rect 3726 56702 3778 56754
rect 3778 56702 3780 56754
rect 3724 56700 3780 56702
rect 3724 56194 3780 56196
rect 3724 56142 3726 56194
rect 3726 56142 3778 56194
rect 3778 56142 3780 56194
rect 3724 56140 3780 56142
rect 64876 67900 64932 67956
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 63532 67058 63588 67060
rect 63532 67006 63534 67058
rect 63534 67006 63586 67058
rect 63586 67006 63588 67058
rect 63532 67004 63588 67006
rect 63420 66946 63476 66948
rect 63420 66894 63422 66946
rect 63422 66894 63474 66946
rect 63474 66894 63476 66946
rect 63420 66892 63476 66894
rect 63980 66946 64036 66948
rect 63980 66894 63982 66946
rect 63982 66894 64034 66946
rect 64034 66894 64036 66946
rect 63980 66892 64036 66894
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 67116 68514 67172 68516
rect 67116 68462 67118 68514
rect 67118 68462 67170 68514
rect 67170 68462 67172 68514
rect 67116 68460 67172 68462
rect 67676 68514 67732 68516
rect 67676 68462 67678 68514
rect 67678 68462 67730 68514
rect 67730 68462 67732 68514
rect 67676 68460 67732 68462
rect 69356 72434 69412 72436
rect 69356 72382 69358 72434
rect 69358 72382 69410 72434
rect 69410 72382 69412 72434
rect 69356 72380 69412 72382
rect 68572 69468 68628 69524
rect 67900 68124 67956 68180
rect 66332 67618 66388 67620
rect 66332 67566 66334 67618
rect 66334 67566 66386 67618
rect 66386 67566 66388 67618
rect 66332 67564 66388 67566
rect 67228 67564 67284 67620
rect 63308 66162 63364 66164
rect 63308 66110 63310 66162
rect 63310 66110 63362 66162
rect 63362 66110 63364 66162
rect 63308 66108 63364 66110
rect 63868 66162 63924 66164
rect 63868 66110 63870 66162
rect 63870 66110 63922 66162
rect 63922 66110 63924 66162
rect 63868 66108 63924 66110
rect 63420 66050 63476 66052
rect 63420 65998 63422 66050
rect 63422 65998 63474 66050
rect 63474 65998 63476 66050
rect 63420 65996 63476 65998
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 62076 65548 62132 65604
rect 4284 65324 4340 65380
rect 4956 65436 5012 65492
rect 4284 65100 4340 65156
rect 4172 64706 4228 64708
rect 4172 64654 4174 64706
rect 4174 64654 4226 64706
rect 4226 64654 4228 64706
rect 4172 64652 4228 64654
rect 4172 62914 4228 62916
rect 4172 62862 4174 62914
rect 4174 62862 4226 62914
rect 4226 62862 4228 62914
rect 4172 62860 4228 62862
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 65884 67058 65940 67060
rect 65884 67006 65886 67058
rect 65886 67006 65938 67058
rect 65938 67006 65940 67058
rect 65884 67004 65940 67006
rect 66108 66780 66164 66836
rect 67452 67170 67508 67172
rect 67452 67118 67454 67170
rect 67454 67118 67506 67170
rect 67506 67118 67508 67170
rect 67452 67116 67508 67118
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 65772 66220 65828 66276
rect 65884 66444 65940 66500
rect 66892 66386 66948 66388
rect 66892 66334 66894 66386
rect 66894 66334 66946 66386
rect 66946 66334 66948 66386
rect 66892 66332 66948 66334
rect 67676 67004 67732 67060
rect 67452 66332 67508 66388
rect 67564 66892 67620 66948
rect 65772 66050 65828 66052
rect 65772 65998 65774 66050
rect 65774 65998 65826 66050
rect 65826 65998 65828 66050
rect 65772 65996 65828 65998
rect 67004 66220 67060 66276
rect 65436 65436 65492 65492
rect 61964 65378 62020 65380
rect 61964 65326 61966 65378
rect 61966 65326 62018 65378
rect 62018 65326 62020 65378
rect 61964 65324 62020 65326
rect 62524 65378 62580 65380
rect 62524 65326 62526 65378
rect 62526 65326 62578 65378
rect 62578 65326 62580 65378
rect 62524 65324 62580 65326
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 65436 64876 65492 64932
rect 65884 65602 65940 65604
rect 65884 65550 65886 65602
rect 65886 65550 65938 65602
rect 65938 65550 65940 65602
rect 65884 65548 65940 65550
rect 66108 65490 66164 65492
rect 66108 65438 66110 65490
rect 66110 65438 66162 65490
rect 66162 65438 66164 65490
rect 66108 65436 66164 65438
rect 66668 65436 66724 65492
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 64652 64764 64708 64820
rect 63756 64706 63812 64708
rect 63756 64654 63758 64706
rect 63758 64654 63810 64706
rect 63810 64654 63812 64706
rect 63756 64652 63812 64654
rect 64316 64706 64372 64708
rect 64316 64654 64318 64706
rect 64318 64654 64370 64706
rect 64370 64654 64372 64706
rect 64316 64652 64372 64654
rect 60732 64594 60788 64596
rect 60732 64542 60734 64594
rect 60734 64542 60786 64594
rect 60786 64542 60788 64594
rect 60732 64540 60788 64542
rect 61740 64594 61796 64596
rect 61740 64542 61742 64594
rect 61742 64542 61794 64594
rect 61794 64542 61796 64594
rect 61740 64540 61796 64542
rect 61852 64482 61908 64484
rect 61852 64430 61854 64482
rect 61854 64430 61906 64482
rect 61906 64430 61908 64482
rect 61852 64428 61908 64430
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 61740 64316 61796 64372
rect 4956 63868 5012 63924
rect 59052 64092 59108 64148
rect 5292 63810 5348 63812
rect 5292 63758 5294 63810
rect 5294 63758 5346 63810
rect 5346 63758 5348 63810
rect 5292 63756 5348 63758
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 4284 62188 4340 62244
rect 4844 62076 4900 62132
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 58492 61628 58548 61684
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 61180 64034 61236 64036
rect 61180 63982 61182 64034
rect 61182 63982 61234 64034
rect 61234 63982 61236 64034
rect 61180 63980 61236 63982
rect 61068 63922 61124 63924
rect 61068 63870 61070 63922
rect 61070 63870 61122 63922
rect 61122 63870 61124 63922
rect 61068 63868 61124 63870
rect 61628 63922 61684 63924
rect 61628 63870 61630 63922
rect 61630 63870 61682 63922
rect 61682 63870 61684 63922
rect 61628 63868 61684 63870
rect 59276 63756 59332 63812
rect 59276 63250 59332 63252
rect 59276 63198 59278 63250
rect 59278 63198 59330 63250
rect 59330 63198 59332 63250
rect 59276 63196 59332 63198
rect 59836 63250 59892 63252
rect 59836 63198 59838 63250
rect 59838 63198 59890 63250
rect 59890 63198 59892 63250
rect 59836 63196 59892 63198
rect 61404 63026 61460 63028
rect 61404 62974 61406 63026
rect 61406 62974 61458 63026
rect 61458 62974 61460 63026
rect 61404 62972 61460 62974
rect 59388 62914 59444 62916
rect 59388 62862 59390 62914
rect 59390 62862 59442 62914
rect 59442 62862 59444 62914
rect 59388 62860 59444 62862
rect 61516 62524 61572 62580
rect 62300 64092 62356 64148
rect 62300 63922 62356 63924
rect 62300 63870 62302 63922
rect 62302 63870 62354 63922
rect 62354 63870 62356 63922
rect 62300 63868 62356 63870
rect 63532 64034 63588 64036
rect 63532 63982 63534 64034
rect 63534 63982 63586 64034
rect 63586 63982 63588 64034
rect 63532 63980 63588 63982
rect 62524 63756 62580 63812
rect 61964 63026 62020 63028
rect 61964 62974 61966 63026
rect 61966 62974 62018 63026
rect 62018 62974 62020 63026
rect 61964 62972 62020 62974
rect 59724 62354 59780 62356
rect 59724 62302 59726 62354
rect 59726 62302 59778 62354
rect 59778 62302 59780 62354
rect 59724 62300 59780 62302
rect 63756 63810 63812 63812
rect 63756 63758 63758 63810
rect 63758 63758 63810 63810
rect 63810 63758 63812 63810
rect 63756 63756 63812 63758
rect 65100 64204 65156 64260
rect 62748 62578 62804 62580
rect 62748 62526 62750 62578
rect 62750 62526 62802 62578
rect 62802 62526 62804 62578
rect 62748 62524 62804 62526
rect 63196 62524 63252 62580
rect 59612 62242 59668 62244
rect 59612 62190 59614 62242
rect 59614 62190 59666 62242
rect 59666 62190 59668 62242
rect 59612 62188 59668 62190
rect 60172 62242 60228 62244
rect 60172 62190 60174 62242
rect 60174 62190 60226 62242
rect 60226 62190 60228 62242
rect 60172 62188 60228 62190
rect 61740 62242 61796 62244
rect 61740 62190 61742 62242
rect 61742 62190 61794 62242
rect 61794 62190 61796 62242
rect 61740 62188 61796 62190
rect 62300 62242 62356 62244
rect 62300 62190 62302 62242
rect 62302 62190 62354 62242
rect 62354 62190 62356 62242
rect 62300 62188 62356 62190
rect 4844 60844 4900 60900
rect 57596 60786 57652 60788
rect 57596 60734 57598 60786
rect 57598 60734 57650 60786
rect 57650 60734 57652 60786
rect 57596 60732 57652 60734
rect 57484 60674 57540 60676
rect 57484 60622 57486 60674
rect 57486 60622 57538 60674
rect 57538 60622 57540 60674
rect 57484 60620 57540 60622
rect 58044 60674 58100 60676
rect 58044 60622 58046 60674
rect 58046 60622 58098 60674
rect 58098 60622 58100 60674
rect 58044 60620 58100 60622
rect 57148 60508 57204 60564
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 4172 59778 4228 59780
rect 4172 59726 4174 59778
rect 4174 59726 4226 59778
rect 4226 59726 4228 59778
rect 4172 59724 4228 59726
rect 59836 61346 59892 61348
rect 59836 61294 59838 61346
rect 59838 61294 59890 61346
rect 59890 61294 59892 61346
rect 59836 61292 59892 61294
rect 60284 61292 60340 61348
rect 61516 61292 61572 61348
rect 60396 60956 60452 61012
rect 59052 60508 59108 60564
rect 60732 60898 60788 60900
rect 60732 60846 60734 60898
rect 60734 60846 60786 60898
rect 60786 60846 60788 60898
rect 60732 60844 60788 60846
rect 61068 60844 61124 60900
rect 60956 60786 61012 60788
rect 60956 60734 60958 60786
rect 60958 60734 61010 60786
rect 61010 60734 61012 60786
rect 60956 60732 61012 60734
rect 59724 60620 59780 60676
rect 60396 60620 60452 60676
rect 59388 60508 59444 60564
rect 59948 60060 60004 60116
rect 57820 59948 57876 60004
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 4476 58826 4532 58828
rect 4284 58716 4340 58772
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 4172 58210 4228 58212
rect 4172 58158 4174 58210
rect 4174 58158 4226 58210
rect 4226 58158 4228 58210
rect 4172 58156 4228 58158
rect 4284 57596 4340 57652
rect 4956 58604 5012 58660
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 5292 58156 5348 58212
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 54572 57650 54628 57652
rect 54572 57598 54574 57650
rect 54574 57598 54626 57650
rect 54626 57598 54628 57650
rect 54572 57596 54628 57598
rect 55132 57650 55188 57652
rect 55132 57598 55134 57650
rect 55134 57598 55186 57650
rect 55186 57598 55188 57650
rect 55132 57596 55188 57598
rect 4956 57484 5012 57540
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 4620 57036 4676 57092
rect 55244 56812 55300 56868
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 53228 56082 53284 56084
rect 53228 56030 53230 56082
rect 53230 56030 53282 56082
rect 53282 56030 53284 56082
rect 53228 56028 53284 56030
rect 4620 55916 4676 55972
rect 53116 55970 53172 55972
rect 53116 55918 53118 55970
rect 53118 55918 53170 55970
rect 53170 55918 53172 55970
rect 53116 55916 53172 55918
rect 53676 55970 53732 55972
rect 53676 55918 53678 55970
rect 53678 55918 53730 55970
rect 53730 55918 53732 55970
rect 53676 55916 53732 55918
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 3948 55356 4004 55412
rect 3724 55074 3780 55076
rect 3724 55022 3726 55074
rect 3726 55022 3778 55074
rect 3778 55022 3780 55074
rect 3724 55020 3780 55022
rect 3724 54738 3780 54740
rect 3724 54686 3726 54738
rect 3726 54686 3778 54738
rect 3778 54686 3780 54738
rect 3724 54684 3780 54686
rect 3612 54460 3668 54516
rect 3388 53676 3444 53732
rect 2156 53004 2212 53060
rect 3724 53506 3780 53508
rect 3724 53454 3726 53506
rect 3726 53454 3778 53506
rect 3778 53454 3780 53506
rect 3724 53452 3780 53454
rect 3500 52892 3556 52948
rect 3724 52834 3780 52836
rect 3724 52782 3726 52834
rect 3726 52782 3778 52834
rect 3778 52782 3780 52834
rect 3724 52780 3780 52782
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 3948 52780 4004 52836
rect 3388 52668 3444 52724
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 2044 52332 2100 52388
rect 1932 51660 1988 51716
rect 3388 51996 3444 52052
rect 2044 51884 2100 51940
rect 3724 51884 3780 51940
rect 2044 50988 2100 51044
rect 2156 51212 2212 51268
rect 1932 50540 1988 50596
rect 2156 50428 2212 50484
rect 1932 49756 1988 49812
rect 3724 51266 3780 51268
rect 3724 51214 3726 51266
rect 3726 51214 3778 51266
rect 3778 51214 3780 51266
rect 3724 51212 3780 51214
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 54460 55356 54516 55412
rect 52332 55244 52388 55300
rect 50764 55186 50820 55188
rect 50764 55134 50766 55186
rect 50766 55134 50818 55186
rect 50818 55134 50820 55186
rect 50764 55132 50820 55134
rect 50652 55020 50708 55076
rect 51212 55074 51268 55076
rect 51212 55022 51214 55074
rect 51214 55022 51266 55074
rect 51266 55022 51268 55074
rect 51212 55020 51268 55022
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 52220 54626 52276 54628
rect 52220 54574 52222 54626
rect 52222 54574 52274 54626
rect 52274 54574 52276 54626
rect 52220 54572 52276 54574
rect 51548 54514 51604 54516
rect 51548 54462 51550 54514
rect 51550 54462 51602 54514
rect 51602 54462 51604 54514
rect 51548 54460 51604 54462
rect 52108 54514 52164 54516
rect 52108 54462 52110 54514
rect 52110 54462 52162 54514
rect 52162 54462 52164 54514
rect 52108 54460 52164 54462
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 54236 55298 54292 55300
rect 54236 55246 54238 55298
rect 54238 55246 54290 55298
rect 54290 55246 54292 55298
rect 54236 55244 54292 55246
rect 55580 56082 55636 56084
rect 55580 56030 55582 56082
rect 55582 56030 55634 56082
rect 55634 56030 55636 56082
rect 55580 56028 55636 56030
rect 54572 55244 54628 55300
rect 53900 54684 53956 54740
rect 52780 54402 52836 54404
rect 52780 54350 52782 54402
rect 52782 54350 52834 54402
rect 52834 54350 52836 54402
rect 52780 54348 52836 54350
rect 53340 54402 53396 54404
rect 53340 54350 53342 54402
rect 53342 54350 53394 54402
rect 53394 54350 53396 54402
rect 53340 54348 53396 54350
rect 48188 53676 48244 53732
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 47740 52946 47796 52948
rect 47740 52894 47742 52946
rect 47742 52894 47794 52946
rect 47794 52894 47796 52946
rect 47740 52892 47796 52894
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 55020 55356 55076 55412
rect 54908 54626 54964 54628
rect 54908 54574 54910 54626
rect 54910 54574 54962 54626
rect 54962 54574 54964 54626
rect 54908 54572 54964 54574
rect 55468 55186 55524 55188
rect 55468 55134 55470 55186
rect 55470 55134 55522 55186
rect 55522 55134 55524 55186
rect 55468 55132 55524 55134
rect 54796 54402 54852 54404
rect 54796 54350 54798 54402
rect 54798 54350 54850 54402
rect 54850 54350 54852 54402
rect 54796 54348 54852 54350
rect 54684 53900 54740 53956
rect 52892 53676 52948 53732
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 48300 52946 48356 52948
rect 48300 52894 48302 52946
rect 48302 52894 48354 52946
rect 48354 52894 48356 52946
rect 48300 52892 48356 52894
rect 54684 53730 54740 53732
rect 54684 53678 54686 53730
rect 54686 53678 54738 53730
rect 54738 53678 54740 53730
rect 54684 53676 54740 53678
rect 50540 52946 50596 52948
rect 50540 52894 50542 52946
rect 50542 52894 50594 52946
rect 50594 52894 50596 52946
rect 50540 52892 50596 52894
rect 50428 52834 50484 52836
rect 50428 52782 50430 52834
rect 50430 52782 50482 52834
rect 50482 52782 50484 52834
rect 50428 52780 50484 52782
rect 50988 52834 51044 52836
rect 50988 52782 50990 52834
rect 50990 52782 51042 52834
rect 51042 52782 51044 52834
rect 50988 52780 51044 52782
rect 48300 52274 48356 52276
rect 48300 52222 48302 52274
rect 48302 52222 48354 52274
rect 48354 52222 48356 52274
rect 48300 52220 48356 52222
rect 48412 51938 48468 51940
rect 48412 51886 48414 51938
rect 48414 51886 48466 51938
rect 48466 51886 48468 51938
rect 48412 51884 48468 51886
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 49532 52668 49588 52724
rect 48860 52274 48916 52276
rect 48860 52222 48862 52274
rect 48862 52222 48914 52274
rect 48914 52222 48916 52274
rect 48860 52220 48916 52222
rect 48524 51436 48580 51492
rect 48972 51996 49028 52052
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 4956 50652 5012 50708
rect 52332 52780 52388 52836
rect 52668 52274 52724 52276
rect 52668 52222 52670 52274
rect 52670 52222 52722 52274
rect 52722 52222 52724 52274
rect 52668 52220 52724 52222
rect 49644 51324 49700 51380
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 52220 51938 52276 51940
rect 52220 51886 52222 51938
rect 52222 51886 52274 51938
rect 52274 51886 52276 51938
rect 52220 51884 52276 51886
rect 52108 51772 52164 51828
rect 51884 51602 51940 51604
rect 51884 51550 51886 51602
rect 51886 51550 51938 51602
rect 51938 51550 51940 51602
rect 51884 51548 51940 51550
rect 52108 51324 52164 51380
rect 52556 52108 52612 52164
rect 52444 51772 52500 51828
rect 3724 50594 3780 50596
rect 3724 50542 3726 50594
rect 3726 50542 3778 50594
rect 3778 50542 3780 50594
rect 3724 50540 3780 50542
rect 49532 50482 49588 50484
rect 49532 50430 49534 50482
rect 49534 50430 49586 50482
rect 49586 50430 49588 50482
rect 49532 50428 49588 50430
rect 50652 50482 50708 50484
rect 50652 50430 50654 50482
rect 50654 50430 50706 50482
rect 50706 50430 50708 50482
rect 50652 50428 50708 50430
rect 50428 50316 50484 50372
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 3612 49868 3668 49924
rect 46732 49922 46788 49924
rect 46732 49870 46734 49922
rect 46734 49870 46786 49922
rect 46786 49870 46788 49922
rect 46732 49868 46788 49870
rect 3500 49756 3556 49812
rect 46620 49810 46676 49812
rect 46620 49758 46622 49810
rect 46622 49758 46674 49810
rect 46674 49758 46676 49810
rect 46620 49756 46676 49758
rect 47180 49810 47236 49812
rect 47180 49758 47182 49810
rect 47182 49758 47234 49810
rect 47234 49758 47236 49810
rect 47180 49756 47236 49758
rect 49420 49756 49476 49812
rect 2044 49644 2100 49700
rect 3724 49698 3780 49700
rect 3724 49646 3726 49698
rect 3726 49646 3778 49698
rect 3778 49646 3780 49698
rect 3724 49644 3780 49646
rect 48188 49698 48244 49700
rect 48188 49646 48190 49698
rect 48190 49646 48242 49698
rect 48242 49646 48244 49698
rect 48188 49644 48244 49646
rect 48748 49698 48804 49700
rect 48748 49646 48750 49698
rect 48750 49646 48802 49698
rect 48802 49646 48804 49698
rect 48748 49644 48804 49646
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 3388 49196 3444 49252
rect 48076 49196 48132 49252
rect 3276 49138 3332 49140
rect 3276 49086 3278 49138
rect 3278 49086 3330 49138
rect 3330 49086 3332 49138
rect 3276 49084 3332 49086
rect 2044 48972 2100 49028
rect 1932 48748 1988 48804
rect 4172 48802 4228 48804
rect 4172 48750 4174 48802
rect 4174 48750 4226 48802
rect 4226 48750 4228 48802
rect 4172 48748 4228 48750
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 1932 48300 1988 48356
rect 3724 47628 3780 47684
rect 2044 46956 2100 47012
rect 3052 46674 3108 46676
rect 3052 46622 3054 46674
rect 3054 46622 3106 46674
rect 3106 46622 3108 46674
rect 3052 46620 3108 46622
rect 3612 46620 3668 46676
rect 1932 46284 1988 46340
rect 2044 45612 2100 45668
rect 3500 45276 3556 45332
rect 48412 49196 48468 49252
rect 50428 49922 50484 49924
rect 50428 49870 50430 49922
rect 50430 49870 50482 49922
rect 50482 49870 50484 49922
rect 50428 49868 50484 49870
rect 48524 48748 48580 48804
rect 48300 48188 48356 48244
rect 4844 48076 4900 48132
rect 5404 48130 5460 48132
rect 5404 48078 5406 48130
rect 5406 48078 5458 48130
rect 5458 48078 5460 48130
rect 5404 48076 5460 48078
rect 47068 48076 47124 48132
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 47404 47346 47460 47348
rect 47404 47294 47406 47346
rect 47406 47294 47458 47346
rect 47458 47294 47460 47346
rect 47404 47292 47460 47294
rect 50092 49756 50148 49812
rect 49644 48802 49700 48804
rect 49644 48750 49646 48802
rect 49646 48750 49698 48802
rect 49698 48750 49700 48802
rect 49644 48748 49700 48750
rect 49868 48242 49924 48244
rect 49868 48190 49870 48242
rect 49870 48190 49922 48242
rect 49922 48190 49924 48242
rect 49868 48188 49924 48190
rect 47740 47292 47796 47348
rect 48076 47346 48132 47348
rect 48076 47294 48078 47346
rect 48078 47294 48130 47346
rect 48130 47294 48132 47346
rect 48076 47292 48132 47294
rect 48860 47292 48916 47348
rect 48412 47234 48468 47236
rect 48412 47182 48414 47234
rect 48414 47182 48466 47234
rect 48466 47182 48468 47234
rect 48412 47180 48468 47182
rect 49644 47346 49700 47348
rect 49644 47294 49646 47346
rect 49646 47294 49698 47346
rect 49698 47294 49700 47346
rect 49644 47292 49700 47294
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 3836 46732 3892 46788
rect 46396 46786 46452 46788
rect 46396 46734 46398 46786
rect 46398 46734 46450 46786
rect 46450 46734 46452 46786
rect 46396 46732 46452 46734
rect 47740 46786 47796 46788
rect 47740 46734 47742 46786
rect 47742 46734 47794 46786
rect 47794 46734 47796 46786
rect 47740 46732 47796 46734
rect 45948 46674 46004 46676
rect 45948 46622 45950 46674
rect 45950 46622 46002 46674
rect 46002 46622 46004 46674
rect 45948 46620 46004 46622
rect 46732 46674 46788 46676
rect 46732 46622 46734 46674
rect 46734 46622 46786 46674
rect 46786 46622 46788 46674
rect 46732 46620 46788 46622
rect 47516 46674 47572 46676
rect 47516 46622 47518 46674
rect 47518 46622 47570 46674
rect 47570 46622 47572 46674
rect 47516 46620 47572 46622
rect 48188 46620 48244 46676
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 46060 45890 46116 45892
rect 46060 45838 46062 45890
rect 46062 45838 46114 45890
rect 46114 45838 46116 45890
rect 46060 45836 46116 45838
rect 46956 45890 47012 45892
rect 46956 45838 46958 45890
rect 46958 45838 47010 45890
rect 47010 45838 47012 45890
rect 46956 45836 47012 45838
rect 47740 45836 47796 45892
rect 47180 45778 47236 45780
rect 47180 45726 47182 45778
rect 47182 45726 47234 45778
rect 47234 45726 47236 45778
rect 47180 45724 47236 45726
rect 3724 45612 3780 45668
rect 45724 45666 45780 45668
rect 45724 45614 45726 45666
rect 45726 45614 45778 45666
rect 45778 45614 45780 45666
rect 45724 45612 45780 45614
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 45612 45500 45668 45556
rect 44380 45330 44436 45332
rect 44380 45278 44382 45330
rect 44382 45278 44434 45330
rect 44434 45278 44436 45330
rect 44380 45276 44436 45278
rect 3612 45164 3668 45220
rect 46172 45218 46228 45220
rect 46172 45166 46174 45218
rect 46174 45166 46226 45218
rect 46226 45166 46228 45218
rect 46172 45164 46228 45166
rect 47404 45218 47460 45220
rect 47404 45166 47406 45218
rect 47406 45166 47458 45218
rect 47458 45166 47460 45218
rect 47404 45164 47460 45166
rect 1932 44940 1988 44996
rect 43932 45106 43988 45108
rect 43932 45054 43934 45106
rect 43934 45054 43986 45106
rect 43986 45054 43988 45106
rect 43932 45052 43988 45054
rect 44716 45106 44772 45108
rect 44716 45054 44718 45106
rect 44718 45054 44770 45106
rect 44770 45054 44772 45106
rect 44716 45052 44772 45054
rect 45388 45106 45444 45108
rect 45388 45054 45390 45106
rect 45390 45054 45442 45106
rect 45442 45054 45444 45106
rect 45388 45052 45444 45054
rect 3052 44940 3108 44996
rect 3612 44994 3668 44996
rect 3612 44942 3614 44994
rect 3614 44942 3666 44994
rect 3666 44942 3668 44994
rect 3612 44940 3668 44942
rect 43708 44940 43764 44996
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 2044 44268 2100 44324
rect 46508 45106 46564 45108
rect 46508 45054 46510 45106
rect 46510 45054 46562 45106
rect 46562 45054 46564 45106
rect 46508 45052 46564 45054
rect 47180 45106 47236 45108
rect 47180 45054 47182 45106
rect 47182 45054 47234 45106
rect 47234 45054 47236 45106
rect 47180 45052 47236 45054
rect 45388 44492 45444 44548
rect 46732 44492 46788 44548
rect 44044 44210 44100 44212
rect 44044 44158 44046 44210
rect 44046 44158 44098 44210
rect 44098 44158 44100 44210
rect 44044 44156 44100 44158
rect 44604 44210 44660 44212
rect 44604 44158 44606 44210
rect 44606 44158 44658 44210
rect 44658 44158 44660 44210
rect 44604 44156 44660 44158
rect 45500 44210 45556 44212
rect 45500 44158 45502 44210
rect 45502 44158 45554 44210
rect 45554 44158 45556 44210
rect 45500 44156 45556 44158
rect 46396 44210 46452 44212
rect 46396 44158 46398 44210
rect 46398 44158 46450 44210
rect 46450 44158 46452 44210
rect 46396 44156 46452 44158
rect 3052 44044 3108 44100
rect 3500 44098 3556 44100
rect 3500 44046 3502 44098
rect 3502 44046 3554 44098
rect 3554 44046 3556 44098
rect 3500 44044 3556 44046
rect 43036 44044 43092 44100
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 45836 44098 45892 44100
rect 45836 44046 45838 44098
rect 45838 44046 45890 44098
rect 45890 44046 45892 44098
rect 45836 44044 45892 44046
rect 44492 43762 44548 43764
rect 44492 43710 44494 43762
rect 44494 43710 44546 43762
rect 44546 43710 44548 43762
rect 44492 43708 44548 43710
rect 1932 43596 1988 43652
rect 42588 43538 42644 43540
rect 42588 43486 42590 43538
rect 42590 43486 42642 43538
rect 42642 43486 42644 43538
rect 42588 43484 42644 43486
rect 43372 43538 43428 43540
rect 43372 43486 43374 43538
rect 43374 43486 43426 43538
rect 43426 43486 43428 43538
rect 43372 43484 43428 43486
rect 44268 43538 44324 43540
rect 44268 43486 44270 43538
rect 44270 43486 44322 43538
rect 44322 43486 44324 43538
rect 44268 43484 44324 43486
rect 44940 43484 44996 43540
rect 3052 43372 3108 43428
rect 3612 43426 3668 43428
rect 3612 43374 3614 43426
rect 3614 43374 3666 43426
rect 3666 43374 3668 43426
rect 3612 43372 3668 43374
rect 42364 43372 42420 43428
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 1932 42924 1988 42980
rect 3052 42588 3108 42644
rect 3500 42642 3556 42644
rect 3500 42590 3502 42642
rect 3502 42590 3554 42642
rect 3554 42590 3556 42642
rect 3500 42588 3556 42590
rect 41804 42588 41860 42644
rect 1932 42252 1988 42308
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 42700 42642 42756 42644
rect 42700 42590 42702 42642
rect 42702 42590 42754 42642
rect 42754 42590 42756 42642
rect 42700 42588 42756 42590
rect 43484 42588 43540 42644
rect 41916 42530 41972 42532
rect 41916 42478 41918 42530
rect 41918 42478 41970 42530
rect 41970 42478 41972 42530
rect 41916 42476 41972 42478
rect 43148 42082 43204 42084
rect 43148 42030 43150 42082
rect 43150 42030 43202 42082
rect 43202 42030 43204 42082
rect 43148 42028 43204 42030
rect 3052 41804 3108 41860
rect 3612 41858 3668 41860
rect 3612 41806 3614 41858
rect 3614 41806 3666 41858
rect 3666 41806 3668 41858
rect 3612 41804 3668 41806
rect 41020 41804 41076 41860
rect 1932 41580 1988 41636
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 1932 40908 1988 40964
rect 42140 41804 42196 41860
rect 42924 41804 42980 41860
rect 3052 40908 3108 40964
rect 3500 40962 3556 40964
rect 3500 40910 3502 40962
rect 3502 40910 3554 40962
rect 3554 40910 3556 40962
rect 3500 40908 3556 40910
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 3052 40402 3108 40404
rect 3052 40350 3054 40402
rect 3054 40350 3106 40402
rect 3106 40350 3108 40402
rect 3052 40348 3108 40350
rect 3612 40402 3668 40404
rect 3612 40350 3614 40402
rect 3614 40350 3666 40402
rect 3666 40350 3668 40402
rect 3612 40348 3668 40350
rect 39452 40348 39508 40404
rect 1932 40290 1988 40292
rect 1932 40238 1934 40290
rect 1934 40238 1986 40290
rect 1986 40238 1988 40290
rect 1932 40236 1988 40238
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 1932 39618 1988 39620
rect 1932 39566 1934 39618
rect 1934 39566 1986 39618
rect 1986 39566 1988 39618
rect 1932 39564 1988 39566
rect 3052 39452 3108 39508
rect 3612 39506 3668 39508
rect 3612 39454 3614 39506
rect 3614 39454 3666 39506
rect 3666 39454 3668 39506
rect 3612 39452 3668 39454
rect 38892 39506 38948 39508
rect 38892 39454 38894 39506
rect 38894 39454 38946 39506
rect 38946 39454 38948 39506
rect 38892 39452 38948 39454
rect 38444 39394 38500 39396
rect 38444 39342 38446 39394
rect 38446 39342 38498 39394
rect 38498 39342 38500 39394
rect 38444 39340 38500 39342
rect 39788 39900 39844 39956
rect 40348 40908 40404 40964
rect 40572 40572 40628 40628
rect 41356 40572 41412 40628
rect 41804 40572 41860 40628
rect 40684 40402 40740 40404
rect 40684 40350 40686 40402
rect 40686 40350 40738 40402
rect 40738 40350 40740 40402
rect 40684 40348 40740 40350
rect 41580 40402 41636 40404
rect 41580 40350 41582 40402
rect 41582 40350 41634 40402
rect 41634 40350 41636 40402
rect 41580 40348 41636 40350
rect 40124 39900 40180 39956
rect 40684 39900 40740 39956
rect 39004 39340 39060 39396
rect 39228 39506 39284 39508
rect 39228 39454 39230 39506
rect 39230 39454 39282 39506
rect 39282 39454 39284 39506
rect 39228 39452 39284 39454
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 1932 38946 1988 38948
rect 1932 38894 1934 38946
rect 1934 38894 1986 38946
rect 1986 38894 1988 38946
rect 1932 38892 1988 38894
rect 3052 38834 3108 38836
rect 3052 38782 3054 38834
rect 3054 38782 3106 38834
rect 3106 38782 3108 38834
rect 3052 38780 3108 38782
rect 3612 38834 3668 38836
rect 3612 38782 3614 38834
rect 3614 38782 3666 38834
rect 3666 38782 3668 38834
rect 3612 38780 3668 38782
rect 38332 38780 38388 38836
rect 38668 38834 38724 38836
rect 38668 38782 38670 38834
rect 38670 38782 38722 38834
rect 38722 38782 38724 38834
rect 38668 38780 38724 38782
rect 37884 38722 37940 38724
rect 37884 38670 37886 38722
rect 37886 38670 37938 38722
rect 37938 38670 37940 38722
rect 37884 38668 37940 38670
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 1932 38220 1988 38276
rect 37996 37938 38052 37940
rect 37996 37886 37998 37938
rect 37998 37886 38050 37938
rect 38050 37886 38052 37938
rect 37996 37884 38052 37886
rect 38892 37884 38948 37940
rect 3052 37772 3108 37828
rect 3612 37826 3668 37828
rect 3612 37774 3614 37826
rect 3614 37774 3666 37826
rect 3666 37774 3668 37826
rect 3612 37772 3668 37774
rect 37660 37826 37716 37828
rect 37660 37774 37662 37826
rect 37662 37774 37714 37826
rect 37714 37774 37716 37826
rect 37660 37772 37716 37774
rect 19836 37658 19892 37660
rect 1932 37548 1988 37604
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 36540 37266 36596 37268
rect 36540 37214 36542 37266
rect 36542 37214 36594 37266
rect 36594 37214 36596 37266
rect 36540 37212 36596 37214
rect 3052 36988 3108 37044
rect 3612 36988 3668 37044
rect 38444 37378 38500 37380
rect 38444 37326 38446 37378
rect 38446 37326 38498 37378
rect 38498 37326 38500 37378
rect 38444 37324 38500 37326
rect 36988 36988 37044 37044
rect 37324 37266 37380 37268
rect 37324 37214 37326 37266
rect 37326 37214 37378 37266
rect 37378 37214 37380 37266
rect 37324 37212 37380 37214
rect 1932 36876 1988 36932
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 1932 36204 1988 36260
rect 35868 36370 35924 36372
rect 35868 36318 35870 36370
rect 35870 36318 35922 36370
rect 35922 36318 35924 36370
rect 35868 36316 35924 36318
rect 36540 36316 36596 36372
rect 3052 36204 3108 36260
rect 3612 36258 3668 36260
rect 3612 36206 3614 36258
rect 3614 36206 3666 36258
rect 3666 36206 3668 36258
rect 3612 36204 3668 36206
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 3052 35756 3108 35812
rect 3612 35756 3668 35812
rect 1932 35532 1988 35588
rect 4844 35532 4900 35588
rect 5404 35586 5460 35588
rect 5404 35534 5406 35586
rect 5406 35534 5458 35586
rect 5458 35534 5460 35586
rect 5404 35532 5460 35534
rect 34300 35532 34356 35588
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 3724 34860 3780 34916
rect 33852 34802 33908 34804
rect 33852 34750 33854 34802
rect 33854 34750 33906 34802
rect 33906 34750 33908 34802
rect 33852 34748 33908 34750
rect 34636 34802 34692 34804
rect 34636 34750 34638 34802
rect 34638 34750 34690 34802
rect 34690 34750 34692 34802
rect 34636 34748 34692 34750
rect 3052 34636 3108 34692
rect 4060 34690 4116 34692
rect 4060 34638 4062 34690
rect 4062 34638 4114 34690
rect 4114 34638 4116 34690
rect 4060 34636 4116 34638
rect 34748 34636 34804 34692
rect 36316 36258 36372 36260
rect 36316 36206 36318 36258
rect 36318 36206 36370 36258
rect 36370 36206 36372 36258
rect 36316 36204 36372 36206
rect 35644 35810 35700 35812
rect 35644 35758 35646 35810
rect 35646 35758 35698 35810
rect 35698 35758 35700 35810
rect 35644 35756 35700 35758
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 1932 34242 1988 34244
rect 1932 34190 1934 34242
rect 1934 34190 1986 34242
rect 1986 34190 1988 34242
rect 1932 34188 1988 34190
rect 3052 33964 3108 34020
rect 3612 34018 3668 34020
rect 3612 33966 3614 34018
rect 3614 33966 3666 34018
rect 3666 33966 3668 34018
rect 3612 33964 3668 33966
rect 34076 34130 34132 34132
rect 34076 34078 34078 34130
rect 34078 34078 34130 34130
rect 34130 34078 34132 34130
rect 34076 34076 34132 34078
rect 34860 34130 34916 34132
rect 34860 34078 34862 34130
rect 34862 34078 34914 34130
rect 34914 34078 34916 34130
rect 34860 34076 34916 34078
rect 33740 33964 33796 34020
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 1932 33516 1988 33572
rect 32508 33292 32564 33348
rect 3052 33180 3108 33236
rect 3612 33234 3668 33236
rect 3612 33182 3614 33234
rect 3614 33182 3666 33234
rect 3666 33182 3668 33234
rect 3612 33180 3668 33182
rect 33180 33346 33236 33348
rect 33180 33294 33182 33346
rect 33182 33294 33234 33346
rect 33234 33294 33236 33346
rect 33180 33292 33236 33294
rect 34076 33346 34132 33348
rect 34076 33294 34078 33346
rect 34078 33294 34130 33346
rect 34130 33294 34132 33346
rect 34076 33292 34132 33294
rect 32956 33234 33012 33236
rect 32956 33182 32958 33234
rect 32958 33182 33010 33234
rect 33010 33182 33012 33234
rect 32956 33180 33012 33182
rect 19836 32954 19892 32956
rect 1932 32844 1988 32900
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 31836 32508 31892 32564
rect 3052 32284 3108 32340
rect 3612 32284 3668 32340
rect 1932 32172 1988 32228
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 1932 31500 1988 31556
rect 31164 31612 31220 31668
rect 3052 31500 3108 31556
rect 3612 31554 3668 31556
rect 3612 31502 3614 31554
rect 3614 31502 3666 31554
rect 3666 31502 3668 31554
rect 3612 31500 3668 31502
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 3052 31052 3108 31108
rect 3612 31052 3668 31108
rect 1932 30828 1988 30884
rect 4844 30828 4900 30884
rect 5404 30882 5460 30884
rect 5404 30830 5406 30882
rect 5406 30830 5458 30882
rect 5458 30830 5460 30882
rect 5404 30828 5460 30830
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 3724 30156 3780 30212
rect 28812 30044 28868 30100
rect 3052 29932 3108 29988
rect 29372 30044 29428 30100
rect 29596 30828 29652 30884
rect 29932 30098 29988 30100
rect 29932 30046 29934 30098
rect 29934 30046 29986 30098
rect 29986 30046 29988 30098
rect 29932 30044 29988 30046
rect 4060 29986 4116 29988
rect 4060 29934 4062 29986
rect 4062 29934 4114 29986
rect 4114 29934 4116 29986
rect 4060 29932 4116 29934
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 1932 29538 1988 29540
rect 1932 29486 1934 29538
rect 1934 29486 1986 29538
rect 1986 29486 1988 29538
rect 1932 29484 1988 29486
rect 28476 29426 28532 29428
rect 28476 29374 28478 29426
rect 28478 29374 28530 29426
rect 28530 29374 28532 29426
rect 28476 29372 28532 29374
rect 3052 29260 3108 29316
rect 3612 29314 3668 29316
rect 3612 29262 3614 29314
rect 3614 29262 3666 29314
rect 3666 29262 3668 29314
rect 3612 29260 3668 29262
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 1932 28812 1988 28868
rect 3052 28642 3108 28644
rect 3052 28590 3054 28642
rect 3054 28590 3106 28642
rect 3106 28590 3108 28642
rect 3052 28588 3108 28590
rect 3612 28642 3668 28644
rect 3612 28590 3614 28642
rect 3614 28590 3666 28642
rect 3666 28590 3668 28642
rect 3612 28588 3668 28590
rect 28252 28588 28308 28644
rect 27692 28476 27748 28532
rect 19836 28250 19892 28252
rect 1932 28140 1988 28196
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 27132 27804 27188 27860
rect 3052 27692 3108 27748
rect 3612 27746 3668 27748
rect 3612 27694 3614 27746
rect 3614 27694 3666 27746
rect 3666 27694 3668 27746
rect 3612 27692 3668 27694
rect 1932 27468 1988 27524
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 3052 27074 3108 27076
rect 3052 27022 3054 27074
rect 3054 27022 3106 27074
rect 3106 27022 3108 27074
rect 3052 27020 3108 27022
rect 3612 27074 3668 27076
rect 3612 27022 3614 27074
rect 3614 27022 3666 27074
rect 3666 27022 3668 27074
rect 3612 27020 3668 27022
rect 26908 27020 26964 27076
rect 26460 26962 26516 26964
rect 26460 26910 26462 26962
rect 26462 26910 26514 26962
rect 26514 26910 26516 26962
rect 26460 26908 26516 26910
rect 1932 26796 1988 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 1932 26124 1988 26180
rect 25788 26290 25844 26292
rect 25788 26238 25790 26290
rect 25790 26238 25842 26290
rect 25842 26238 25844 26290
rect 25788 26236 25844 26238
rect 4844 26124 4900 26180
rect 5404 26178 5460 26180
rect 5404 26126 5406 26178
rect 5406 26126 5458 26178
rect 5458 26126 5460 26178
rect 5404 26124 5460 26126
rect 24332 26124 24388 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 3724 25452 3780 25508
rect 3052 25340 3108 25396
rect 4060 25394 4116 25396
rect 4060 25342 4062 25394
rect 4062 25342 4114 25394
rect 4114 25342 4116 25394
rect 4060 25340 4116 25342
rect 2940 25228 2996 25284
rect 3612 25282 3668 25284
rect 3612 25230 3614 25282
rect 3614 25230 3666 25282
rect 3666 25230 3668 25282
rect 3612 25228 3668 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 24668 25116 24724 25172
rect 25564 25506 25620 25508
rect 25564 25454 25566 25506
rect 25566 25454 25618 25506
rect 25618 25454 25620 25506
rect 25564 25452 25620 25454
rect 25228 25394 25284 25396
rect 25228 25342 25230 25394
rect 25230 25342 25282 25394
rect 25282 25342 25284 25394
rect 25228 25340 25284 25342
rect 26572 26290 26628 26292
rect 26572 26238 26574 26290
rect 26574 26238 26626 26290
rect 26626 26238 26628 26290
rect 26572 26236 26628 26238
rect 27580 27692 27636 27748
rect 28588 28530 28644 28532
rect 28588 28478 28590 28530
rect 28590 28478 28642 28530
rect 28642 28478 28644 28530
rect 28588 28476 28644 28478
rect 27804 27858 27860 27860
rect 27804 27806 27806 27858
rect 27806 27806 27858 27858
rect 27858 27806 27860 27858
rect 27804 27804 27860 27806
rect 28588 27858 28644 27860
rect 28588 27806 28590 27858
rect 28590 27806 28642 27858
rect 28642 27806 28644 27858
rect 28588 27804 28644 27806
rect 27244 26962 27300 26964
rect 27244 26910 27246 26962
rect 27246 26910 27298 26962
rect 27298 26910 27300 26962
rect 27244 26908 27300 26910
rect 27020 25788 27076 25844
rect 27132 26236 27188 26292
rect 26460 25506 26516 25508
rect 26460 25454 26462 25506
rect 26462 25454 26514 25506
rect 26514 25454 26516 25506
rect 26460 25452 26516 25454
rect 26236 25228 26292 25284
rect 25004 25116 25060 25172
rect 25900 25116 25956 25172
rect 20044 25060 20100 25062
rect 1932 24834 1988 24836
rect 1932 24782 1934 24834
rect 1934 24782 1986 24834
rect 1986 24782 1988 24834
rect 1932 24780 1988 24782
rect 22764 24722 22820 24724
rect 22764 24670 22766 24722
rect 22766 24670 22818 24722
rect 22818 24670 22820 24722
rect 22764 24668 22820 24670
rect 23100 24722 23156 24724
rect 23100 24670 23102 24722
rect 23102 24670 23154 24722
rect 23154 24670 23156 24722
rect 23100 24668 23156 24670
rect 3052 24444 3108 24500
rect 3612 24444 3668 24500
rect 23996 24722 24052 24724
rect 23996 24670 23998 24722
rect 23998 24670 24050 24722
rect 24050 24670 24052 24722
rect 23996 24668 24052 24670
rect 23660 24444 23716 24500
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 1932 24108 1988 24164
rect 3052 23660 3108 23716
rect 3612 23714 3668 23716
rect 3612 23662 3614 23714
rect 3614 23662 3666 23714
rect 3666 23662 3668 23714
rect 3612 23660 3668 23662
rect 19836 23546 19892 23548
rect 1932 23436 1988 23492
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 3052 22988 3108 23044
rect 3612 23042 3668 23044
rect 3612 22990 3614 23042
rect 3614 22990 3666 23042
rect 3666 22990 3668 23042
rect 3612 22988 3668 22990
rect 22764 23154 22820 23156
rect 22764 23102 22766 23154
rect 22766 23102 22818 23154
rect 22818 23102 22820 23154
rect 22764 23100 22820 23102
rect 23660 23714 23716 23716
rect 23660 23662 23662 23714
rect 23662 23662 23714 23714
rect 23714 23662 23716 23714
rect 23660 23660 23716 23662
rect 23884 23266 23940 23268
rect 23884 23214 23886 23266
rect 23886 23214 23938 23266
rect 23938 23214 23940 23266
rect 23884 23212 23940 23214
rect 23100 23100 23156 23156
rect 23660 23154 23716 23156
rect 23660 23102 23662 23154
rect 23662 23102 23714 23154
rect 23714 23102 23716 23154
rect 23660 23100 23716 23102
rect 22428 22988 22484 23044
rect 1932 22764 1988 22820
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 1932 22092 1988 22148
rect 3052 22092 3108 22148
rect 3612 22146 3668 22148
rect 3612 22094 3614 22146
rect 3614 22094 3666 22146
rect 3666 22094 3668 22146
rect 3612 22092 3668 22094
rect 22092 22146 22148 22148
rect 22092 22094 22094 22146
rect 22094 22094 22146 22146
rect 22146 22094 22148 22146
rect 22092 22092 22148 22094
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 22652 21810 22708 21812
rect 22652 21758 22654 21810
rect 22654 21758 22706 21810
rect 22706 21758 22708 21810
rect 22652 21756 22708 21758
rect 23324 22146 23380 22148
rect 23324 22094 23326 22146
rect 23326 22094 23378 22146
rect 23378 22094 23380 22146
rect 23324 22092 23380 22094
rect 24332 22876 24388 22932
rect 23100 21756 23156 21812
rect 1932 21420 1988 21476
rect 2940 20860 2996 20916
rect 3612 20914 3668 20916
rect 3612 20862 3614 20914
rect 3614 20862 3666 20914
rect 3666 20862 3668 20914
rect 3612 20860 3668 20862
rect 4844 21420 4900 21476
rect 5404 21474 5460 21476
rect 5404 21422 5406 21474
rect 5406 21422 5458 21474
rect 5458 21422 5460 21474
rect 5404 21420 5460 21422
rect 19628 21420 19684 21476
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 3724 20748 3780 20804
rect 3052 20636 3108 20692
rect 4060 20690 4116 20692
rect 4060 20638 4062 20690
rect 4062 20638 4114 20690
rect 4114 20638 4116 20690
rect 4060 20636 4116 20638
rect 22092 21586 22148 21588
rect 22092 21534 22094 21586
rect 22094 21534 22146 21586
rect 22146 21534 22148 21586
rect 22092 21532 22148 21534
rect 23100 21586 23156 21588
rect 23100 21534 23102 21586
rect 23102 21534 23154 21586
rect 23154 21534 23156 21586
rect 23100 21532 23156 21534
rect 21756 20860 21812 20916
rect 20972 20748 21028 20804
rect 21868 20802 21924 20804
rect 21868 20750 21870 20802
rect 21870 20750 21922 20802
rect 21922 20750 21924 20802
rect 21868 20748 21924 20750
rect 22764 20802 22820 20804
rect 22764 20750 22766 20802
rect 22766 20750 22818 20802
rect 22818 20750 22820 20802
rect 22764 20748 22820 20750
rect 21644 20690 21700 20692
rect 21644 20638 21646 20690
rect 21646 20638 21698 20690
rect 21698 20638 21700 20690
rect 21644 20636 21700 20638
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 1932 20130 1988 20132
rect 1932 20078 1934 20130
rect 1934 20078 1986 20130
rect 1986 20078 1988 20130
rect 1932 20076 1988 20078
rect 19516 20018 19572 20020
rect 19516 19966 19518 20018
rect 19518 19966 19570 20018
rect 19570 19966 19572 20018
rect 19516 19964 19572 19966
rect 20300 20018 20356 20020
rect 20300 19966 20302 20018
rect 20302 19966 20354 20018
rect 20354 19966 20356 20018
rect 20300 19964 20356 19966
rect 3052 19852 3108 19908
rect 3612 19906 3668 19908
rect 3612 19854 3614 19906
rect 3614 19854 3666 19906
rect 3666 19854 3668 19906
rect 3612 19852 3668 19854
rect 19628 19852 19684 19908
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 1932 19404 1988 19460
rect 3052 18844 3108 18900
rect 18284 19010 18340 19012
rect 18284 18958 18286 19010
rect 18286 18958 18338 19010
rect 18338 18958 18340 19010
rect 18284 18956 18340 18958
rect 3612 18844 3668 18900
rect 18732 18844 18788 18900
rect 18956 18956 19012 19012
rect 1932 18732 1988 18788
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 3052 18284 3108 18340
rect 3612 18338 3668 18340
rect 3612 18286 3614 18338
rect 3614 18286 3666 18338
rect 3666 18286 3668 18338
rect 3612 18284 3668 18286
rect 1932 18060 1988 18116
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 1932 17388 1988 17444
rect 18620 18284 18676 18340
rect 3052 17276 3108 17332
rect 3612 17276 3668 17332
rect 3052 16940 3108 16996
rect 3612 16940 3668 16996
rect 1932 16716 1988 16772
rect 4844 16882 4900 16884
rect 4844 16830 4846 16882
rect 4846 16830 4898 16882
rect 4898 16830 4900 16882
rect 4844 16828 4900 16830
rect 5404 16882 5460 16884
rect 5404 16830 5406 16882
rect 5406 16830 5458 16882
rect 5458 16830 5460 16882
rect 5404 16828 5460 16830
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 3724 16044 3780 16100
rect 3052 15820 3108 15876
rect 4060 15874 4116 15876
rect 4060 15822 4062 15874
rect 4062 15822 4114 15874
rect 4114 15822 4116 15874
rect 4060 15820 4116 15822
rect 15820 16828 15876 16884
rect 16044 16882 16100 16884
rect 16044 16830 16046 16882
rect 16046 16830 16098 16882
rect 16098 16830 16100 16882
rect 16044 16828 16100 16830
rect 17612 17276 17668 17332
rect 16604 16994 16660 16996
rect 16604 16942 16606 16994
rect 16606 16942 16658 16994
rect 16658 16942 16660 16994
rect 16604 16940 16660 16942
rect 16380 16828 16436 16884
rect 16716 16828 16772 16884
rect 15708 15820 15764 15876
rect 1932 15426 1988 15428
rect 1932 15374 1934 15426
rect 1934 15374 1986 15426
rect 1986 15374 1988 15426
rect 1932 15372 1988 15374
rect 3052 15148 3108 15204
rect 3612 15202 3668 15204
rect 3612 15150 3614 15202
rect 3614 15150 3666 15202
rect 3666 15150 3668 15202
rect 3612 15148 3668 15150
rect 14700 15148 14756 15204
rect 16380 15314 16436 15316
rect 16380 15262 16382 15314
rect 16382 15262 16434 15314
rect 16434 15262 16436 15314
rect 16380 15260 16436 15262
rect 15036 15148 15092 15204
rect 15484 15202 15540 15204
rect 15484 15150 15486 15202
rect 15486 15150 15538 15202
rect 15538 15150 15540 15202
rect 15484 15148 15540 15150
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 1932 14700 1988 14756
rect 3052 14252 3108 14308
rect 3612 14306 3668 14308
rect 3612 14254 3614 14306
rect 3614 14254 3666 14306
rect 3666 14254 3668 14306
rect 3612 14252 3668 14254
rect 14028 14306 14084 14308
rect 14028 14254 14030 14306
rect 14030 14254 14082 14306
rect 14082 14254 14084 14306
rect 14028 14252 14084 14254
rect 14364 14252 14420 14308
rect 14812 14306 14868 14308
rect 14812 14254 14814 14306
rect 14814 14254 14866 14306
rect 14866 14254 14868 14306
rect 14812 14252 14868 14254
rect 1932 14028 1988 14084
rect 3052 13580 3108 13636
rect 3612 13634 3668 13636
rect 3612 13582 3614 13634
rect 3614 13582 3666 13634
rect 3666 13582 3668 13634
rect 3612 13580 3668 13582
rect 12012 13468 12068 13524
rect 1932 13356 1988 13412
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 1932 12684 1988 12740
rect 3052 12684 3108 12740
rect 3612 12738 3668 12740
rect 3612 12686 3614 12738
rect 3614 12686 3666 12738
rect 3666 12686 3668 12738
rect 3612 12684 3668 12686
rect 3052 12236 3108 12292
rect 3612 12236 3668 12292
rect 1932 12012 1988 12068
rect 3052 11452 3108 11508
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4060 11506 4116 11508
rect 4060 11454 4062 11506
rect 4062 11454 4114 11506
rect 4114 11454 4116 11506
rect 4060 11452 4116 11454
rect 3724 11340 3780 11396
rect 13692 13746 13748 13748
rect 13692 13694 13694 13746
rect 13694 13694 13746 13746
rect 13746 13694 13748 13746
rect 13692 13692 13748 13694
rect 14140 13746 14196 13748
rect 14140 13694 14142 13746
rect 14142 13694 14194 13746
rect 14194 13694 14196 13746
rect 14140 13692 14196 13694
rect 13356 13580 13412 13636
rect 12796 13468 12852 13524
rect 14028 13468 14084 13524
rect 12460 12684 12516 12740
rect 12236 12290 12292 12292
rect 12236 12238 12238 12290
rect 12238 12238 12290 12290
rect 12290 12238 12292 12290
rect 12236 12236 12292 12238
rect 12572 12178 12628 12180
rect 12572 12126 12574 12178
rect 12574 12126 12626 12178
rect 12626 12126 12628 12178
rect 12572 12124 12628 12126
rect 11340 11452 11396 11508
rect 13468 12290 13524 12292
rect 13468 12238 13470 12290
rect 13470 12238 13522 12290
rect 13522 12238 13524 12290
rect 13468 12236 13524 12238
rect 12908 12124 12964 12180
rect 13244 12178 13300 12180
rect 13244 12126 13246 12178
rect 13246 12126 13298 12178
rect 13298 12126 13300 12178
rect 13244 12124 13300 12126
rect 13916 12124 13972 12180
rect 11788 11340 11844 11396
rect 12572 11394 12628 11396
rect 12572 11342 12574 11394
rect 12574 11342 12626 11394
rect 12626 11342 12628 11394
rect 12572 11340 12628 11342
rect 4844 11228 4900 11284
rect 10668 11282 10724 11284
rect 10668 11230 10670 11282
rect 10670 11230 10722 11282
rect 10722 11230 10724 11282
rect 10668 11228 10724 11230
rect 1932 10722 1988 10724
rect 1932 10670 1934 10722
rect 1934 10670 1986 10722
rect 1986 10670 1988 10722
rect 1932 10668 1988 10670
rect 3052 10668 3108 10724
rect 10108 10722 10164 10724
rect 10108 10670 10110 10722
rect 10110 10670 10162 10722
rect 10162 10670 10164 10722
rect 10108 10668 10164 10670
rect 11452 10722 11508 10724
rect 11452 10670 11454 10722
rect 11454 10670 11506 10722
rect 11506 10670 11508 10722
rect 11452 10668 11508 10670
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 1932 9996 1988 10052
rect 3052 9660 3108 9716
rect 9436 9714 9492 9716
rect 9436 9662 9438 9714
rect 9438 9662 9490 9714
rect 9490 9662 9492 9714
rect 9436 9660 9492 9662
rect 9660 9660 9716 9716
rect 1932 9324 1988 9380
rect 3052 9100 3108 9156
rect 8652 9154 8708 9156
rect 8652 9102 8654 9154
rect 8654 9102 8706 9154
rect 8706 9102 8708 9154
rect 8652 9100 8708 9102
rect 8988 9042 9044 9044
rect 8988 8990 8990 9042
rect 8990 8990 9042 9042
rect 9042 8990 9044 9042
rect 8988 8988 9044 8990
rect 1932 8652 1988 8708
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 3052 8092 3108 8148
rect 8092 8146 8148 8148
rect 8092 8094 8094 8146
rect 8094 8094 8146 8146
rect 8146 8094 8148 8146
rect 8092 8092 8148 8094
rect 8428 8146 8484 8148
rect 8428 8094 8430 8146
rect 8430 8094 8482 8146
rect 8482 8094 8484 8146
rect 8428 8092 8484 8094
rect 1932 7980 1988 8036
rect 3052 7532 3108 7588
rect 1932 7308 1988 7364
rect 3052 6748 3108 6804
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 3724 6636 3780 6692
rect 7420 7586 7476 7588
rect 7420 7534 7422 7586
rect 7422 7534 7474 7586
rect 7474 7534 7476 7586
rect 7420 7532 7476 7534
rect 8764 7586 8820 7588
rect 8764 7534 8766 7586
rect 8766 7534 8818 7586
rect 8818 7534 8820 7586
rect 8764 7532 8820 7534
rect 6524 6748 6580 6804
rect 6860 6748 6916 6804
rect 7644 7474 7700 7476
rect 7644 7422 7646 7474
rect 7646 7422 7698 7474
rect 7698 7422 7700 7474
rect 7644 7420 7700 7422
rect 4844 6524 4900 6580
rect 5740 6636 5796 6692
rect 1932 6018 1988 6020
rect 1932 5966 1934 6018
rect 1934 5966 1986 6018
rect 1986 5966 1988 6018
rect 1932 5964 1988 5966
rect 3052 5964 3108 6020
rect 4620 6018 4676 6020
rect 4620 5966 4622 6018
rect 4622 5966 4674 6018
rect 4674 5966 4676 6018
rect 4620 5964 4676 5966
rect 1932 5292 1988 5348
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4620 5180 4676 5236
rect 5516 5180 5572 5236
rect 4172 4732 4228 4788
rect 3052 4508 3108 4564
rect 4620 4562 4676 4564
rect 4620 4510 4622 4562
rect 4622 4510 4674 4562
rect 4674 4510 4676 4562
rect 4620 4508 4676 4510
rect 5068 4956 5124 5012
rect 4956 4898 5012 4900
rect 4956 4846 4958 4898
rect 4958 4846 5010 4898
rect 5010 4846 5012 4898
rect 4956 4844 5012 4846
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 5292 4732 5348 4788
rect 3948 3442 4004 3444
rect 3948 3390 3950 3442
rect 3950 3390 4002 3442
rect 4002 3390 4004 3442
rect 3948 3388 4004 3390
rect 6300 6690 6356 6692
rect 6300 6638 6302 6690
rect 6302 6638 6354 6690
rect 6354 6638 6356 6690
rect 6300 6636 6356 6638
rect 6972 6690 7028 6692
rect 6972 6638 6974 6690
rect 6974 6638 7026 6690
rect 7026 6638 7028 6690
rect 6972 6636 7028 6638
rect 7308 6636 7364 6692
rect 6076 6578 6132 6580
rect 6076 6526 6078 6578
rect 6078 6526 6130 6578
rect 6130 6526 6132 6578
rect 6076 6524 6132 6526
rect 6412 5010 6468 5012
rect 6412 4958 6414 5010
rect 6414 4958 6466 5010
rect 6466 4958 6468 5010
rect 6412 4956 6468 4958
rect 6860 4732 6916 4788
rect 7308 5964 7364 6020
rect 6748 4620 6804 4676
rect 5740 3442 5796 3444
rect 5740 3390 5742 3442
rect 5742 3390 5794 3442
rect 5794 3390 5796 3442
rect 5740 3388 5796 3390
rect 8428 7474 8484 7476
rect 8428 7422 8430 7474
rect 8430 7422 8482 7474
rect 8482 7422 8484 7474
rect 8428 7420 8484 7422
rect 7868 6748 7924 6804
rect 8204 6076 8260 6132
rect 8652 6018 8708 6020
rect 8652 5966 8654 6018
rect 8654 5966 8706 6018
rect 8706 5966 8708 6018
rect 8652 5964 8708 5966
rect 7980 3612 8036 3668
rect 8092 4172 8148 4228
rect 7868 3442 7924 3444
rect 7868 3390 7870 3442
rect 7870 3390 7922 3442
rect 7922 3390 7924 3442
rect 7868 3388 7924 3390
rect 8316 4172 8372 4228
rect 8652 3612 8708 3668
rect 8988 8092 9044 8148
rect 9436 8034 9492 8036
rect 9436 7982 9438 8034
rect 9438 7982 9490 8034
rect 9490 7982 9492 8034
rect 9436 7980 9492 7982
rect 10220 9154 10276 9156
rect 10220 9102 10222 9154
rect 10222 9102 10274 9154
rect 10274 9102 10276 9154
rect 10220 9100 10276 9102
rect 9884 9042 9940 9044
rect 9884 8990 9886 9042
rect 9886 8990 9938 9042
rect 9938 8990 9940 9042
rect 9884 8988 9940 8990
rect 10556 9714 10612 9716
rect 10556 9662 10558 9714
rect 10558 9662 10610 9714
rect 10610 9662 10612 9714
rect 10556 9660 10612 9662
rect 10892 9602 10948 9604
rect 10892 9550 10894 9602
rect 10894 9550 10946 9602
rect 10946 9550 10948 9602
rect 10892 9548 10948 9550
rect 10444 5010 10500 5012
rect 10444 4958 10446 5010
rect 10446 4958 10498 5010
rect 10498 4958 10500 5010
rect 10444 4956 10500 4958
rect 9660 4338 9716 4340
rect 9660 4286 9662 4338
rect 9662 4286 9714 4338
rect 9714 4286 9716 4338
rect 9660 4284 9716 4286
rect 9548 3666 9604 3668
rect 9548 3614 9550 3666
rect 9550 3614 9602 3666
rect 9602 3614 9604 3666
rect 9548 3612 9604 3614
rect 9324 3388 9380 3444
rect 9996 3442 10052 3444
rect 9996 3390 9998 3442
rect 9998 3390 10050 3442
rect 10050 3390 10052 3442
rect 9996 3388 10052 3390
rect 11116 4956 11172 5012
rect 11228 5740 11284 5796
rect 11900 11170 11956 11172
rect 11900 11118 11902 11170
rect 11902 11118 11954 11170
rect 11954 11118 11956 11170
rect 11900 11116 11956 11118
rect 11900 5794 11956 5796
rect 11900 5742 11902 5794
rect 11902 5742 11954 5794
rect 11954 5742 11956 5794
rect 11900 5740 11956 5742
rect 11340 4956 11396 5012
rect 10892 3442 10948 3444
rect 10892 3390 10894 3442
rect 10894 3390 10946 3442
rect 10946 3390 10948 3442
rect 10892 3388 10948 3390
rect 12460 5010 12516 5012
rect 12460 4958 12462 5010
rect 12462 4958 12514 5010
rect 12514 4958 12516 5010
rect 12460 4956 12516 4958
rect 12460 4732 12516 4788
rect 13580 11394 13636 11396
rect 13580 11342 13582 11394
rect 13582 11342 13634 11394
rect 13634 11342 13636 11394
rect 13580 11340 13636 11342
rect 12796 11282 12852 11284
rect 12796 11230 12798 11282
rect 12798 11230 12850 11282
rect 12850 11230 12852 11282
rect 12796 11228 12852 11230
rect 12684 5740 12740 5796
rect 13468 4956 13524 5012
rect 11676 3442 11732 3444
rect 11676 3390 11678 3442
rect 11678 3390 11730 3442
rect 11730 3390 11732 3442
rect 11676 3388 11732 3390
rect 13916 5794 13972 5796
rect 13916 5742 13918 5794
rect 13918 5742 13970 5794
rect 13970 5742 13972 5794
rect 13916 5740 13972 5742
rect 13692 5010 13748 5012
rect 13692 4958 13694 5010
rect 13694 4958 13746 5010
rect 13746 4958 13748 5010
rect 13692 4956 13748 4958
rect 18844 17554 18900 17556
rect 18844 17502 18846 17554
rect 18846 17502 18898 17554
rect 18898 17502 18900 17554
rect 18844 17500 18900 17502
rect 18732 17052 18788 17108
rect 20188 18396 20244 18452
rect 20860 20018 20916 20020
rect 20860 19966 20862 20018
rect 20862 19966 20914 20018
rect 20914 19966 20916 20018
rect 20860 19964 20916 19966
rect 20860 19010 20916 19012
rect 20860 18958 20862 19010
rect 20862 18958 20914 19010
rect 20914 18958 20916 19010
rect 20860 18956 20916 18958
rect 20860 18620 20916 18676
rect 20524 18396 20580 18452
rect 20300 17666 20356 17668
rect 20300 17614 20302 17666
rect 20302 17614 20354 17666
rect 20354 17614 20356 17666
rect 20300 17612 20356 17614
rect 21196 20242 21252 20244
rect 21196 20190 21198 20242
rect 21198 20190 21250 20242
rect 21250 20190 21252 20242
rect 21196 20188 21252 20190
rect 23660 21586 23716 21588
rect 23660 21534 23662 21586
rect 23662 21534 23714 21586
rect 23714 21534 23716 21586
rect 23660 21532 23716 21534
rect 23212 20802 23268 20804
rect 23212 20750 23214 20802
rect 23214 20750 23266 20802
rect 23266 20750 23268 20802
rect 23212 20748 23268 20750
rect 23548 20578 23604 20580
rect 23548 20526 23550 20578
rect 23550 20526 23602 20578
rect 23602 20526 23604 20578
rect 23548 20524 23604 20526
rect 24892 24668 24948 24724
rect 26124 24834 26180 24836
rect 26124 24782 26126 24834
rect 26126 24782 26178 24834
rect 26178 24782 26180 24834
rect 26124 24780 26180 24782
rect 25676 23714 25732 23716
rect 25676 23662 25678 23714
rect 25678 23662 25730 23714
rect 25730 23662 25732 23714
rect 25676 23660 25732 23662
rect 24220 21756 24276 21812
rect 23996 21698 24052 21700
rect 23996 21646 23998 21698
rect 23998 21646 24050 21698
rect 24050 21646 24052 21698
rect 23996 21644 24052 21646
rect 23884 21532 23940 21588
rect 21644 20018 21700 20020
rect 21644 19966 21646 20018
rect 21646 19966 21698 20018
rect 21698 19966 21700 20018
rect 21644 19964 21700 19966
rect 21980 19122 22036 19124
rect 21980 19070 21982 19122
rect 21982 19070 22034 19122
rect 22034 19070 22036 19122
rect 21980 19068 22036 19070
rect 21532 18674 21588 18676
rect 21532 18622 21534 18674
rect 21534 18622 21586 18674
rect 21586 18622 21588 18674
rect 21532 18620 21588 18622
rect 21084 18396 21140 18452
rect 18508 16994 18564 16996
rect 18508 16942 18510 16994
rect 18510 16942 18562 16994
rect 18562 16942 18564 16994
rect 18508 16940 18564 16942
rect 18732 16828 18788 16884
rect 17052 15260 17108 15316
rect 17052 15036 17108 15092
rect 16940 14252 16996 14308
rect 16828 13692 16884 13748
rect 16044 5852 16100 5908
rect 15820 5010 15876 5012
rect 15820 4958 15822 5010
rect 15822 4958 15874 5010
rect 15874 4958 15876 5010
rect 15820 4956 15876 4958
rect 14476 4732 14532 4788
rect 13804 3442 13860 3444
rect 13804 3390 13806 3442
rect 13806 3390 13858 3442
rect 13858 3390 13860 3442
rect 13804 3388 13860 3390
rect 14700 3442 14756 3444
rect 14700 3390 14702 3442
rect 14702 3390 14754 3442
rect 14754 3390 14756 3442
rect 14700 3388 14756 3390
rect 15372 3388 15428 3444
rect 16716 5794 16772 5796
rect 16716 5742 16718 5794
rect 16718 5742 16770 5794
rect 16770 5742 16772 5794
rect 16716 5740 16772 5742
rect 16604 5628 16660 5684
rect 16716 5234 16772 5236
rect 16716 5182 16718 5234
rect 16718 5182 16770 5234
rect 16770 5182 16772 5234
rect 16716 5180 16772 5182
rect 17052 5740 17108 5796
rect 18284 15372 18340 15428
rect 18844 16098 18900 16100
rect 18844 16046 18846 16098
rect 18846 16046 18898 16098
rect 18898 16046 18900 16098
rect 18844 16044 18900 16046
rect 19292 17052 19348 17108
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20188 17276 20244 17332
rect 20044 17220 20100 17222
rect 20860 17388 20916 17444
rect 20860 17164 20916 17220
rect 19180 16882 19236 16884
rect 19180 16830 19182 16882
rect 19182 16830 19234 16882
rect 19234 16830 19236 16882
rect 19180 16828 19236 16830
rect 18508 15820 18564 15876
rect 18508 15260 18564 15316
rect 17724 15036 17780 15092
rect 20412 16882 20468 16884
rect 20412 16830 20414 16882
rect 20414 16830 20466 16882
rect 20466 16830 20468 16882
rect 20412 16828 20468 16830
rect 19516 16156 19572 16212
rect 20748 16716 20804 16772
rect 20188 15986 20244 15988
rect 20188 15934 20190 15986
rect 20190 15934 20242 15986
rect 20242 15934 20244 15986
rect 20188 15932 20244 15934
rect 19404 15820 19460 15876
rect 19740 15874 19796 15876
rect 19740 15822 19742 15874
rect 19742 15822 19794 15874
rect 19794 15822 19796 15874
rect 19740 15820 19796 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 17276 5628 17332 5684
rect 17948 5628 18004 5684
rect 17164 5180 17220 5236
rect 17388 4956 17444 5012
rect 17836 5010 17892 5012
rect 17836 4958 17838 5010
rect 17838 4958 17890 5010
rect 17890 4958 17892 5010
rect 17836 4956 17892 4958
rect 17612 3442 17668 3444
rect 17612 3390 17614 3442
rect 17614 3390 17666 3442
rect 17666 3390 17668 3442
rect 17612 3388 17668 3390
rect 18060 3388 18116 3444
rect 18396 5906 18452 5908
rect 18396 5854 18398 5906
rect 18398 5854 18450 5906
rect 18450 5854 18452 5906
rect 18396 5852 18452 5854
rect 19068 15260 19124 15316
rect 19628 15148 19684 15204
rect 19404 5964 19460 6020
rect 18732 4956 18788 5012
rect 19516 5180 19572 5236
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20300 6018 20356 6020
rect 20300 5966 20302 6018
rect 20302 5966 20354 6018
rect 20354 5966 20356 6018
rect 20300 5964 20356 5966
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19852 4450 19908 4452
rect 19852 4398 19854 4450
rect 19854 4398 19906 4450
rect 19906 4398 19908 4450
rect 19852 4396 19908 4398
rect 21084 17106 21140 17108
rect 21084 17054 21086 17106
rect 21086 17054 21138 17106
rect 21138 17054 21140 17106
rect 21084 17052 21140 17054
rect 21196 16716 21252 16772
rect 21532 17612 21588 17668
rect 21980 17164 22036 17220
rect 22428 17164 22484 17220
rect 22316 16770 22372 16772
rect 22316 16718 22318 16770
rect 22318 16718 22370 16770
rect 22370 16718 22372 16770
rect 22316 16716 22372 16718
rect 23100 17164 23156 17220
rect 22652 16098 22708 16100
rect 22652 16046 22654 16098
rect 22654 16046 22706 16098
rect 22706 16046 22708 16098
rect 22652 16044 22708 16046
rect 22652 15708 22708 15764
rect 20972 5068 21028 5124
rect 21980 5234 22036 5236
rect 21980 5182 21982 5234
rect 21982 5182 22034 5234
rect 22034 5182 22036 5234
rect 21980 5180 22036 5182
rect 21644 5122 21700 5124
rect 21644 5070 21646 5122
rect 21646 5070 21698 5122
rect 21698 5070 21700 5122
rect 21644 5068 21700 5070
rect 21308 4396 21364 4452
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21868 3500 21924 3556
rect 23324 17052 23380 17108
rect 23212 16770 23268 16772
rect 23212 16718 23214 16770
rect 23214 16718 23266 16770
rect 23266 16718 23268 16770
rect 23212 16716 23268 16718
rect 23660 16882 23716 16884
rect 23660 16830 23662 16882
rect 23662 16830 23714 16882
rect 23714 16830 23716 16882
rect 23660 16828 23716 16830
rect 23436 15708 23492 15764
rect 26684 25282 26740 25284
rect 26684 25230 26686 25282
rect 26686 25230 26738 25282
rect 26738 25230 26740 25282
rect 26684 25228 26740 25230
rect 24556 22764 24612 22820
rect 24444 21586 24500 21588
rect 24444 21534 24446 21586
rect 24446 21534 24498 21586
rect 24498 21534 24500 21586
rect 24444 21532 24500 21534
rect 22540 3554 22596 3556
rect 22540 3502 22542 3554
rect 22542 3502 22594 3554
rect 22594 3502 22596 3554
rect 22540 3500 22596 3502
rect 24444 17164 24500 17220
rect 24220 16828 24276 16884
rect 25228 17276 25284 17332
rect 24892 16882 24948 16884
rect 24892 16830 24894 16882
rect 24894 16830 24946 16882
rect 24946 16830 24948 16882
rect 24892 16828 24948 16830
rect 24332 15708 24388 15764
rect 24332 13356 24388 13412
rect 24108 4172 24164 4228
rect 23324 3500 23380 3556
rect 23436 3442 23492 3444
rect 23436 3390 23438 3442
rect 23438 3390 23490 3442
rect 23490 3390 23492 3442
rect 23436 3388 23492 3390
rect 26012 17388 26068 17444
rect 25676 17164 25732 17220
rect 26124 17276 26180 17332
rect 25900 16882 25956 16884
rect 25900 16830 25902 16882
rect 25902 16830 25954 16882
rect 25954 16830 25956 16882
rect 25900 16828 25956 16830
rect 26572 17276 26628 17332
rect 26684 16882 26740 16884
rect 26684 16830 26686 16882
rect 26686 16830 26738 16882
rect 26738 16830 26740 16882
rect 26684 16828 26740 16830
rect 25340 13356 25396 13412
rect 26572 6524 26628 6580
rect 24780 4284 24836 4340
rect 26012 4338 26068 4340
rect 26012 4286 26014 4338
rect 26014 4286 26066 4338
rect 26066 4286 26068 4338
rect 26012 4284 26068 4286
rect 25564 4226 25620 4228
rect 25564 4174 25566 4226
rect 25566 4174 25618 4226
rect 25618 4174 25620 4226
rect 25564 4172 25620 4174
rect 26124 4172 26180 4228
rect 25340 3442 25396 3444
rect 25340 3390 25342 3442
rect 25342 3390 25394 3442
rect 25394 3390 25396 3442
rect 25340 3388 25396 3390
rect 27356 26290 27412 26292
rect 27356 26238 27358 26290
rect 27358 26238 27410 26290
rect 27410 26238 27412 26290
rect 27356 26236 27412 26238
rect 27916 26962 27972 26964
rect 27916 26910 27918 26962
rect 27918 26910 27970 26962
rect 27970 26910 27972 26962
rect 27916 26908 27972 26910
rect 28252 26850 28308 26852
rect 28252 26798 28254 26850
rect 28254 26798 28306 26850
rect 28306 26798 28308 26850
rect 28252 26796 28308 26798
rect 27692 26402 27748 26404
rect 27692 26350 27694 26402
rect 27694 26350 27746 26402
rect 27746 26350 27748 26402
rect 27692 26348 27748 26350
rect 27580 26012 27636 26068
rect 27356 25900 27412 25956
rect 27468 25788 27524 25844
rect 27580 25506 27636 25508
rect 27580 25454 27582 25506
rect 27582 25454 27634 25506
rect 27634 25454 27636 25506
rect 27580 25452 27636 25454
rect 26796 4226 26852 4228
rect 26796 4174 26798 4226
rect 26798 4174 26850 4226
rect 26850 4174 26852 4226
rect 26796 4172 26852 4174
rect 30940 31106 30996 31108
rect 30940 31054 30942 31106
rect 30942 31054 30994 31106
rect 30994 31054 30996 31106
rect 30940 31052 30996 31054
rect 31612 31554 31668 31556
rect 31612 31502 31614 31554
rect 31614 31502 31666 31554
rect 31666 31502 31668 31554
rect 31612 31500 31668 31502
rect 31276 30994 31332 30996
rect 31276 30942 31278 30994
rect 31278 30942 31330 30994
rect 31330 30942 31332 30994
rect 31276 30940 31332 30942
rect 30492 30098 30548 30100
rect 30492 30046 30494 30098
rect 30494 30046 30546 30098
rect 30546 30046 30548 30098
rect 30492 30044 30548 30046
rect 30940 30044 30996 30100
rect 30044 29932 30100 29988
rect 30828 29986 30884 29988
rect 30828 29934 30830 29986
rect 30830 29934 30882 29986
rect 30882 29934 30884 29986
rect 30828 29932 30884 29934
rect 30380 29538 30436 29540
rect 30380 29486 30382 29538
rect 30382 29486 30434 29538
rect 30434 29486 30436 29538
rect 30380 29484 30436 29486
rect 28924 29260 28980 29316
rect 29260 29426 29316 29428
rect 29260 29374 29262 29426
rect 29262 29374 29314 29426
rect 29314 29374 29316 29426
rect 29260 29372 29316 29374
rect 28924 27970 28980 27972
rect 28924 27918 28926 27970
rect 28926 27918 28978 27970
rect 28978 27918 28980 27970
rect 28924 27916 28980 27918
rect 28812 26962 28868 26964
rect 28812 26910 28814 26962
rect 28814 26910 28866 26962
rect 28866 26910 28868 26962
rect 28812 26908 28868 26910
rect 30044 29426 30100 29428
rect 30044 29374 30046 29426
rect 30046 29374 30098 29426
rect 30098 29374 30100 29426
rect 30044 29372 30100 29374
rect 29372 28476 29428 28532
rect 29596 28530 29652 28532
rect 29596 28478 29598 28530
rect 29598 28478 29650 28530
rect 29650 28478 29652 28530
rect 29596 28476 29652 28478
rect 29932 28418 29988 28420
rect 29932 28366 29934 28418
rect 29934 28366 29986 28418
rect 29986 28366 29988 28418
rect 29932 28364 29988 28366
rect 29820 27858 29876 27860
rect 29820 27806 29822 27858
rect 29822 27806 29874 27858
rect 29874 27806 29876 27858
rect 29820 27804 29876 27806
rect 28028 6578 28084 6580
rect 28028 6526 28030 6578
rect 28030 6526 28082 6578
rect 28082 6526 28084 6578
rect 28028 6524 28084 6526
rect 27692 5964 27748 6020
rect 27468 3442 27524 3444
rect 27468 3390 27470 3442
rect 27470 3390 27522 3442
rect 27522 3390 27524 3442
rect 27468 3388 27524 3390
rect 28364 5010 28420 5012
rect 28364 4958 28366 5010
rect 28366 4958 28418 5010
rect 28418 4958 28420 5010
rect 28364 4956 28420 4958
rect 28700 6018 28756 6020
rect 28700 5966 28702 6018
rect 28702 5966 28754 6018
rect 28754 5966 28756 6018
rect 28700 5964 28756 5966
rect 29596 5964 29652 6020
rect 29484 5852 29540 5908
rect 30380 6018 30436 6020
rect 30380 5966 30382 6018
rect 30382 5966 30434 6018
rect 30434 5966 30436 6018
rect 30380 5964 30436 5966
rect 29932 5010 29988 5012
rect 29932 4958 29934 5010
rect 29934 4958 29986 5010
rect 29986 4958 29988 5010
rect 29932 4956 29988 4958
rect 29820 4450 29876 4452
rect 29820 4398 29822 4450
rect 29822 4398 29874 4450
rect 29874 4398 29876 4450
rect 29820 4396 29876 4398
rect 31052 5964 31108 6020
rect 31388 30098 31444 30100
rect 31388 30046 31390 30098
rect 31390 30046 31442 30098
rect 31442 30046 31444 30098
rect 31388 30044 31444 30046
rect 31724 30098 31780 30100
rect 31724 30046 31726 30098
rect 31726 30046 31778 30098
rect 31778 30046 31780 30098
rect 31724 30044 31780 30046
rect 32284 32284 32340 32340
rect 31948 31778 32004 31780
rect 31948 31726 31950 31778
rect 31950 31726 32002 31778
rect 32002 31726 32004 31778
rect 31948 31724 32004 31726
rect 32284 31106 32340 31108
rect 32284 31054 32286 31106
rect 32286 31054 32338 31106
rect 32338 31054 32340 31106
rect 32284 31052 32340 31054
rect 32060 30994 32116 30996
rect 32060 30942 32062 30994
rect 32062 30942 32114 30994
rect 32114 30942 32116 30994
rect 32060 30940 32116 30942
rect 31500 29314 31556 29316
rect 31500 29262 31502 29314
rect 31502 29262 31554 29314
rect 31554 29262 31556 29314
rect 31500 29260 31556 29262
rect 30828 4396 30884 4452
rect 29708 3442 29764 3444
rect 29708 3390 29710 3442
rect 29710 3390 29762 3442
rect 29762 3390 29764 3442
rect 29708 3388 29764 3390
rect 34412 33122 34468 33124
rect 34412 33070 34414 33122
rect 34414 33070 34466 33122
rect 34466 33070 34468 33122
rect 34412 33068 34468 33070
rect 33964 32674 34020 32676
rect 33964 32622 33966 32674
rect 33966 32622 34018 32674
rect 34018 32622 34020 32674
rect 33964 32620 34020 32622
rect 32508 32562 32564 32564
rect 32508 32510 32510 32562
rect 32510 32510 32562 32562
rect 32562 32510 32564 32562
rect 32508 32508 32564 32510
rect 33628 32562 33684 32564
rect 33628 32510 33630 32562
rect 33630 32510 33682 32562
rect 33682 32510 33684 32562
rect 33628 32508 33684 32510
rect 32844 31778 32900 31780
rect 32844 31726 32846 31778
rect 32846 31726 32898 31778
rect 32898 31726 32900 31778
rect 32844 31724 32900 31726
rect 33964 31778 34020 31780
rect 33964 31726 33966 31778
rect 33966 31726 34018 31778
rect 34018 31726 34020 31778
rect 33964 31724 34020 31726
rect 33068 31554 33124 31556
rect 33068 31502 33070 31554
rect 33070 31502 33122 31554
rect 33122 31502 33124 31554
rect 33068 31500 33124 31502
rect 32732 30994 32788 30996
rect 32732 30942 32734 30994
rect 32734 30942 32786 30994
rect 32786 30942 32788 30994
rect 32732 30940 32788 30942
rect 31612 5404 31668 5460
rect 31388 3442 31444 3444
rect 31388 3390 31390 3442
rect 31390 3390 31442 3442
rect 31442 3390 31444 3442
rect 31388 3388 31444 3390
rect 32396 5404 32452 5460
rect 33516 5404 33572 5460
rect 34860 5964 34916 6020
rect 32284 4284 32340 4340
rect 33516 4338 33572 4340
rect 33516 4286 33518 4338
rect 33518 4286 33570 4338
rect 33570 4286 33572 4338
rect 33516 4284 33572 4286
rect 32844 4172 32900 4228
rect 33964 4226 34020 4228
rect 33964 4174 33966 4226
rect 33966 4174 34018 4226
rect 34018 4174 34020 4226
rect 33964 4172 34020 4174
rect 33180 3442 33236 3444
rect 33180 3390 33182 3442
rect 33182 3390 33234 3442
rect 33234 3390 33236 3442
rect 33180 3388 33236 3390
rect 34412 3442 34468 3444
rect 34412 3390 34414 3442
rect 34414 3390 34466 3442
rect 34466 3390 34468 3442
rect 34412 3388 34468 3390
rect 35980 35698 36036 35700
rect 35980 35646 35982 35698
rect 35982 35646 36034 35698
rect 36034 35646 36036 35698
rect 35980 35644 36036 35646
rect 36988 35810 37044 35812
rect 36988 35758 36990 35810
rect 36990 35758 37042 35810
rect 37042 35758 37044 35810
rect 36988 35756 37044 35758
rect 36540 35532 36596 35588
rect 35420 35420 35476 35476
rect 36092 35420 36148 35476
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35308 34748 35364 34804
rect 35084 34242 35140 34244
rect 35084 34190 35086 34242
rect 35086 34190 35138 34242
rect 35138 34190 35140 34242
rect 35084 34188 35140 34190
rect 36428 34802 36484 34804
rect 36428 34750 36430 34802
rect 36430 34750 36482 34802
rect 36482 34750 36484 34802
rect 36428 34748 36484 34750
rect 35532 34690 35588 34692
rect 35532 34638 35534 34690
rect 35534 34638 35586 34690
rect 35586 34638 35588 34690
rect 35532 34636 35588 34638
rect 36204 34130 36260 34132
rect 36204 34078 36206 34130
rect 36206 34078 36258 34130
rect 36258 34078 36260 34130
rect 36204 34076 36260 34078
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 6018 35252 6020
rect 35196 5966 35198 6018
rect 35198 5966 35250 6018
rect 35250 5966 35252 6018
rect 35196 5964 35252 5966
rect 36652 35698 36708 35700
rect 36652 35646 36654 35698
rect 36654 35646 36706 35698
rect 36706 35646 36708 35698
rect 36652 35644 36708 35646
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35644 5068 35700 5124
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35532 3500 35588 3556
rect 35196 3442 35252 3444
rect 35196 3390 35198 3442
rect 35198 3390 35250 3442
rect 35250 3390 35252 3442
rect 35196 3388 35252 3390
rect 36316 5068 36372 5124
rect 38108 37266 38164 37268
rect 38108 37214 38110 37266
rect 38110 37214 38162 37266
rect 38162 37214 38164 37266
rect 38108 37212 38164 37214
rect 39116 37826 39172 37828
rect 39116 37774 39118 37826
rect 39118 37774 39170 37826
rect 39170 37774 39172 37826
rect 39116 37772 39172 37774
rect 37884 36258 37940 36260
rect 37884 36206 37886 36258
rect 37886 36206 37938 36258
rect 37938 36206 37940 36258
rect 37884 36204 37940 36206
rect 37884 35698 37940 35700
rect 37884 35646 37886 35698
rect 37886 35646 37938 35698
rect 37938 35646 37940 35698
rect 37884 35644 37940 35646
rect 38332 35698 38388 35700
rect 38332 35646 38334 35698
rect 38334 35646 38386 35698
rect 38386 35646 38388 35698
rect 38332 35644 38388 35646
rect 37436 35586 37492 35588
rect 37436 35534 37438 35586
rect 37438 35534 37490 35586
rect 37490 35534 37492 35586
rect 37436 35532 37492 35534
rect 37436 35308 37492 35364
rect 37436 5122 37492 5124
rect 37436 5070 37438 5122
rect 37438 5070 37490 5122
rect 37490 5070 37492 5122
rect 37436 5068 37492 5070
rect 38108 5740 38164 5796
rect 37996 4732 38052 4788
rect 38780 5794 38836 5796
rect 38780 5742 38782 5794
rect 38782 5742 38834 5794
rect 38834 5742 38836 5794
rect 38780 5740 38836 5742
rect 38892 5180 38948 5236
rect 37884 3666 37940 3668
rect 37884 3614 37886 3666
rect 37886 3614 37938 3666
rect 37938 3614 37940 3666
rect 37884 3612 37940 3614
rect 36204 3500 36260 3556
rect 36988 3554 37044 3556
rect 36988 3502 36990 3554
rect 36990 3502 37042 3554
rect 37042 3502 37044 3554
rect 36988 3500 37044 3502
rect 36876 3388 36932 3444
rect 38220 4732 38276 4788
rect 38668 4732 38724 4788
rect 38892 3612 38948 3668
rect 38332 3442 38388 3444
rect 38332 3390 38334 3442
rect 38334 3390 38386 3442
rect 38386 3390 38388 3442
rect 38332 3388 38388 3390
rect 39788 39506 39844 39508
rect 39788 39454 39790 39506
rect 39790 39454 39842 39506
rect 39842 39454 39844 39506
rect 39788 39452 39844 39454
rect 40124 39394 40180 39396
rect 40124 39342 40126 39394
rect 40126 39342 40178 39394
rect 40178 39342 40180 39394
rect 40124 39340 40180 39342
rect 39676 38946 39732 38948
rect 39676 38894 39678 38946
rect 39678 38894 39730 38946
rect 39730 38894 39732 38946
rect 39676 38892 39732 38894
rect 39452 38834 39508 38836
rect 39452 38782 39454 38834
rect 39454 38782 39506 38834
rect 39506 38782 39508 38834
rect 39452 38780 39508 38782
rect 41020 39564 41076 39620
rect 40012 37938 40068 37940
rect 40012 37886 40014 37938
rect 40014 37886 40066 37938
rect 40066 37886 40068 37938
rect 40012 37884 40068 37886
rect 39340 37266 39396 37268
rect 39340 37214 39342 37266
rect 39342 37214 39394 37266
rect 39394 37214 39396 37266
rect 39340 37212 39396 37214
rect 39676 5234 39732 5236
rect 39676 5182 39678 5234
rect 39678 5182 39730 5234
rect 39730 5182 39732 5234
rect 39676 5180 39732 5182
rect 40236 4732 40292 4788
rect 40124 3612 40180 3668
rect 39564 3388 39620 3444
rect 41580 4956 41636 5012
rect 41468 4732 41524 4788
rect 42476 40962 42532 40964
rect 42476 40910 42478 40962
rect 42478 40910 42530 40962
rect 42530 40910 42532 40962
rect 42476 40908 42532 40910
rect 42140 40572 42196 40628
rect 42364 40626 42420 40628
rect 42364 40574 42366 40626
rect 42366 40574 42418 40626
rect 42418 40574 42420 40626
rect 42364 40572 42420 40574
rect 41916 40514 41972 40516
rect 41916 40462 41918 40514
rect 41918 40462 41970 40514
rect 41970 40462 41972 40514
rect 41916 40460 41972 40462
rect 42812 40402 42868 40404
rect 42812 40350 42814 40402
rect 42814 40350 42866 40402
rect 42866 40350 42868 40402
rect 42812 40348 42868 40350
rect 44268 42642 44324 42644
rect 44268 42590 44270 42642
rect 44270 42590 44322 42642
rect 44322 42590 44324 42642
rect 44268 42588 44324 42590
rect 43708 42530 43764 42532
rect 43708 42478 43710 42530
rect 43710 42478 43762 42530
rect 43762 42478 43764 42530
rect 43708 42476 43764 42478
rect 43596 41858 43652 41860
rect 43596 41806 43598 41858
rect 43598 41806 43650 41858
rect 43650 41806 43652 41858
rect 43596 41804 43652 41806
rect 42924 5180 42980 5236
rect 41580 3388 41636 3444
rect 42812 4956 42868 5012
rect 43708 5234 43764 5236
rect 43708 5182 43710 5234
rect 43710 5182 43762 5234
rect 43762 5182 43764 5234
rect 43708 5180 43764 5182
rect 44828 4956 44884 5012
rect 43596 3612 43652 3668
rect 42924 3500 42980 3556
rect 42812 3442 42868 3444
rect 42812 3390 42814 3442
rect 42814 3390 42866 3442
rect 42866 3390 42868 3442
rect 42812 3388 42868 3390
rect 44268 3500 44324 3556
rect 44380 4172 44436 4228
rect 43708 3442 43764 3444
rect 43708 3390 43710 3442
rect 43710 3390 43762 3442
rect 43762 3390 43764 3442
rect 43708 3388 43764 3390
rect 46732 5964 46788 6020
rect 45612 5010 45668 5012
rect 45612 4958 45614 5010
rect 45614 4958 45666 5010
rect 45666 4958 45668 5010
rect 45612 4956 45668 4958
rect 45388 4172 45444 4228
rect 45724 4172 45780 4228
rect 46284 4172 46340 4228
rect 45948 3612 46004 3668
rect 45612 3388 45668 3444
rect 47292 6018 47348 6020
rect 47292 5966 47294 6018
rect 47294 5966 47346 6018
rect 47346 5966 47348 6018
rect 47292 5964 47348 5966
rect 47740 5180 47796 5236
rect 47852 45052 47908 45108
rect 47516 4226 47572 4228
rect 47516 4174 47518 4226
rect 47518 4174 47570 4226
rect 47570 4174 47572 4226
rect 47516 4172 47572 4174
rect 47628 4060 47684 4116
rect 46844 3666 46900 3668
rect 46844 3614 46846 3666
rect 46846 3614 46898 3666
rect 46898 3614 46900 3666
rect 46844 3612 46900 3614
rect 48972 5740 49028 5796
rect 48748 5234 48804 5236
rect 48748 5182 48750 5234
rect 48750 5182 48802 5234
rect 48802 5182 48804 5234
rect 48748 5180 48804 5182
rect 47852 3612 47908 3668
rect 48300 5068 48356 5124
rect 48188 3442 48244 3444
rect 48188 3390 48190 3442
rect 48190 3390 48242 3442
rect 48242 3390 48244 3442
rect 48188 3388 48244 3390
rect 48748 4060 48804 4116
rect 48860 3666 48916 3668
rect 48860 3614 48862 3666
rect 48862 3614 48914 3666
rect 48914 3614 48916 3666
rect 48860 3612 48916 3614
rect 49644 5794 49700 5796
rect 49644 5742 49646 5794
rect 49646 5742 49698 5794
rect 49698 5742 49700 5794
rect 49644 5740 49700 5742
rect 49644 5122 49700 5124
rect 49644 5070 49646 5122
rect 49646 5070 49698 5122
rect 49698 5070 49700 5122
rect 49644 5068 49700 5070
rect 50652 49810 50708 49812
rect 50652 49758 50654 49810
rect 50654 49758 50706 49810
rect 50706 49758 50708 49810
rect 50652 49756 50708 49758
rect 51772 50594 51828 50596
rect 51772 50542 51774 50594
rect 51774 50542 51826 50594
rect 51826 50542 51828 50594
rect 51772 50540 51828 50542
rect 52332 50594 52388 50596
rect 52332 50542 52334 50594
rect 52334 50542 52386 50594
rect 52386 50542 52388 50594
rect 52332 50540 52388 50542
rect 50988 49756 51044 49812
rect 50652 49196 50708 49252
rect 51548 49698 51604 49700
rect 51548 49646 51550 49698
rect 51550 49646 51602 49698
rect 51602 49646 51604 49698
rect 51548 49644 51604 49646
rect 51212 49196 51268 49252
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50204 47346 50260 47348
rect 50204 47294 50206 47346
rect 50206 47294 50258 47346
rect 50258 47294 50260 47346
rect 50204 47292 50260 47294
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 49980 5852 50036 5908
rect 49868 4284 49924 4340
rect 49644 4172 49700 4228
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 50540 5906 50596 5908
rect 50540 5854 50542 5906
rect 50542 5854 50594 5906
rect 50594 5854 50596 5906
rect 50540 5852 50596 5854
rect 51212 5906 51268 5908
rect 51212 5854 51214 5906
rect 51214 5854 51266 5906
rect 51266 5854 51268 5906
rect 51212 5852 51268 5854
rect 50764 5292 50820 5348
rect 50988 5180 51044 5236
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 50540 4060 50596 4116
rect 50204 3724 50260 3780
rect 50316 3612 50372 3668
rect 49868 3442 49924 3444
rect 49868 3390 49870 3442
rect 49870 3390 49922 3442
rect 49922 3390 49924 3442
rect 49868 3388 49924 3390
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 51996 49698 52052 49700
rect 51996 49646 51998 49698
rect 51998 49646 52050 49698
rect 52050 49646 52052 49698
rect 51996 49644 52052 49646
rect 52780 51884 52836 51940
rect 52444 6524 52500 6580
rect 53116 52946 53172 52948
rect 53116 52894 53118 52946
rect 53118 52894 53170 52946
rect 53170 52894 53172 52946
rect 53116 52892 53172 52894
rect 52892 51548 52948 51604
rect 53340 52834 53396 52836
rect 53340 52782 53342 52834
rect 53342 52782 53394 52834
rect 53394 52782 53396 52834
rect 53340 52780 53396 52782
rect 53676 52780 53732 52836
rect 53676 51938 53732 51940
rect 53676 51886 53678 51938
rect 53678 51886 53730 51938
rect 53730 51886 53732 51938
rect 53676 51884 53732 51886
rect 53340 51602 53396 51604
rect 53340 51550 53342 51602
rect 53342 51550 53394 51602
rect 53394 51550 53396 51602
rect 53340 51548 53396 51550
rect 53676 51548 53732 51604
rect 53788 51436 53844 51492
rect 53452 50370 53508 50372
rect 53452 50318 53454 50370
rect 53454 50318 53506 50370
rect 53506 50318 53508 50370
rect 53452 50316 53508 50318
rect 53676 17052 53732 17108
rect 53676 14306 53732 14308
rect 53676 14254 53678 14306
rect 53678 14254 53730 14306
rect 53730 14254 53732 14306
rect 53676 14252 53732 14254
rect 53004 6412 53060 6468
rect 52780 6300 52836 6356
rect 51996 6188 52052 6244
rect 53004 6188 53060 6244
rect 53340 6188 53396 6244
rect 51660 5292 51716 5348
rect 51996 5234 52052 5236
rect 51996 5182 51998 5234
rect 51998 5182 52050 5234
rect 52050 5182 52052 5234
rect 51996 5180 52052 5182
rect 53004 4956 53060 5012
rect 51548 4338 51604 4340
rect 51548 4286 51550 4338
rect 51550 4286 51602 4338
rect 51602 4286 51604 4338
rect 51548 4284 51604 4286
rect 52220 4226 52276 4228
rect 52220 4174 52222 4226
rect 52222 4174 52274 4226
rect 52274 4174 52276 4226
rect 52220 4172 52276 4174
rect 52108 3724 52164 3780
rect 52780 3724 52836 3780
rect 51660 3500 51716 3556
rect 52332 3388 52388 3444
rect 54908 53506 54964 53508
rect 54908 53454 54910 53506
rect 54910 53454 54962 53506
rect 54962 53454 54964 53506
rect 54908 53452 54964 53454
rect 54124 52834 54180 52836
rect 54124 52782 54126 52834
rect 54126 52782 54178 52834
rect 54178 52782 54180 52834
rect 54124 52780 54180 52782
rect 54012 52668 54068 52724
rect 54236 52386 54292 52388
rect 54236 52334 54238 52386
rect 54238 52334 54290 52386
rect 54290 52334 54292 52386
rect 54236 52332 54292 52334
rect 55692 55410 55748 55412
rect 55692 55358 55694 55410
rect 55694 55358 55746 55410
rect 55746 55358 55748 55410
rect 55692 55356 55748 55358
rect 55244 54348 55300 54404
rect 54124 17666 54180 17668
rect 54124 17614 54126 17666
rect 54126 17614 54178 17666
rect 54178 17614 54180 17666
rect 54124 17612 54180 17614
rect 54124 15148 54180 15204
rect 53900 5964 53956 6020
rect 54236 6524 54292 6580
rect 54908 18508 54964 18564
rect 55132 18284 55188 18340
rect 54572 16882 54628 16884
rect 54572 16830 54574 16882
rect 54574 16830 54626 16882
rect 54626 16830 54628 16882
rect 54572 16828 54628 16830
rect 54572 13746 54628 13748
rect 54572 13694 54574 13746
rect 54574 13694 54626 13746
rect 54626 13694 54628 13746
rect 54572 13692 54628 13694
rect 55132 17052 55188 17108
rect 55132 14252 55188 14308
rect 55020 13692 55076 13748
rect 54348 6188 54404 6244
rect 54460 6300 54516 6356
rect 53564 5010 53620 5012
rect 53564 4958 53566 5010
rect 53566 4958 53618 5010
rect 53618 4958 53620 5010
rect 53564 4956 53620 4958
rect 55356 54290 55412 54292
rect 55356 54238 55358 54290
rect 55358 54238 55410 54290
rect 55410 54238 55412 54290
rect 55356 54236 55412 54238
rect 55580 53506 55636 53508
rect 55580 53454 55582 53506
rect 55582 53454 55634 53506
rect 55634 53454 55636 53506
rect 55580 53452 55636 53454
rect 58044 60002 58100 60004
rect 58044 59950 58046 60002
rect 58046 59950 58098 60002
rect 58098 59950 58100 60002
rect 58044 59948 58100 59950
rect 58156 59890 58212 59892
rect 58156 59838 58158 59890
rect 58158 59838 58210 59890
rect 58210 59838 58212 59890
rect 58156 59836 58212 59838
rect 59612 59500 59668 59556
rect 60172 59890 60228 59892
rect 60172 59838 60174 59890
rect 60174 59838 60226 59890
rect 60226 59838 60228 59890
rect 60172 59836 60228 59838
rect 59948 59500 60004 59556
rect 60284 59724 60340 59780
rect 58380 59218 58436 59220
rect 58380 59166 58382 59218
rect 58382 59166 58434 59218
rect 58434 59166 58436 59218
rect 58380 59164 58436 59166
rect 58940 59218 58996 59220
rect 58940 59166 58942 59218
rect 58942 59166 58994 59218
rect 58994 59166 58996 59218
rect 58940 59164 58996 59166
rect 57372 59052 57428 59108
rect 57260 58434 57316 58436
rect 57260 58382 57262 58434
rect 57262 58382 57314 58434
rect 57314 58382 57316 58434
rect 57260 58380 57316 58382
rect 56700 58210 56756 58212
rect 56700 58158 56702 58210
rect 56702 58158 56754 58210
rect 56754 58158 56756 58210
rect 56700 58156 56756 58158
rect 58156 58434 58212 58436
rect 58156 58382 58158 58434
rect 58158 58382 58210 58434
rect 58210 58382 58212 58434
rect 58156 58380 58212 58382
rect 57148 58156 57204 58212
rect 56140 57650 56196 57652
rect 56140 57598 56142 57650
rect 56142 57598 56194 57650
rect 56194 57598 56196 57650
rect 56140 57596 56196 57598
rect 56028 57538 56084 57540
rect 56028 57486 56030 57538
rect 56030 57486 56082 57538
rect 56082 57486 56084 57538
rect 56028 57484 56084 57486
rect 56588 57538 56644 57540
rect 56588 57486 56590 57538
rect 56590 57486 56642 57538
rect 56642 57486 56644 57538
rect 56588 57484 56644 57486
rect 55916 57036 55972 57092
rect 56140 56754 56196 56756
rect 56140 56702 56142 56754
rect 56142 56702 56194 56754
rect 56194 56702 56196 56754
rect 56140 56700 56196 56702
rect 56588 56754 56644 56756
rect 56588 56702 56590 56754
rect 56590 56702 56642 56754
rect 56642 56702 56644 56754
rect 56588 56700 56644 56702
rect 56700 56252 56756 56308
rect 56700 56082 56756 56084
rect 56700 56030 56702 56082
rect 56702 56030 56754 56082
rect 56754 56030 56756 56082
rect 56700 56028 56756 56030
rect 57596 56866 57652 56868
rect 57596 56814 57598 56866
rect 57598 56814 57650 56866
rect 57650 56814 57652 56866
rect 57596 56812 57652 56814
rect 55916 55298 55972 55300
rect 55916 55246 55918 55298
rect 55918 55246 55970 55298
rect 55970 55246 55972 55298
rect 55916 55244 55972 55246
rect 56588 55244 56644 55300
rect 56364 55132 56420 55188
rect 55916 54290 55972 54292
rect 55916 54238 55918 54290
rect 55918 54238 55970 54290
rect 55970 54238 55972 54290
rect 55916 54236 55972 54238
rect 55468 49532 55524 49588
rect 55692 51324 55748 51380
rect 55580 18562 55636 18564
rect 55580 18510 55582 18562
rect 55582 18510 55634 18562
rect 55634 18510 55636 18562
rect 55580 18508 55636 18510
rect 56924 55186 56980 55188
rect 56924 55134 56926 55186
rect 56926 55134 56978 55186
rect 56978 55134 56980 55186
rect 56924 55132 56980 55134
rect 56700 54626 56756 54628
rect 56700 54574 56702 54626
rect 56702 54574 56754 54626
rect 56754 54574 56756 54626
rect 56700 54572 56756 54574
rect 56252 51548 56308 51604
rect 56588 51490 56644 51492
rect 56588 51438 56590 51490
rect 56590 51438 56642 51490
rect 56642 51438 56644 51490
rect 56588 51436 56644 51438
rect 56252 51378 56308 51380
rect 56252 51326 56254 51378
rect 56254 51326 56306 51378
rect 56306 51326 56308 51378
rect 56252 51324 56308 51326
rect 58044 57650 58100 57652
rect 58044 57598 58046 57650
rect 58046 57598 58098 57650
rect 58098 57598 58100 57650
rect 58044 57596 58100 57598
rect 57820 56978 57876 56980
rect 57820 56926 57822 56978
rect 57822 56926 57874 56978
rect 57874 56926 57876 56978
rect 57820 56924 57876 56926
rect 57820 56306 57876 56308
rect 57820 56254 57822 56306
rect 57822 56254 57874 56306
rect 57874 56254 57876 56306
rect 57820 56252 57876 56254
rect 57820 56028 57876 56084
rect 57708 55970 57764 55972
rect 57708 55918 57710 55970
rect 57710 55918 57762 55970
rect 57762 55918 57764 55970
rect 57708 55916 57764 55918
rect 57260 55186 57316 55188
rect 57260 55134 57262 55186
rect 57262 55134 57314 55186
rect 57314 55134 57316 55186
rect 57260 55132 57316 55134
rect 57372 54626 57428 54628
rect 57372 54574 57374 54626
rect 57374 54574 57426 54626
rect 57426 54574 57428 54626
rect 57372 54572 57428 54574
rect 57596 53900 57652 53956
rect 57484 52556 57540 52612
rect 57036 51548 57092 51604
rect 56924 51324 56980 51380
rect 56924 49532 56980 49588
rect 55804 18284 55860 18340
rect 55580 17666 55636 17668
rect 55580 17614 55582 17666
rect 55582 17614 55634 17666
rect 55634 17614 55636 17666
rect 55580 17612 55636 17614
rect 55356 17442 55412 17444
rect 55356 17390 55358 17442
rect 55358 17390 55410 17442
rect 55410 17390 55412 17442
rect 55356 17388 55412 17390
rect 56140 17666 56196 17668
rect 56140 17614 56142 17666
rect 56142 17614 56194 17666
rect 56194 17614 56196 17666
rect 56140 17612 56196 17614
rect 56700 17612 56756 17668
rect 56028 17388 56084 17444
rect 55356 16828 55412 16884
rect 56364 15426 56420 15428
rect 56364 15374 56366 15426
rect 56366 15374 56418 15426
rect 56418 15374 56420 15426
rect 56364 15372 56420 15374
rect 56028 15314 56084 15316
rect 56028 15262 56030 15314
rect 56030 15262 56082 15314
rect 56082 15262 56084 15314
rect 56028 15260 56084 15262
rect 55356 15148 55412 15204
rect 56140 14530 56196 14532
rect 56140 14478 56142 14530
rect 56142 14478 56194 14530
rect 56194 14478 56196 14530
rect 56140 14476 56196 14478
rect 56364 14306 56420 14308
rect 56364 14254 56366 14306
rect 56366 14254 56418 14306
rect 56418 14254 56420 14306
rect 56364 14252 56420 14254
rect 55692 13858 55748 13860
rect 55692 13806 55694 13858
rect 55694 13806 55746 13858
rect 55746 13806 55748 13858
rect 55692 13804 55748 13806
rect 55356 13746 55412 13748
rect 55356 13694 55358 13746
rect 55358 13694 55410 13746
rect 55410 13694 55412 13746
rect 55356 13692 55412 13694
rect 56812 14530 56868 14532
rect 56812 14478 56814 14530
rect 56814 14478 56866 14530
rect 56866 14478 56868 14530
rect 56812 14476 56868 14478
rect 56700 13468 56756 13524
rect 55804 6412 55860 6468
rect 55020 5180 55076 5236
rect 53676 4172 53732 4228
rect 53564 3666 53620 3668
rect 53564 3614 53566 3666
rect 53566 3614 53618 3666
rect 53618 3614 53620 3666
rect 53564 3612 53620 3614
rect 54012 3500 54068 3556
rect 54348 3612 54404 3668
rect 55356 6300 55412 6356
rect 57484 13468 57540 13524
rect 56924 6188 56980 6244
rect 57372 6300 57428 6356
rect 57820 13692 57876 13748
rect 58044 57372 58100 57428
rect 58044 56812 58100 56868
rect 58044 55132 58100 55188
rect 58044 53900 58100 53956
rect 58492 57650 58548 57652
rect 58492 57598 58494 57650
rect 58494 57598 58546 57650
rect 58546 57598 58548 57650
rect 58492 57596 58548 57598
rect 59276 58156 59332 58212
rect 59164 57596 59220 57652
rect 58268 56924 58324 56980
rect 58940 56754 58996 56756
rect 58940 56702 58942 56754
rect 58942 56702 58994 56754
rect 58994 56702 58996 56754
rect 58940 56700 58996 56702
rect 59500 56754 59556 56756
rect 59500 56702 59502 56754
rect 59502 56702 59554 56754
rect 59554 56702 59556 56754
rect 59500 56700 59556 56702
rect 58268 56082 58324 56084
rect 58268 56030 58270 56082
rect 58270 56030 58322 56082
rect 58322 56030 58324 56082
rect 58268 56028 58324 56030
rect 58828 56028 58884 56084
rect 57932 6636 57988 6692
rect 58604 55916 58660 55972
rect 58044 6412 58100 6468
rect 57708 6300 57764 6356
rect 58156 6188 58212 6244
rect 59276 52274 59332 52276
rect 59276 52222 59278 52274
rect 59278 52222 59330 52274
rect 59330 52222 59332 52274
rect 59276 52220 59332 52222
rect 59388 52162 59444 52164
rect 59388 52110 59390 52162
rect 59390 52110 59442 52162
rect 59442 52110 59444 52162
rect 59388 52108 59444 52110
rect 59164 6412 59220 6468
rect 56364 5964 56420 6020
rect 55916 5234 55972 5236
rect 55916 5182 55918 5234
rect 55918 5182 55970 5234
rect 55970 5182 55972 5234
rect 55916 5180 55972 5182
rect 55468 4226 55524 4228
rect 55468 4174 55470 4226
rect 55470 4174 55522 4226
rect 55522 4174 55524 4226
rect 55468 4172 55524 4174
rect 55804 3500 55860 3556
rect 55692 3442 55748 3444
rect 55692 3390 55694 3442
rect 55694 3390 55746 3442
rect 55746 3390 55748 3442
rect 55692 3388 55748 3390
rect 56364 3388 56420 3444
rect 59612 6300 59668 6356
rect 59836 58210 59892 58212
rect 59836 58158 59838 58210
rect 59838 58158 59890 58210
rect 59890 58158 59892 58210
rect 59836 58156 59892 58158
rect 60620 60002 60676 60004
rect 60620 59950 60622 60002
rect 60622 59950 60674 60002
rect 60674 59950 60676 60002
rect 60620 59948 60676 59950
rect 62188 61346 62244 61348
rect 62188 61294 62190 61346
rect 62190 61294 62242 61346
rect 62242 61294 62244 61346
rect 62188 61292 62244 61294
rect 62412 61010 62468 61012
rect 62412 60958 62414 61010
rect 62414 60958 62466 61010
rect 62466 60958 62468 61010
rect 62412 60956 62468 60958
rect 62636 60898 62692 60900
rect 62636 60846 62638 60898
rect 62638 60846 62690 60898
rect 62690 60846 62692 60898
rect 62636 60844 62692 60846
rect 61180 60674 61236 60676
rect 61180 60622 61182 60674
rect 61182 60622 61234 60674
rect 61234 60622 61236 60674
rect 61180 60620 61236 60622
rect 62188 60674 62244 60676
rect 62188 60622 62190 60674
rect 62190 60622 62242 60674
rect 62242 60622 62244 60674
rect 62188 60620 62244 60622
rect 62524 60674 62580 60676
rect 62524 60622 62526 60674
rect 62526 60622 62578 60674
rect 62578 60622 62580 60674
rect 62524 60620 62580 60622
rect 61404 60562 61460 60564
rect 61404 60510 61406 60562
rect 61406 60510 61458 60562
rect 61458 60510 61460 60562
rect 61404 60508 61460 60510
rect 61068 60060 61124 60116
rect 62748 60396 62804 60452
rect 61516 59890 61572 59892
rect 61516 59838 61518 59890
rect 61518 59838 61570 59890
rect 61570 59838 61572 59890
rect 61516 59836 61572 59838
rect 62076 59890 62132 59892
rect 62076 59838 62078 59890
rect 62078 59838 62130 59890
rect 62130 59838 62132 59890
rect 62076 59836 62132 59838
rect 61404 59778 61460 59780
rect 61404 59726 61406 59778
rect 61406 59726 61458 59778
rect 61458 59726 61460 59778
rect 61404 59724 61460 59726
rect 61292 59052 61348 59108
rect 61852 59106 61908 59108
rect 61852 59054 61854 59106
rect 61854 59054 61906 59106
rect 61906 59054 61908 59106
rect 61852 59052 61908 59054
rect 62748 59052 62804 59108
rect 63420 62914 63476 62916
rect 63420 62862 63422 62914
rect 63422 62862 63474 62914
rect 63474 62862 63476 62914
rect 63420 62860 63476 62862
rect 63532 61740 63588 61796
rect 63644 62860 63700 62916
rect 63196 60620 63252 60676
rect 62860 57762 62916 57764
rect 62860 57710 62862 57762
rect 62862 57710 62914 57762
rect 62914 57710 62916 57762
rect 62860 57708 62916 57710
rect 62748 57426 62804 57428
rect 62748 57374 62750 57426
rect 62750 57374 62802 57426
rect 62802 57374 62804 57426
rect 62748 57372 62804 57374
rect 59948 52162 60004 52164
rect 59948 52110 59950 52162
rect 59950 52110 60002 52162
rect 60002 52110 60004 52162
rect 59948 52108 60004 52110
rect 61404 53788 61460 53844
rect 60508 52444 60564 52500
rect 60060 6300 60116 6356
rect 60284 6636 60340 6692
rect 59724 6188 59780 6244
rect 57708 4172 57764 4228
rect 57372 3666 57428 3668
rect 57372 3614 57374 3666
rect 57374 3614 57426 3666
rect 57426 3614 57428 3666
rect 57372 3612 57428 3614
rect 58156 3500 58212 3556
rect 58380 3500 58436 3556
rect 61068 6188 61124 6244
rect 59164 3388 59220 3444
rect 59948 4226 60004 4228
rect 59948 4174 59950 4226
rect 59950 4174 60002 4226
rect 60002 4174 60004 4226
rect 59948 4172 60004 4174
rect 59724 3724 59780 3780
rect 60396 3612 60452 3668
rect 60956 5180 61012 5236
rect 62076 6300 62132 6356
rect 61516 6188 61572 6244
rect 62860 6188 62916 6244
rect 62076 5234 62132 5236
rect 62076 5182 62078 5234
rect 62078 5182 62130 5234
rect 62130 5182 62132 5234
rect 62076 5180 62132 5182
rect 61740 3724 61796 3780
rect 61852 4172 61908 4228
rect 61292 3500 61348 3556
rect 63308 60060 63364 60116
rect 63308 57708 63364 57764
rect 63756 62578 63812 62580
rect 63756 62526 63758 62578
rect 63758 62526 63810 62578
rect 63810 62526 63812 62578
rect 63756 62524 63812 62526
rect 63980 62354 64036 62356
rect 63980 62302 63982 62354
rect 63982 62302 64034 62354
rect 64034 62302 64036 62354
rect 63980 62300 64036 62302
rect 63644 60396 63700 60452
rect 63756 61628 63812 61684
rect 63532 6300 63588 6356
rect 63196 4284 63252 4340
rect 62972 4226 63028 4228
rect 62972 4174 62974 4226
rect 62974 4174 63026 4226
rect 63026 4174 63028 4226
rect 62972 4172 63028 4174
rect 63084 3666 63140 3668
rect 63084 3614 63086 3666
rect 63086 3614 63138 3666
rect 63138 3614 63140 3666
rect 63084 3612 63140 3614
rect 62524 3500 62580 3556
rect 64428 62242 64484 62244
rect 64428 62190 64430 62242
rect 64430 62190 64482 62242
rect 64482 62190 64484 62242
rect 64428 62188 64484 62190
rect 64540 60674 64596 60676
rect 64540 60622 64542 60674
rect 64542 60622 64594 60674
rect 64594 60622 64596 60674
rect 64540 60620 64596 60622
rect 64428 60562 64484 60564
rect 64428 60510 64430 60562
rect 64430 60510 64482 60562
rect 64482 60510 64484 60562
rect 64428 60508 64484 60510
rect 65324 64482 65380 64484
rect 65324 64430 65326 64482
rect 65326 64430 65378 64482
rect 65378 64430 65380 64482
rect 65324 64428 65380 64430
rect 65436 64092 65492 64148
rect 65548 64540 65604 64596
rect 65324 63868 65380 63924
rect 65772 64876 65828 64932
rect 66444 64988 66500 65044
rect 66332 64204 66388 64260
rect 65772 64146 65828 64148
rect 65772 64094 65774 64146
rect 65774 64094 65826 64146
rect 65826 64094 65828 64146
rect 65772 64092 65828 64094
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 65996 62914 66052 62916
rect 65996 62862 65998 62914
rect 65998 62862 66050 62914
rect 66050 62862 66052 62914
rect 65996 62860 66052 62862
rect 67116 65100 67172 65156
rect 66892 64540 66948 64596
rect 66668 64204 66724 64260
rect 66668 63922 66724 63924
rect 66668 63870 66670 63922
rect 66670 63870 66722 63922
rect 66722 63870 66724 63922
rect 66668 63868 66724 63870
rect 66668 62860 66724 62916
rect 67004 62914 67060 62916
rect 67004 62862 67006 62914
rect 67006 62862 67058 62914
rect 67058 62862 67060 62914
rect 67004 62860 67060 62862
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 65324 60674 65380 60676
rect 65324 60622 65326 60674
rect 65326 60622 65378 60674
rect 65378 60622 65380 60674
rect 65324 60620 65380 60622
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 66556 60172 66612 60228
rect 66444 60002 66500 60004
rect 66444 59950 66446 60002
rect 66446 59950 66498 60002
rect 66498 59950 66500 60002
rect 66444 59948 66500 59950
rect 64204 6188 64260 6244
rect 63756 4396 63812 4452
rect 63868 4338 63924 4340
rect 63868 4286 63870 4338
rect 63870 4286 63922 4338
rect 63922 4286 63924 4338
rect 63868 4284 63924 4286
rect 63756 4060 63812 4116
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 66668 49138 66724 49140
rect 66668 49086 66670 49138
rect 66670 49086 66722 49138
rect 66722 49086 66724 49138
rect 66668 49084 66724 49086
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 66780 6412 66836 6468
rect 65436 6188 65492 6244
rect 65772 6300 65828 6356
rect 64540 4338 64596 4340
rect 64540 4286 64542 4338
rect 64542 4286 64594 4338
rect 64594 4286 64596 4338
rect 64540 4284 64596 4286
rect 64428 3388 64484 3444
rect 66332 6188 66388 6244
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 66780 6188 66836 6244
rect 66556 5180 66612 5236
rect 65772 4172 65828 4228
rect 65212 3500 65268 3556
rect 66108 4060 66164 4116
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 66444 3442 66500 3444
rect 66444 3390 66446 3442
rect 66446 3390 66498 3442
rect 66498 3390 66500 3442
rect 66444 3388 66500 3390
rect 67340 64594 67396 64596
rect 67340 64542 67342 64594
rect 67342 64542 67394 64594
rect 67394 64542 67396 64594
rect 67340 64540 67396 64542
rect 67340 63922 67396 63924
rect 67340 63870 67342 63922
rect 67342 63870 67394 63922
rect 67394 63870 67396 63922
rect 67340 63868 67396 63870
rect 67116 60172 67172 60228
rect 68460 68124 68516 68180
rect 68124 67058 68180 67060
rect 68124 67006 68126 67058
rect 68126 67006 68178 67058
rect 68178 67006 68180 67058
rect 68124 67004 68180 67006
rect 68236 66946 68292 66948
rect 68236 66894 68238 66946
rect 68238 66894 68290 66946
rect 68290 66894 68292 66946
rect 68236 66892 68292 66894
rect 67788 66220 67844 66276
rect 68348 66498 68404 66500
rect 68348 66446 68350 66498
rect 68350 66446 68402 66498
rect 68402 66446 68404 66498
rect 68348 66444 68404 66446
rect 68236 66220 68292 66276
rect 67676 65436 67732 65492
rect 67676 64146 67732 64148
rect 67676 64094 67678 64146
rect 67678 64094 67730 64146
rect 67730 64094 67732 64146
rect 67676 64092 67732 64094
rect 67116 49138 67172 49140
rect 67116 49086 67118 49138
rect 67118 49086 67170 49138
rect 67170 49086 67172 49138
rect 67116 49084 67172 49086
rect 67228 48802 67284 48804
rect 67228 48750 67230 48802
rect 67230 48750 67282 48802
rect 67282 48750 67284 48802
rect 67228 48748 67284 48750
rect 67676 6636 67732 6692
rect 67004 6188 67060 6244
rect 67116 6412 67172 6468
rect 67340 6188 67396 6244
rect 67228 5740 67284 5796
rect 68012 65490 68068 65492
rect 68012 65438 68014 65490
rect 68014 65438 68066 65490
rect 68066 65438 68068 65490
rect 68012 65436 68068 65438
rect 68124 65378 68180 65380
rect 68124 65326 68126 65378
rect 68126 65326 68178 65378
rect 68178 65326 68180 65378
rect 68124 65324 68180 65326
rect 68012 64092 68068 64148
rect 68124 64988 68180 65044
rect 68236 64540 68292 64596
rect 68684 65548 68740 65604
rect 68796 65324 68852 65380
rect 71820 73164 71876 73220
rect 69692 72380 69748 72436
rect 70140 72434 70196 72436
rect 70140 72382 70142 72434
rect 70142 72382 70194 72434
rect 70194 72382 70196 72434
rect 70140 72380 70196 72382
rect 72156 72546 72212 72548
rect 72156 72494 72158 72546
rect 72158 72494 72210 72546
rect 72210 72494 72212 72546
rect 72156 72492 72212 72494
rect 72380 72492 72436 72548
rect 69468 72322 69524 72324
rect 69468 72270 69470 72322
rect 69470 72270 69522 72322
rect 69522 72270 69524 72322
rect 69468 72268 69524 72270
rect 69580 71932 69636 71988
rect 74956 75068 75012 75124
rect 73836 73442 73892 73444
rect 73836 73390 73838 73442
rect 73838 73390 73890 73442
rect 73890 73390 73892 73442
rect 73836 73388 73892 73390
rect 73612 73106 73668 73108
rect 73612 73054 73614 73106
rect 73614 73054 73666 73106
rect 73666 73054 73668 73106
rect 73612 73052 73668 73054
rect 73612 72604 73668 72660
rect 73052 72546 73108 72548
rect 73052 72494 73054 72546
rect 73054 72494 73106 72546
rect 73106 72494 73108 72546
rect 73052 72492 73108 72494
rect 71260 71874 71316 71876
rect 71260 71822 71262 71874
rect 71262 71822 71314 71874
rect 71314 71822 71316 71874
rect 71260 71820 71316 71822
rect 71596 71874 71652 71876
rect 71596 71822 71598 71874
rect 71598 71822 71650 71874
rect 71650 71822 71652 71874
rect 71596 71820 71652 71822
rect 72268 71820 72324 71876
rect 70812 71762 70868 71764
rect 70812 71710 70814 71762
rect 70814 71710 70866 71762
rect 70866 71710 70868 71762
rect 70812 71708 70868 71710
rect 71932 71708 71988 71764
rect 70588 71596 70644 71652
rect 70140 70866 70196 70868
rect 70140 70814 70142 70866
rect 70142 70814 70194 70866
rect 70194 70814 70196 70866
rect 70140 70812 70196 70814
rect 70700 71260 70756 71316
rect 69916 70306 69972 70308
rect 69916 70254 69918 70306
rect 69918 70254 69970 70306
rect 69970 70254 69972 70306
rect 69916 70252 69972 70254
rect 69468 70194 69524 70196
rect 69468 70142 69470 70194
rect 69470 70142 69522 70194
rect 69522 70142 69524 70194
rect 69468 70140 69524 70142
rect 70252 70194 70308 70196
rect 70252 70142 70254 70194
rect 70254 70142 70306 70194
rect 70306 70142 70308 70194
rect 70252 70140 70308 70142
rect 69580 70028 69636 70084
rect 69356 69186 69412 69188
rect 69356 69134 69358 69186
rect 69358 69134 69410 69186
rect 69410 69134 69412 69186
rect 69356 69132 69412 69134
rect 69692 69298 69748 69300
rect 69692 69246 69694 69298
rect 69694 69246 69746 69298
rect 69746 69246 69748 69298
rect 69692 69244 69748 69246
rect 70252 69298 70308 69300
rect 70252 69246 70254 69298
rect 70254 69246 70306 69298
rect 70306 69246 70308 69298
rect 70252 69244 70308 69246
rect 70924 70866 70980 70868
rect 70924 70814 70926 70866
rect 70926 70814 70978 70866
rect 70978 70814 70980 70866
rect 70924 70812 70980 70814
rect 71596 70866 71652 70868
rect 71596 70814 71598 70866
rect 71598 70814 71650 70866
rect 71650 70814 71652 70866
rect 71596 70812 71652 70814
rect 72268 70700 72324 70756
rect 72380 70812 72436 70868
rect 71260 70588 71316 70644
rect 70924 70194 70980 70196
rect 70924 70142 70926 70194
rect 70926 70142 70978 70194
rect 70978 70142 70980 70194
rect 70924 70140 70980 70142
rect 69580 68236 69636 68292
rect 69356 66444 69412 66500
rect 69244 65548 69300 65604
rect 68236 62466 68292 62468
rect 68236 62414 68238 62466
rect 68238 62414 68290 62466
rect 68290 62414 68292 62466
rect 68236 62412 68292 62414
rect 68124 62242 68180 62244
rect 68124 62190 68126 62242
rect 68126 62190 68178 62242
rect 68178 62190 68180 62242
rect 68124 62188 68180 62190
rect 68684 62466 68740 62468
rect 68684 62414 68686 62466
rect 68686 62414 68738 62466
rect 68738 62414 68740 62466
rect 68684 62412 68740 62414
rect 68572 49026 68628 49028
rect 68572 48974 68574 49026
rect 68574 48974 68626 49026
rect 68626 48974 68628 49026
rect 68572 48972 68628 48974
rect 68348 48860 68404 48916
rect 67900 48636 67956 48692
rect 68124 48802 68180 48804
rect 68124 48750 68126 48802
rect 68126 48750 68178 48802
rect 68178 48750 68180 48802
rect 68124 48748 68180 48750
rect 68012 5794 68068 5796
rect 68012 5742 68014 5794
rect 68014 5742 68066 5794
rect 68066 5742 68068 5794
rect 68012 5740 68068 5742
rect 67788 5516 67844 5572
rect 68684 6690 68740 6692
rect 68684 6638 68686 6690
rect 68686 6638 68738 6690
rect 68738 6638 68740 6690
rect 68684 6636 68740 6638
rect 69356 64092 69412 64148
rect 69468 49138 69524 49140
rect 69468 49086 69470 49138
rect 69470 49086 69522 49138
rect 69522 49086 69524 49138
rect 69468 49084 69524 49086
rect 69356 49026 69412 49028
rect 69356 48974 69358 49026
rect 69358 48974 69410 49026
rect 69410 48974 69412 49026
rect 69356 48972 69412 48974
rect 68908 48636 68964 48692
rect 69356 6690 69412 6692
rect 69356 6638 69358 6690
rect 69358 6638 69410 6690
rect 69410 6638 69412 6690
rect 69356 6636 69412 6638
rect 68796 5852 68852 5908
rect 68124 5404 68180 5460
rect 67788 5234 67844 5236
rect 67788 5182 67790 5234
rect 67790 5182 67842 5234
rect 67842 5182 67844 5234
rect 67788 5180 67844 5182
rect 68012 5180 68068 5236
rect 66892 4284 66948 4340
rect 67452 4396 67508 4452
rect 67340 4226 67396 4228
rect 67340 4174 67342 4226
rect 67342 4174 67394 4226
rect 67394 4174 67396 4226
rect 67340 4172 67396 4174
rect 67452 3612 67508 3668
rect 68460 5068 68516 5124
rect 68236 4338 68292 4340
rect 68236 4286 68238 4338
rect 68238 4286 68290 4338
rect 68290 4286 68292 4338
rect 68236 4284 68292 4286
rect 68348 3666 68404 3668
rect 68348 3614 68350 3666
rect 68350 3614 68402 3666
rect 68402 3614 68404 3666
rect 68348 3612 68404 3614
rect 69244 5068 69300 5124
rect 69356 5516 69412 5572
rect 68908 4338 68964 4340
rect 68908 4286 68910 4338
rect 68910 4286 68962 4338
rect 68962 4286 68964 4338
rect 68908 4284 68964 4286
rect 69132 3724 69188 3780
rect 70028 48914 70084 48916
rect 70028 48862 70030 48914
rect 70030 48862 70082 48914
rect 70082 48862 70084 48914
rect 70028 48860 70084 48862
rect 70140 5906 70196 5908
rect 70140 5854 70142 5906
rect 70142 5854 70194 5906
rect 70194 5854 70196 5906
rect 70140 5852 70196 5854
rect 70812 5906 70868 5908
rect 70812 5854 70814 5906
rect 70814 5854 70866 5906
rect 70866 5854 70868 5906
rect 70812 5852 70868 5854
rect 70140 5234 70196 5236
rect 70140 5182 70142 5234
rect 70142 5182 70194 5234
rect 70194 5182 70196 5234
rect 70140 5180 70196 5182
rect 70028 3724 70084 3780
rect 69916 3612 69972 3668
rect 71708 70194 71764 70196
rect 71708 70142 71710 70194
rect 71710 70142 71762 70194
rect 71762 70142 71764 70194
rect 71708 70140 71764 70142
rect 71148 69298 71204 69300
rect 71148 69246 71150 69298
rect 71150 69246 71202 69298
rect 71202 69246 71204 69298
rect 71148 69244 71204 69246
rect 72156 50706 72212 50708
rect 72156 50654 72158 50706
rect 72158 50654 72210 50706
rect 72210 50654 72212 50706
rect 72156 50652 72212 50654
rect 70924 4172 70980 4228
rect 71260 3666 71316 3668
rect 71260 3614 71262 3666
rect 71262 3614 71314 3666
rect 71314 3614 71316 3666
rect 71260 3612 71316 3614
rect 71148 3388 71204 3444
rect 71932 4226 71988 4228
rect 71932 4174 71934 4226
rect 71934 4174 71986 4226
rect 71986 4174 71988 4226
rect 71932 4172 71988 4174
rect 72828 70754 72884 70756
rect 72828 70702 72830 70754
rect 72830 70702 72882 70754
rect 72882 70702 72884 70754
rect 72828 70700 72884 70702
rect 72940 69522 72996 69524
rect 72940 69470 72942 69522
rect 72942 69470 72994 69522
rect 72994 69470 72996 69522
rect 72940 69468 72996 69470
rect 72940 64818 72996 64820
rect 72940 64766 72942 64818
rect 72942 64766 72994 64818
rect 72994 64766 72996 64818
rect 72940 64764 72996 64766
rect 72940 59836 72996 59892
rect 72604 50706 72660 50708
rect 72604 50654 72606 50706
rect 72606 50654 72658 50706
rect 72658 50654 72660 50706
rect 72604 50652 72660 50654
rect 72716 49980 72772 50036
rect 72604 49756 72660 49812
rect 72604 48860 72660 48916
rect 73052 48636 73108 48692
rect 72492 4396 72548 4452
rect 73500 72492 73556 72548
rect 73276 72434 73332 72436
rect 73276 72382 73278 72434
rect 73278 72382 73330 72434
rect 73330 72382 73332 72434
rect 73276 72380 73332 72382
rect 75516 74508 75572 74564
rect 74172 72658 74228 72660
rect 74172 72606 74174 72658
rect 74174 72606 74226 72658
rect 74226 72606 74228 72658
rect 74172 72604 74228 72606
rect 73836 72268 73892 72324
rect 73388 71986 73444 71988
rect 73388 71934 73390 71986
rect 73390 71934 73442 71986
rect 73442 71934 73444 71986
rect 73388 71932 73444 71934
rect 73948 71932 74004 71988
rect 74060 72268 74116 72324
rect 73276 70700 73332 70756
rect 74396 70754 74452 70756
rect 74396 70702 74398 70754
rect 74398 70702 74450 70754
rect 74450 70702 74452 70754
rect 74396 70700 74452 70702
rect 73500 50706 73556 50708
rect 73500 50654 73502 50706
rect 73502 50654 73554 50706
rect 73554 50654 73556 50706
rect 73500 50652 73556 50654
rect 73612 49810 73668 49812
rect 73612 49758 73614 49810
rect 73614 49758 73666 49810
rect 73666 49758 73668 49810
rect 73612 49756 73668 49758
rect 73388 4396 73444 4452
rect 74172 70476 74228 70532
rect 76300 74002 76356 74004
rect 76300 73950 76302 74002
rect 76302 73950 76354 74002
rect 76354 73950 76356 74002
rect 76300 73948 76356 73950
rect 74956 73330 75012 73332
rect 74956 73278 74958 73330
rect 74958 73278 75010 73330
rect 75010 73278 75012 73330
rect 74956 73276 75012 73278
rect 77308 74002 77364 74004
rect 77308 73950 77310 74002
rect 77310 73950 77362 74002
rect 77362 73950 77364 74002
rect 77308 73948 77364 73950
rect 75516 73164 75572 73220
rect 74956 71260 75012 71316
rect 74844 70476 74900 70532
rect 75964 71820 76020 71876
rect 75068 70588 75124 70644
rect 75404 70700 75460 70756
rect 74956 70028 75012 70084
rect 74956 69356 75012 69412
rect 74284 69132 74340 69188
rect 74508 69132 74564 69188
rect 75068 68236 75124 68292
rect 74956 67954 75012 67956
rect 74956 67902 74958 67954
rect 74958 67902 75010 67954
rect 75010 67902 75012 67954
rect 74956 67900 75012 67902
rect 75180 67116 75236 67172
rect 74956 64988 75012 65044
rect 74284 64428 74340 64484
rect 74508 64428 74564 64484
rect 75180 65100 75236 65156
rect 75068 64652 75124 64708
rect 74956 64316 75012 64372
rect 74620 60620 74676 60676
rect 74284 59724 74340 59780
rect 74508 59724 74564 59780
rect 74732 59164 74788 59220
rect 75180 61292 75236 61348
rect 75068 60172 75124 60228
rect 74956 60114 75012 60116
rect 74956 60062 74958 60114
rect 74958 60062 75010 60114
rect 75010 60062 75012 60114
rect 74956 60060 75012 60062
rect 74844 58156 74900 58212
rect 74956 56978 75012 56980
rect 74956 56926 74958 56978
rect 74958 56926 75010 56978
rect 75010 56926 75012 56978
rect 74956 56924 75012 56926
rect 75180 56700 75236 56756
rect 75068 56252 75124 56308
rect 75068 54684 75124 54740
rect 74844 54572 74900 54628
rect 75068 53900 75124 53956
rect 74956 53842 75012 53844
rect 74956 53790 74958 53842
rect 74958 53790 75010 53842
rect 75010 53790 75012 53842
rect 74956 53788 75012 53790
rect 75180 52780 75236 52836
rect 75068 52108 75124 52164
rect 74060 50706 74116 50708
rect 74060 50654 74062 50706
rect 74062 50654 74114 50706
rect 74114 50654 74116 50706
rect 74060 50652 74116 50654
rect 73836 50034 73892 50036
rect 73836 49982 73838 50034
rect 73838 49982 73890 50034
rect 73890 49982 73892 50034
rect 73836 49980 73892 49982
rect 75180 50540 75236 50596
rect 75068 49644 75124 49700
rect 74844 49196 74900 49252
rect 74956 49138 75012 49140
rect 74956 49086 74958 49138
rect 74958 49086 75010 49138
rect 75010 49086 75012 49138
rect 74956 49084 75012 49086
rect 74060 48636 74116 48692
rect 74284 46956 74340 47012
rect 75180 47292 75236 47348
rect 74956 46956 75012 47012
rect 74508 46844 74564 46900
rect 74284 45724 74340 45780
rect 74396 45666 74452 45668
rect 74396 45614 74398 45666
rect 74398 45614 74450 45666
rect 74450 45614 74452 45666
rect 74396 45612 74452 45614
rect 74956 45612 75012 45668
rect 74508 45276 74564 45332
rect 74508 44044 74564 44100
rect 74396 43708 74452 43764
rect 74956 43708 75012 43764
rect 74396 42700 74452 42756
rect 74956 42754 75012 42756
rect 74956 42702 74958 42754
rect 74958 42702 75010 42754
rect 75010 42702 75012 42754
rect 74956 42700 75012 42702
rect 74508 42476 74564 42532
rect 74396 42028 74452 42084
rect 74396 41132 74452 41188
rect 74956 41186 75012 41188
rect 74956 41134 74958 41186
rect 74958 41134 75010 41186
rect 75010 41134 75012 41186
rect 74956 41132 75012 41134
rect 74508 40908 74564 40964
rect 74396 40460 74452 40516
rect 74508 39564 74564 39620
rect 74508 39394 74564 39396
rect 74508 39342 74510 39394
rect 74510 39342 74562 39394
rect 74562 39342 74564 39394
rect 74508 39340 74564 39342
rect 74956 39340 75012 39396
rect 74508 38946 74564 38948
rect 74508 38894 74510 38946
rect 74510 38894 74562 38946
rect 74562 38894 74564 38946
rect 74508 38892 74564 38894
rect 74956 38892 75012 38948
rect 74508 37826 74564 37828
rect 74508 37774 74510 37826
rect 74510 37774 74562 37826
rect 74562 37774 74564 37826
rect 74508 37772 74564 37774
rect 74956 37772 75012 37828
rect 74508 37378 74564 37380
rect 74508 37326 74510 37378
rect 74510 37326 74562 37378
rect 74562 37326 74564 37378
rect 74508 37324 74564 37326
rect 74956 37324 75012 37380
rect 74508 36258 74564 36260
rect 74508 36206 74510 36258
rect 74510 36206 74562 36258
rect 74562 36206 74564 36258
rect 74508 36204 74564 36206
rect 74956 36204 75012 36260
rect 74508 35810 74564 35812
rect 74508 35758 74510 35810
rect 74510 35758 74562 35810
rect 74562 35758 74564 35810
rect 74508 35756 74564 35758
rect 74956 35756 75012 35812
rect 74508 34802 74564 34804
rect 74508 34750 74510 34802
rect 74510 34750 74562 34802
rect 74562 34750 74564 34802
rect 74508 34748 74564 34750
rect 74956 34748 75012 34804
rect 74508 34242 74564 34244
rect 74508 34190 74510 34242
rect 74510 34190 74562 34242
rect 74562 34190 74564 34242
rect 74508 34188 74564 34190
rect 74956 34188 75012 34244
rect 74508 33122 74564 33124
rect 74508 33070 74510 33122
rect 74510 33070 74562 33122
rect 74562 33070 74564 33122
rect 74508 33068 74564 33070
rect 74956 33068 75012 33124
rect 74508 32674 74564 32676
rect 74508 32622 74510 32674
rect 74510 32622 74562 32674
rect 74562 32622 74564 32674
rect 74508 32620 74564 32622
rect 74956 32620 75012 32676
rect 74508 31554 74564 31556
rect 74508 31502 74510 31554
rect 74510 31502 74562 31554
rect 74562 31502 74564 31554
rect 74508 31500 74564 31502
rect 74956 31500 75012 31556
rect 74508 31106 74564 31108
rect 74508 31054 74510 31106
rect 74510 31054 74562 31106
rect 74562 31054 74564 31106
rect 74508 31052 74564 31054
rect 74956 31052 75012 31108
rect 74508 30098 74564 30100
rect 74508 30046 74510 30098
rect 74510 30046 74562 30098
rect 74562 30046 74564 30098
rect 74508 30044 74564 30046
rect 74956 30044 75012 30100
rect 74508 29538 74564 29540
rect 74508 29486 74510 29538
rect 74510 29486 74562 29538
rect 74562 29486 74564 29538
rect 74508 29484 74564 29486
rect 74956 29484 75012 29540
rect 74508 28364 74564 28420
rect 74956 28364 75012 28420
rect 74508 27970 74564 27972
rect 74508 27918 74510 27970
rect 74510 27918 74562 27970
rect 74562 27918 74564 27970
rect 74508 27916 74564 27918
rect 74956 27916 75012 27972
rect 74508 26796 74564 26852
rect 74956 26796 75012 26852
rect 74508 26402 74564 26404
rect 74508 26350 74510 26402
rect 74510 26350 74562 26402
rect 74562 26350 74564 26402
rect 74508 26348 74564 26350
rect 74956 26348 75012 26404
rect 74508 25282 74564 25284
rect 74508 25230 74510 25282
rect 74510 25230 74562 25282
rect 74562 25230 74564 25282
rect 74508 25228 74564 25230
rect 74956 25228 75012 25284
rect 74508 24722 74564 24724
rect 74508 24670 74510 24722
rect 74510 24670 74562 24722
rect 74562 24670 74564 24722
rect 74508 24668 74564 24670
rect 74956 24722 75012 24724
rect 74956 24670 74958 24722
rect 74958 24670 75010 24722
rect 75010 24670 75012 24722
rect 74956 24668 75012 24670
rect 74508 23714 74564 23716
rect 74508 23662 74510 23714
rect 74510 23662 74562 23714
rect 74562 23662 74564 23714
rect 74508 23660 74564 23662
rect 74956 23660 75012 23716
rect 74508 23266 74564 23268
rect 74508 23214 74510 23266
rect 74510 23214 74562 23266
rect 74562 23214 74564 23266
rect 74508 23212 74564 23214
rect 74956 23212 75012 23268
rect 74508 22146 74564 22148
rect 74508 22094 74510 22146
rect 74510 22094 74562 22146
rect 74562 22094 74564 22146
rect 74508 22092 74564 22094
rect 74956 22092 75012 22148
rect 74508 21698 74564 21700
rect 74508 21646 74510 21698
rect 74510 21646 74562 21698
rect 74562 21646 74564 21698
rect 74508 21644 74564 21646
rect 74956 21644 75012 21700
rect 74508 20578 74564 20580
rect 74508 20526 74510 20578
rect 74510 20526 74562 20578
rect 74562 20526 74564 20578
rect 74508 20524 74564 20526
rect 74956 20524 75012 20580
rect 73500 4956 73556 5012
rect 74508 19122 74564 19124
rect 74508 19070 74510 19122
rect 74510 19070 74562 19122
rect 74562 19070 74564 19122
rect 74508 19068 74564 19070
rect 74956 19068 75012 19124
rect 74396 18956 74452 19012
rect 74508 18450 74564 18452
rect 74508 18398 74510 18450
rect 74510 18398 74562 18450
rect 74562 18398 74564 18450
rect 74508 18396 74564 18398
rect 74956 18450 75012 18452
rect 74956 18398 74958 18450
rect 74958 18398 75010 18450
rect 75010 18398 75012 18450
rect 74956 18396 75012 18398
rect 74508 17554 74564 17556
rect 74508 17502 74510 17554
rect 74510 17502 74562 17554
rect 74562 17502 74564 17554
rect 74508 17500 74564 17502
rect 74956 17500 75012 17556
rect 74508 16994 74564 16996
rect 74508 16942 74510 16994
rect 74510 16942 74562 16994
rect 74562 16942 74564 16994
rect 74508 16940 74564 16942
rect 74956 16940 75012 16996
rect 74508 16098 74564 16100
rect 74508 16046 74510 16098
rect 74510 16046 74562 16098
rect 74562 16046 74564 16098
rect 74508 16044 74564 16046
rect 74956 16098 75012 16100
rect 74956 16046 74958 16098
rect 74958 16046 75010 16098
rect 75010 16046 75012 16098
rect 74956 16044 75012 16046
rect 74508 15426 74564 15428
rect 74508 15374 74510 15426
rect 74510 15374 74562 15426
rect 74562 15374 74564 15426
rect 74508 15372 74564 15374
rect 74956 15372 75012 15428
rect 74508 14306 74564 14308
rect 74508 14254 74510 14306
rect 74510 14254 74562 14306
rect 74562 14254 74564 14306
rect 74508 14252 74564 14254
rect 74956 14252 75012 14308
rect 74508 13858 74564 13860
rect 74508 13806 74510 13858
rect 74510 13806 74562 13858
rect 74562 13806 74564 13858
rect 74508 13804 74564 13806
rect 74956 13804 75012 13860
rect 74396 13692 74452 13748
rect 74508 12290 74564 12292
rect 74508 12238 74510 12290
rect 74510 12238 74562 12290
rect 74562 12238 74564 12290
rect 74508 12236 74564 12238
rect 74956 12236 75012 12292
rect 74508 11282 74564 11284
rect 74508 11230 74510 11282
rect 74510 11230 74562 11282
rect 74562 11230 74564 11282
rect 74508 11228 74564 11230
rect 74956 11228 75012 11284
rect 74508 10722 74564 10724
rect 74508 10670 74510 10722
rect 74510 10670 74562 10722
rect 74562 10670 74564 10722
rect 74508 10668 74564 10670
rect 74956 10668 75012 10724
rect 74508 9602 74564 9604
rect 74508 9550 74510 9602
rect 74510 9550 74562 9602
rect 74562 9550 74564 9602
rect 74508 9548 74564 9550
rect 74956 9548 75012 9604
rect 74508 9154 74564 9156
rect 74508 9102 74510 9154
rect 74510 9102 74562 9154
rect 74562 9102 74564 9154
rect 74508 9100 74564 9102
rect 74956 9100 75012 9156
rect 74508 8034 74564 8036
rect 74508 7982 74510 8034
rect 74510 7982 74562 8034
rect 74562 7982 74564 8034
rect 74508 7980 74564 7982
rect 74956 7980 75012 8036
rect 74508 7586 74564 7588
rect 74508 7534 74510 7586
rect 74510 7534 74562 7586
rect 74562 7534 74564 7586
rect 74508 7532 74564 7534
rect 74956 7532 75012 7588
rect 74508 6076 74564 6132
rect 74956 6076 75012 6132
rect 75068 5010 75124 5012
rect 75068 4958 75070 5010
rect 75070 4958 75122 5010
rect 75122 4958 75124 5010
rect 75068 4956 75124 4958
rect 74508 4508 74564 4564
rect 74396 4450 74452 4452
rect 74396 4398 74398 4450
rect 74398 4398 74450 4450
rect 74450 4398 74452 4450
rect 74396 4396 74452 4398
rect 77868 72492 77924 72548
rect 76748 72380 76804 72436
rect 76748 71762 76804 71764
rect 76748 71710 76750 71762
rect 76750 71710 76802 71762
rect 76802 71710 76804 71762
rect 76748 71708 76804 71710
rect 77868 71148 77924 71204
rect 76300 70866 76356 70868
rect 76300 70814 76302 70866
rect 76302 70814 76354 70866
rect 76354 70814 76356 70866
rect 76300 70812 76356 70814
rect 77308 70812 77364 70868
rect 76076 70588 76132 70644
rect 75516 69804 75572 69860
rect 76300 69298 76356 69300
rect 76300 69246 76302 69298
rect 76302 69246 76354 69298
rect 76354 69246 76356 69298
rect 76300 69244 76356 69246
rect 76300 68738 76356 68740
rect 76300 68686 76302 68738
rect 76302 68686 76354 68738
rect 76354 68686 76356 68738
rect 76300 68684 76356 68686
rect 77308 69244 77364 69300
rect 76860 68684 76916 68740
rect 76748 67788 76804 67844
rect 76300 67730 76356 67732
rect 76300 67678 76302 67730
rect 76302 67678 76354 67730
rect 76354 67678 76356 67730
rect 76300 67676 76356 67678
rect 76300 67170 76356 67172
rect 76300 67118 76302 67170
rect 76302 67118 76354 67170
rect 76354 67118 76356 67170
rect 76300 67116 76356 67118
rect 76860 67116 76916 67172
rect 76300 65996 76356 66052
rect 77308 67730 77364 67732
rect 77308 67678 77310 67730
rect 77310 67678 77362 67730
rect 77362 67678 77364 67730
rect 77308 67676 77364 67678
rect 77532 68460 77588 68516
rect 77420 67116 77476 67172
rect 76972 66444 77028 66500
rect 76860 65548 76916 65604
rect 77308 66050 77364 66052
rect 77308 65998 77310 66050
rect 77310 65998 77362 66050
rect 77362 65998 77364 66050
rect 77308 65996 77364 65998
rect 77420 65772 77476 65828
rect 76300 64594 76356 64596
rect 76300 64542 76302 64594
rect 76302 64542 76354 64594
rect 76354 64542 76356 64594
rect 76300 64540 76356 64542
rect 76300 63756 76356 63812
rect 77308 64540 77364 64596
rect 76860 63756 76916 63812
rect 76748 63084 76804 63140
rect 76300 63026 76356 63028
rect 76300 62974 76302 63026
rect 76302 62974 76354 63026
rect 76354 62974 76356 63026
rect 76300 62972 76356 62974
rect 76300 61458 76356 61460
rect 76300 61406 76302 61458
rect 76302 61406 76354 61458
rect 76354 61406 76356 61458
rect 76300 61404 76356 61406
rect 77308 62972 77364 63028
rect 77532 63868 77588 63924
rect 77420 62412 77476 62468
rect 77084 61740 77140 61796
rect 76972 60508 77028 60564
rect 77196 61404 77252 61460
rect 76300 59890 76356 59892
rect 76300 59838 76302 59890
rect 76302 59838 76354 59890
rect 76354 59838 76356 59890
rect 76300 59836 76356 59838
rect 76300 58322 76356 58324
rect 76300 58270 76302 58322
rect 76302 58270 76354 58322
rect 76354 58270 76356 58322
rect 76300 58268 76356 58270
rect 76300 57762 76356 57764
rect 76300 57710 76302 57762
rect 76302 57710 76354 57762
rect 76354 57710 76356 57762
rect 76300 57708 76356 57710
rect 77420 61068 77476 61124
rect 77308 59836 77364 59892
rect 77196 59052 77252 59108
rect 76972 58380 77028 58436
rect 77308 58268 77364 58324
rect 76860 57708 76916 57764
rect 77420 57708 77476 57764
rect 76748 57260 76804 57316
rect 76300 56754 76356 56756
rect 76300 56702 76302 56754
rect 76302 56702 76354 56754
rect 76354 56702 76356 56754
rect 76300 56700 76356 56702
rect 76300 56194 76356 56196
rect 76300 56142 76302 56194
rect 76302 56142 76354 56194
rect 76354 56142 76356 56194
rect 76300 56140 76356 56142
rect 76860 56194 76916 56196
rect 76860 56142 76862 56194
rect 76862 56142 76914 56194
rect 76914 56142 76916 56194
rect 76860 56140 76916 56142
rect 76972 55692 77028 55748
rect 77308 56700 77364 56756
rect 77420 56364 77476 56420
rect 77308 55468 77364 55524
rect 76300 55186 76356 55188
rect 76300 55134 76302 55186
rect 76302 55134 76354 55186
rect 76354 55134 76356 55186
rect 76300 55132 76356 55134
rect 76300 54626 76356 54628
rect 76300 54574 76302 54626
rect 76302 54574 76354 54626
rect 76354 54574 76356 54626
rect 76300 54572 76356 54574
rect 76860 54572 76916 54628
rect 76300 53618 76356 53620
rect 76300 53566 76302 53618
rect 76302 53566 76354 53618
rect 76354 53566 76356 53618
rect 76300 53564 76356 53566
rect 76972 54348 77028 54404
rect 77308 55132 77364 55188
rect 77308 53788 77364 53844
rect 76860 53228 76916 53284
rect 77308 53564 77364 53620
rect 76300 53058 76356 53060
rect 76300 53006 76302 53058
rect 76302 53006 76354 53058
rect 76354 53006 76356 53058
rect 76300 53004 76356 53006
rect 76860 53004 76916 53060
rect 76300 52050 76356 52052
rect 76300 51998 76302 52050
rect 76302 51998 76354 52050
rect 76354 51998 76356 52050
rect 76300 51996 76356 51998
rect 77308 52332 77364 52388
rect 76860 51660 76916 51716
rect 77308 51996 77364 52052
rect 76300 51490 76356 51492
rect 76300 51438 76302 51490
rect 76302 51438 76354 51490
rect 76354 51438 76356 51490
rect 76300 51436 76356 51438
rect 76860 51436 76916 51492
rect 76300 50482 76356 50484
rect 76300 50430 76302 50482
rect 76302 50430 76354 50482
rect 76354 50430 76356 50482
rect 76300 50428 76356 50430
rect 77308 50988 77364 51044
rect 76860 50316 76916 50372
rect 77308 50482 77364 50484
rect 77308 50430 77310 50482
rect 77310 50430 77362 50482
rect 77362 50430 77364 50482
rect 77308 50428 77364 50430
rect 76300 49922 76356 49924
rect 76300 49870 76302 49922
rect 76302 49870 76354 49922
rect 76354 49870 76356 49922
rect 76300 49868 76356 49870
rect 76860 49868 76916 49924
rect 77308 49644 77364 49700
rect 76860 48972 76916 49028
rect 76300 48914 76356 48916
rect 76300 48862 76302 48914
rect 76302 48862 76354 48914
rect 76354 48862 76356 48914
rect 76300 48860 76356 48862
rect 77308 48860 77364 48916
rect 77308 48300 77364 48356
rect 75964 47068 76020 47124
rect 77868 47628 77924 47684
rect 76748 47180 76804 47236
rect 77196 47234 77252 47236
rect 77196 47182 77198 47234
rect 77198 47182 77250 47234
rect 77250 47182 77252 47234
rect 77196 47180 77252 47182
rect 76076 46284 76132 46340
rect 75964 45612 76020 45668
rect 76076 44940 76132 44996
rect 75964 44268 76020 44324
rect 76076 43708 76132 43764
rect 76076 42924 76132 42980
rect 76076 42252 76132 42308
rect 76076 41580 76132 41636
rect 76076 40908 76132 40964
rect 76076 40402 76132 40404
rect 76076 40350 76078 40402
rect 76078 40350 76130 40402
rect 76130 40350 76132 40402
rect 76076 40348 76132 40350
rect 76076 39618 76132 39620
rect 76076 39566 76078 39618
rect 76078 39566 76130 39618
rect 76130 39566 76132 39618
rect 76076 39564 76132 39566
rect 76076 38946 76132 38948
rect 76076 38894 76078 38946
rect 76078 38894 76130 38946
rect 76130 38894 76132 38946
rect 76076 38892 76132 38894
rect 76076 38220 76132 38276
rect 76076 37548 76132 37604
rect 76076 36876 76132 36932
rect 76076 36204 76132 36260
rect 76076 35532 76132 35588
rect 77868 34860 77924 34916
rect 76748 34636 76804 34692
rect 77196 34690 77252 34692
rect 77196 34638 77198 34690
rect 77198 34638 77250 34690
rect 77250 34638 77252 34690
rect 77196 34636 77252 34638
rect 76076 34242 76132 34244
rect 76076 34190 76078 34242
rect 76078 34190 76130 34242
rect 76130 34190 76132 34242
rect 76076 34188 76132 34190
rect 76076 33516 76132 33572
rect 76076 32844 76132 32900
rect 76076 31890 76132 31892
rect 76076 31838 76078 31890
rect 76078 31838 76130 31890
rect 76130 31838 76132 31890
rect 76076 31836 76132 31838
rect 76076 31500 76132 31556
rect 76076 30828 76132 30884
rect 77868 30268 77924 30324
rect 76748 29932 76804 29988
rect 77196 29986 77252 29988
rect 77196 29934 77198 29986
rect 77198 29934 77250 29986
rect 77250 29934 77252 29986
rect 77196 29932 77252 29934
rect 76076 29538 76132 29540
rect 76076 29486 76078 29538
rect 76078 29486 76130 29538
rect 76130 29486 76132 29538
rect 76076 29484 76132 29486
rect 76076 28812 76132 28868
rect 76076 28140 76132 28196
rect 76076 27468 76132 27524
rect 76076 26796 76132 26852
rect 76076 26124 76132 26180
rect 77868 25452 77924 25508
rect 77196 24892 77252 24948
rect 76076 24834 76132 24836
rect 76076 24782 76078 24834
rect 76078 24782 76130 24834
rect 76130 24782 76132 24834
rect 76076 24780 76132 24782
rect 76076 24108 76132 24164
rect 76076 23436 76132 23492
rect 76076 22764 76132 22820
rect 76076 22092 76132 22148
rect 76076 21420 76132 21476
rect 77868 20748 77924 20804
rect 77196 20188 77252 20244
rect 76076 20130 76132 20132
rect 76076 20078 76078 20130
rect 76078 20078 76130 20130
rect 76130 20078 76132 20130
rect 76076 20076 76132 20078
rect 76076 19404 76132 19460
rect 76076 18732 76132 18788
rect 76076 18060 76132 18116
rect 76076 17388 76132 17444
rect 76076 16716 76132 16772
rect 77868 16044 77924 16100
rect 76748 15820 76804 15876
rect 77196 15874 77252 15876
rect 77196 15822 77198 15874
rect 77198 15822 77250 15874
rect 77250 15822 77252 15874
rect 77196 15820 77252 15822
rect 76076 15426 76132 15428
rect 76076 15374 76078 15426
rect 76078 15374 76130 15426
rect 76130 15374 76132 15426
rect 76076 15372 76132 15374
rect 76076 14700 76132 14756
rect 76076 14028 76132 14084
rect 76076 13356 76132 13412
rect 76076 12684 76132 12740
rect 76076 12012 76132 12068
rect 77868 11340 77924 11396
rect 76748 11116 76804 11172
rect 77196 11170 77252 11172
rect 77196 11118 77198 11170
rect 77198 11118 77250 11170
rect 77250 11118 77252 11170
rect 77196 11116 77252 11118
rect 76076 10722 76132 10724
rect 76076 10670 76078 10722
rect 76078 10670 76130 10722
rect 76130 10670 76132 10722
rect 76076 10668 76132 10670
rect 76076 9996 76132 10052
rect 76076 9324 76132 9380
rect 76076 8370 76132 8372
rect 76076 8318 76078 8370
rect 76078 8318 76130 8370
rect 76130 8318 76132 8370
rect 76076 8316 76132 8318
rect 76076 7980 76132 8036
rect 76076 7308 76132 7364
rect 77868 6748 77924 6804
rect 76748 6524 76804 6580
rect 77196 6578 77252 6580
rect 77196 6526 77198 6578
rect 77198 6526 77250 6578
rect 77250 6526 77252 6578
rect 77196 6524 77252 6526
rect 76076 6018 76132 6020
rect 76076 5966 76078 6018
rect 76078 5966 76130 6018
rect 76130 5966 76132 6018
rect 76076 5964 76132 5966
rect 77868 5292 77924 5348
rect 76524 4844 76580 4900
rect 74172 3724 74228 3780
rect 75628 3724 75684 3780
rect 72716 3388 72772 3444
rect 73836 3612 73892 3668
rect 73388 3442 73444 3444
rect 73388 3390 73390 3442
rect 73390 3390 73442 3442
rect 73442 3390 73444 3442
rect 73388 3388 73444 3390
rect 76300 3724 76356 3780
rect 74508 3388 74564 3444
rect 75068 3442 75124 3444
rect 75068 3390 75070 3442
rect 75070 3390 75122 3442
rect 75122 3390 75124 3442
rect 75068 3388 75124 3390
rect 76972 3666 77028 3668
rect 76972 3614 76974 3666
rect 76974 3614 77026 3666
rect 77026 3614 77028 3666
rect 76972 3612 77028 3614
rect 76412 3388 76468 3444
<< metal3 >>
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 73714 75068 73724 75124
rect 73780 75068 74956 75124
rect 75012 75068 75022 75124
rect 3042 74844 3052 74900
rect 3108 74844 3612 74900
rect 3668 74844 3678 74900
rect 0 74564 800 74592
rect 79200 74564 80000 74592
rect 0 74508 2044 74564
rect 2100 74508 2110 74564
rect 75506 74508 75516 74564
rect 75572 74508 80000 74564
rect 0 74480 800 74508
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 79200 74480 80000 74508
rect 2258 73948 2268 74004
rect 2324 73948 4172 74004
rect 4228 73948 4238 74004
rect 76290 73948 76300 74004
rect 76356 73948 77308 74004
rect 77364 73948 77374 74004
rect 0 73892 800 73920
rect 2268 73892 2324 73948
rect 0 73836 2324 73892
rect 77308 73892 77364 73948
rect 79200 73892 80000 73920
rect 77308 73836 80000 73892
rect 0 73808 800 73836
rect 79200 73808 80000 73836
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 3490 73500 3500 73556
rect 3556 73500 68908 73556
rect 68964 73500 68974 73556
rect 69010 73388 69020 73444
rect 69076 73388 73836 73444
rect 73892 73388 73902 73444
rect 3042 73276 3052 73332
rect 3108 73276 3836 73332
rect 3892 73276 3902 73332
rect 72482 73276 72492 73332
rect 72548 73276 74956 73332
rect 75012 73276 75022 73332
rect 0 73220 800 73248
rect 79200 73220 80000 73248
rect 0 73164 1932 73220
rect 1988 73164 1998 73220
rect 4834 73164 4844 73220
rect 4900 73164 5404 73220
rect 5460 73164 71820 73220
rect 71876 73164 71886 73220
rect 75506 73164 75516 73220
rect 75572 73164 80000 73220
rect 0 73136 800 73164
rect 79200 73136 80000 73164
rect 68450 73052 68460 73108
rect 68516 73052 73612 73108
rect 73668 73052 73678 73108
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 3602 72604 3612 72660
rect 3668 72604 8428 72660
rect 73602 72604 73612 72660
rect 73668 72604 74172 72660
rect 74228 72604 74238 72660
rect 0 72548 800 72576
rect 0 72492 3724 72548
rect 3780 72492 3790 72548
rect 0 72464 800 72492
rect 8372 72324 8428 72604
rect 79200 72548 80000 72576
rect 72146 72492 72156 72548
rect 72212 72492 72380 72548
rect 72436 72492 73052 72548
rect 73108 72492 73500 72548
rect 73556 72492 73566 72548
rect 77858 72492 77868 72548
rect 77924 72492 80000 72548
rect 79200 72464 80000 72492
rect 69346 72380 69356 72436
rect 69412 72380 69692 72436
rect 69748 72380 70140 72436
rect 70196 72380 70206 72436
rect 73266 72380 73276 72436
rect 73332 72380 76748 72436
rect 76804 72380 76814 72436
rect 3042 72268 3052 72324
rect 3108 72268 3948 72324
rect 4004 72268 4014 72324
rect 8372 72268 69468 72324
rect 69524 72268 69534 72324
rect 73826 72268 73836 72324
rect 73892 72268 74060 72324
rect 74116 72268 74126 72324
rect 3826 72156 3836 72212
rect 3892 72156 8428 72212
rect 0 71876 800 71904
rect 8372 71876 8428 72156
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 69570 71932 69580 71988
rect 69636 71932 73388 71988
rect 73444 71932 73948 71988
rect 74004 71932 74014 71988
rect 79200 71876 80000 71904
rect 0 71820 2044 71876
rect 2100 71820 2110 71876
rect 8372 71820 71260 71876
rect 71316 71820 71326 71876
rect 71586 71820 71596 71876
rect 71652 71820 72268 71876
rect 72324 71820 72334 71876
rect 75954 71820 75964 71876
rect 76020 71820 80000 71876
rect 0 71792 800 71820
rect 71596 71764 71652 71820
rect 79200 71792 80000 71820
rect 3042 71708 3052 71764
rect 3108 71708 3612 71764
rect 3668 71708 3678 71764
rect 70802 71708 70812 71764
rect 70868 71708 71652 71764
rect 71922 71708 71932 71764
rect 71988 71708 76748 71764
rect 76804 71708 76814 71764
rect 4834 71596 4844 71652
rect 4900 71596 5404 71652
rect 5460 71596 70588 71652
rect 70644 71596 70654 71652
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 70690 71260 70700 71316
rect 70756 71260 74956 71316
rect 75012 71260 75022 71316
rect 0 71204 800 71232
rect 79200 71204 80000 71232
rect 0 71148 3724 71204
rect 3780 71148 3790 71204
rect 77858 71148 77868 71204
rect 77924 71148 80000 71204
rect 0 71120 800 71148
rect 79200 71120 80000 71148
rect 3378 70924 3388 70980
rect 3444 70924 3836 70980
rect 3892 70924 3902 70980
rect 70130 70812 70140 70868
rect 70196 70812 70924 70868
rect 70980 70812 71596 70868
rect 71652 70812 72380 70868
rect 72436 70812 72446 70868
rect 76290 70812 76300 70868
rect 76356 70812 77308 70868
rect 77364 70812 77374 70868
rect 2146 70700 2156 70756
rect 2212 70700 3724 70756
rect 3780 70700 3790 70756
rect 72258 70700 72268 70756
rect 72324 70700 72828 70756
rect 72884 70700 73276 70756
rect 73332 70700 73342 70756
rect 74386 70700 74396 70756
rect 74452 70700 75404 70756
rect 75460 70700 75470 70756
rect 71250 70588 71260 70644
rect 71316 70588 75068 70644
rect 75124 70588 75134 70644
rect 76066 70588 76076 70644
rect 76132 70588 76142 70644
rect 0 70532 800 70560
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 76076 70532 76132 70588
rect 79200 70532 80000 70560
rect 0 70476 1820 70532
rect 1876 70476 1886 70532
rect 74162 70476 74172 70532
rect 74228 70476 74844 70532
rect 74900 70476 74910 70532
rect 76076 70476 80000 70532
rect 0 70448 800 70476
rect 79200 70448 80000 70476
rect 1922 70252 1932 70308
rect 1988 70252 3724 70308
rect 3780 70252 3790 70308
rect 3938 70252 3948 70308
rect 4004 70252 69916 70308
rect 69972 70252 69982 70308
rect 69458 70140 69468 70196
rect 69524 70140 70252 70196
rect 70308 70140 70924 70196
rect 70980 70140 71708 70196
rect 71764 70140 71774 70196
rect 69570 70028 69580 70084
rect 69636 70028 74956 70084
rect 75012 70028 75022 70084
rect 3378 69916 3388 69972
rect 3444 69916 4060 69972
rect 4116 69916 4126 69972
rect 0 69860 800 69888
rect 79200 69860 80000 69888
rect 0 69804 2044 69860
rect 2100 69804 2110 69860
rect 75506 69804 75516 69860
rect 75572 69804 80000 69860
rect 0 69776 800 69804
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 79200 69776 80000 69804
rect 68562 69468 68572 69524
rect 68628 69468 72940 69524
rect 72996 69468 73006 69524
rect 66770 69356 66780 69412
rect 66836 69356 74956 69412
rect 75012 69356 75022 69412
rect 1698 69244 1708 69300
rect 1764 69244 2268 69300
rect 2324 69244 4172 69300
rect 4228 69244 4238 69300
rect 69682 69244 69692 69300
rect 69748 69244 70252 69300
rect 70308 69244 71148 69300
rect 71204 69244 71214 69300
rect 76290 69244 76300 69300
rect 76356 69244 77308 69300
rect 77364 69244 77374 69300
rect 0 69188 800 69216
rect 79200 69188 80000 69216
rect 0 69132 2156 69188
rect 2212 69132 2222 69188
rect 3042 69132 3052 69188
rect 3108 69132 69356 69188
rect 69412 69132 69422 69188
rect 74274 69132 74284 69188
rect 74340 69132 74508 69188
rect 74564 69132 80000 69188
rect 0 69104 800 69132
rect 79200 69104 80000 69132
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 2258 68684 2268 68740
rect 2324 68684 3724 68740
rect 3780 68684 3790 68740
rect 76290 68684 76300 68740
rect 76356 68684 76860 68740
rect 76916 68684 76926 68740
rect 3826 68572 3836 68628
rect 3892 68572 8428 68628
rect 0 68516 800 68544
rect 8372 68516 8428 68572
rect 79200 68516 80000 68544
rect 0 68460 3948 68516
rect 4004 68460 4014 68516
rect 8372 68460 67116 68516
rect 67172 68460 67676 68516
rect 67732 68460 67742 68516
rect 77522 68460 77532 68516
rect 77588 68460 80000 68516
rect 0 68432 800 68460
rect 79200 68432 80000 68460
rect 5282 68348 5292 68404
rect 5348 68348 67956 68404
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 67900 68180 67956 68348
rect 69570 68236 69580 68292
rect 69636 68236 75068 68292
rect 75124 68236 75134 68292
rect 67890 68124 67900 68180
rect 67956 68124 68460 68180
rect 68516 68124 68526 68180
rect 64866 67900 64876 67956
rect 64932 67900 74956 67956
rect 75012 67900 75022 67956
rect 0 67844 800 67872
rect 79200 67844 80000 67872
rect 0 67788 1820 67844
rect 1876 67788 1886 67844
rect 76738 67788 76748 67844
rect 76804 67788 80000 67844
rect 0 67760 800 67788
rect 79200 67760 80000 67788
rect 2258 67676 2268 67732
rect 2324 67676 4172 67732
rect 4228 67676 4238 67732
rect 76290 67676 76300 67732
rect 76356 67676 77308 67732
rect 77364 67676 77374 67732
rect 4050 67564 4060 67620
rect 4116 67564 66332 67620
rect 66388 67564 67228 67620
rect 67284 67564 67294 67620
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 1708 67340 2156 67396
rect 2212 67340 2222 67396
rect 0 67172 800 67200
rect 1708 67172 1764 67340
rect 79200 67172 80000 67200
rect 0 67116 1092 67172
rect 1708 67116 1988 67172
rect 67442 67116 67452 67172
rect 67508 67116 75180 67172
rect 75236 67116 75246 67172
rect 76290 67116 76300 67172
rect 76356 67116 76860 67172
rect 76916 67116 76926 67172
rect 77410 67116 77420 67172
rect 77476 67116 80000 67172
rect 0 67088 800 67116
rect 1036 67060 1092 67116
rect 1036 67004 1708 67060
rect 1764 67004 1774 67060
rect 0 66500 800 66528
rect 1932 66500 1988 67116
rect 79200 67088 80000 67116
rect 2146 67004 2156 67060
rect 2212 67004 3724 67060
rect 3780 67004 3790 67060
rect 63522 67004 63532 67060
rect 63588 67004 65884 67060
rect 65940 67004 65950 67060
rect 67666 67004 67676 67060
rect 67732 67004 68124 67060
rect 68180 67004 68190 67060
rect 3826 66892 3836 66948
rect 3892 66892 63420 66948
rect 63476 66892 63980 66948
rect 64036 66892 64046 66948
rect 67554 66892 67564 66948
rect 67620 66892 68236 66948
rect 68292 66892 68302 66948
rect 65772 66780 66108 66836
rect 66164 66780 66174 66836
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 0 66444 1988 66500
rect 65772 66500 65828 66780
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 79200 66500 80000 66528
rect 65772 66444 65884 66500
rect 65940 66444 65950 66500
rect 68338 66444 68348 66500
rect 68404 66444 69356 66500
rect 69412 66444 69422 66500
rect 76962 66444 76972 66500
rect 77028 66444 80000 66500
rect 0 66416 800 66444
rect 79200 66416 80000 66444
rect 66882 66332 66892 66388
rect 66948 66332 67452 66388
rect 67508 66332 67518 66388
rect 65762 66220 65772 66276
rect 65828 66220 67004 66276
rect 67060 66220 67070 66276
rect 67778 66220 67788 66276
rect 67844 66220 68236 66276
rect 68292 66220 68302 66276
rect 3602 66108 3612 66164
rect 3668 66108 63308 66164
rect 63364 66108 63868 66164
rect 63924 66108 63934 66164
rect 2034 65996 2044 66052
rect 2100 65996 3724 66052
rect 3780 65996 3790 66052
rect 63410 65996 63420 66052
rect 63476 65996 65772 66052
rect 65828 65996 65838 66052
rect 76290 65996 76300 66052
rect 76356 65996 77308 66052
rect 77364 65996 77374 66052
rect 0 65828 800 65856
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 79200 65828 80000 65856
rect 0 65772 2268 65828
rect 2324 65772 2334 65828
rect 77410 65772 77420 65828
rect 77476 65772 80000 65828
rect 0 65744 800 65772
rect 79200 65744 80000 65772
rect 62066 65548 62076 65604
rect 62132 65548 65884 65604
rect 65940 65548 65950 65604
rect 68674 65548 68684 65604
rect 68740 65548 69244 65604
rect 69300 65548 69310 65604
rect 76850 65548 76860 65604
rect 76916 65548 76926 65604
rect 3378 65436 3388 65492
rect 3444 65436 4956 65492
rect 5012 65436 5022 65492
rect 65426 65436 65436 65492
rect 65492 65436 66108 65492
rect 66164 65436 66668 65492
rect 66724 65436 66734 65492
rect 67666 65436 67676 65492
rect 67732 65436 68012 65492
rect 68068 65436 68078 65492
rect 1810 65324 1820 65380
rect 1876 65324 3724 65380
rect 3780 65324 3790 65380
rect 4274 65324 4284 65380
rect 4340 65324 61964 65380
rect 62020 65324 62524 65380
rect 62580 65324 62590 65380
rect 68114 65324 68124 65380
rect 68180 65324 68796 65380
rect 68852 65324 68862 65380
rect 0 65156 800 65184
rect 76860 65156 76916 65548
rect 79200 65156 80000 65184
rect 0 65100 2156 65156
rect 2212 65100 2222 65156
rect 3378 65100 3388 65156
rect 3444 65100 4284 65156
rect 4340 65100 4350 65156
rect 66444 65100 67116 65156
rect 67172 65100 75180 65156
rect 75236 65100 75246 65156
rect 76860 65100 80000 65156
rect 0 65072 800 65100
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 66444 65044 66500 65100
rect 79200 65072 80000 65100
rect 66434 64988 66444 65044
rect 66500 64988 66510 65044
rect 68114 64988 68124 65044
rect 68180 64988 74956 65044
rect 75012 64988 75022 65044
rect 65426 64876 65436 64932
rect 65492 64876 65772 64932
rect 65828 64876 65838 64932
rect 64642 64764 64652 64820
rect 64708 64764 72940 64820
rect 72996 64764 73006 64820
rect 1922 64652 1932 64708
rect 1988 64652 4172 64708
rect 4228 64652 4238 64708
rect 63746 64652 63756 64708
rect 63812 64652 64316 64708
rect 64372 64652 75068 64708
rect 75124 64652 75134 64708
rect 3490 64540 3500 64596
rect 3556 64540 60732 64596
rect 60788 64540 61740 64596
rect 61796 64540 61806 64596
rect 65538 64540 65548 64596
rect 65604 64540 66892 64596
rect 66948 64540 66958 64596
rect 67330 64540 67340 64596
rect 67396 64540 68236 64596
rect 68292 64540 68302 64596
rect 76290 64540 76300 64596
rect 76356 64540 77308 64596
rect 77364 64540 77374 64596
rect 0 64484 800 64512
rect 79200 64484 80000 64512
rect 0 64428 2044 64484
rect 2100 64428 2110 64484
rect 61842 64428 61852 64484
rect 61908 64428 65324 64484
rect 65380 64428 65390 64484
rect 74274 64428 74284 64484
rect 74340 64428 74508 64484
rect 74564 64428 80000 64484
rect 0 64400 800 64428
rect 79200 64400 80000 64428
rect 61730 64316 61740 64372
rect 61796 64316 74956 64372
rect 75012 64316 75022 64372
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 2034 64204 2044 64260
rect 2100 64204 3724 64260
rect 3780 64204 3790 64260
rect 65090 64204 65100 64260
rect 65156 64204 66332 64260
rect 66388 64204 66668 64260
rect 66724 64204 66734 64260
rect 59042 64092 59052 64148
rect 59108 64092 62300 64148
rect 62356 64092 62366 64148
rect 65426 64092 65436 64148
rect 65492 64092 65772 64148
rect 65828 64092 65838 64148
rect 67666 64092 67676 64148
rect 67732 64092 68012 64148
rect 68068 64092 69356 64148
rect 69412 64092 69422 64148
rect 61170 63980 61180 64036
rect 61236 63980 63532 64036
rect 63588 63980 63598 64036
rect 4946 63868 4956 63924
rect 5012 63868 61068 63924
rect 61124 63868 61628 63924
rect 61684 63868 61694 63924
rect 62290 63868 62300 63924
rect 62356 63868 65324 63924
rect 65380 63868 65390 63924
rect 66658 63868 66668 63924
rect 66724 63868 67340 63924
rect 67396 63868 67406 63924
rect 77522 63868 77532 63924
rect 77588 63868 77598 63924
rect 0 63812 800 63840
rect 77532 63812 77588 63868
rect 79200 63812 80000 63840
rect 0 63756 3948 63812
rect 4004 63756 4014 63812
rect 5282 63756 5292 63812
rect 5348 63756 59276 63812
rect 59332 63756 59342 63812
rect 62514 63756 62524 63812
rect 62580 63756 63756 63812
rect 63812 63756 63822 63812
rect 76290 63756 76300 63812
rect 76356 63756 76860 63812
rect 76916 63756 76926 63812
rect 77532 63756 80000 63812
rect 0 63728 800 63756
rect 79200 63728 80000 63756
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 59266 63196 59276 63252
rect 59332 63196 59836 63252
rect 59892 63196 59902 63252
rect 0 63140 800 63168
rect 79200 63140 80000 63168
rect 0 63084 1820 63140
rect 1876 63084 1886 63140
rect 76738 63084 76748 63140
rect 76804 63084 80000 63140
rect 0 63056 800 63084
rect 79200 63056 80000 63084
rect 3714 62972 3724 63028
rect 3780 62972 61404 63028
rect 61460 62972 61964 63028
rect 62020 62972 62030 63028
rect 76290 62972 76300 63028
rect 76356 62972 77308 63028
rect 77364 62972 77374 63028
rect 2146 62860 2156 62916
rect 2212 62860 4172 62916
rect 4228 62860 4238 62916
rect 59378 62860 59388 62916
rect 59444 62860 63420 62916
rect 63476 62860 63486 62916
rect 63634 62860 63644 62916
rect 63700 62860 65996 62916
rect 66052 62860 66668 62916
rect 66724 62860 67004 62916
rect 67060 62860 67070 62916
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 1708 62636 1932 62692
rect 1988 62636 1998 62692
rect 0 62468 800 62496
rect 1708 62468 1764 62636
rect 61506 62524 61516 62580
rect 61572 62524 62748 62580
rect 62804 62524 62814 62580
rect 63186 62524 63196 62580
rect 63252 62524 63756 62580
rect 63812 62524 63822 62580
rect 79200 62468 80000 62496
rect 0 62412 1764 62468
rect 1922 62412 1932 62468
rect 1988 62412 3724 62468
rect 3780 62412 3790 62468
rect 68226 62412 68236 62468
rect 68292 62412 68684 62468
rect 68740 62412 68750 62468
rect 77410 62412 77420 62468
rect 77476 62412 80000 62468
rect 0 62384 800 62412
rect 79200 62384 80000 62412
rect 59714 62300 59724 62356
rect 59780 62300 63980 62356
rect 64036 62300 64046 62356
rect 4274 62188 4284 62244
rect 4340 62188 59612 62244
rect 59668 62188 60172 62244
rect 60228 62188 60238 62244
rect 61730 62188 61740 62244
rect 61796 62188 62300 62244
rect 62356 62188 62366 62244
rect 64418 62188 64428 62244
rect 64484 62188 68124 62244
rect 68180 62188 68190 62244
rect 3490 62076 3500 62132
rect 3556 62076 4844 62132
rect 4900 62076 4910 62132
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 0 61796 800 61824
rect 79200 61796 80000 61824
rect 0 61740 2044 61796
rect 2100 61740 2110 61796
rect 63522 61740 63532 61796
rect 63588 61740 63812 61796
rect 77074 61740 77084 61796
rect 77140 61740 80000 61796
rect 0 61712 800 61740
rect 63756 61684 63812 61740
rect 79200 61712 80000 61740
rect 3266 61628 3276 61684
rect 3332 61628 58492 61684
rect 58548 61628 58558 61684
rect 63746 61628 63756 61684
rect 63812 61628 63822 61684
rect 3602 61404 3612 61460
rect 3668 61404 8428 61460
rect 76290 61404 76300 61460
rect 76356 61404 77196 61460
rect 77252 61404 77262 61460
rect 8372 61348 8428 61404
rect 2034 61292 2044 61348
rect 2100 61292 3724 61348
rect 3780 61292 3790 61348
rect 8372 61292 59836 61348
rect 59892 61292 60284 61348
rect 60340 61292 60350 61348
rect 61506 61292 61516 61348
rect 61572 61292 62188 61348
rect 62244 61292 75180 61348
rect 75236 61292 75246 61348
rect 0 61124 800 61152
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 79200 61124 80000 61152
rect 0 61068 2156 61124
rect 2212 61068 2222 61124
rect 77410 61068 77420 61124
rect 77476 61068 80000 61124
rect 0 61040 800 61068
rect 79200 61040 80000 61068
rect 60386 60956 60396 61012
rect 60452 60956 62412 61012
rect 62468 60956 62478 61012
rect 4834 60844 4844 60900
rect 4900 60844 8428 60900
rect 60722 60844 60732 60900
rect 60788 60844 61068 60900
rect 61124 60844 62636 60900
rect 62692 60844 62702 60900
rect 8372 60676 8428 60844
rect 57586 60732 57596 60788
rect 57652 60732 60956 60788
rect 61012 60732 61022 60788
rect 2146 60620 2156 60676
rect 2212 60620 3724 60676
rect 3780 60620 3790 60676
rect 8372 60620 57484 60676
rect 57540 60620 58044 60676
rect 58100 60620 58110 60676
rect 59714 60620 59724 60676
rect 59780 60620 60396 60676
rect 60452 60620 61180 60676
rect 61236 60620 62188 60676
rect 62244 60620 62254 60676
rect 62514 60620 62524 60676
rect 62580 60620 63196 60676
rect 63252 60620 63262 60676
rect 64530 60620 64540 60676
rect 64596 60620 65324 60676
rect 65380 60620 74620 60676
rect 74676 60620 74686 60676
rect 57138 60508 57148 60564
rect 57204 60508 59052 60564
rect 59108 60508 59388 60564
rect 59444 60508 59454 60564
rect 61394 60508 61404 60564
rect 61460 60508 64428 60564
rect 64484 60508 64494 60564
rect 76962 60508 76972 60564
rect 77028 60508 77038 60564
rect 0 60452 800 60480
rect 76972 60452 77028 60508
rect 79200 60452 80000 60480
rect 0 60396 1820 60452
rect 1876 60396 1886 60452
rect 62738 60396 62748 60452
rect 62804 60396 63644 60452
rect 63700 60396 63710 60452
rect 76972 60396 80000 60452
rect 0 60368 800 60396
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 79200 60368 80000 60396
rect 66546 60172 66556 60228
rect 66612 60172 67116 60228
rect 67172 60172 75068 60228
rect 75124 60172 75134 60228
rect 59938 60060 59948 60116
rect 60004 60060 61068 60116
rect 61124 60060 61134 60116
rect 63298 60060 63308 60116
rect 63364 60060 74956 60116
rect 75012 60060 75022 60116
rect 3826 59948 3836 60004
rect 3892 59948 8428 60004
rect 8372 59892 8428 59948
rect 55412 59948 57820 60004
rect 57876 59948 58044 60004
rect 58100 59948 58110 60004
rect 60610 59948 60620 60004
rect 60676 59948 66444 60004
rect 66500 59948 66510 60004
rect 55412 59892 55468 59948
rect 8372 59836 55468 59892
rect 58146 59836 58156 59892
rect 58212 59836 60172 59892
rect 60228 59836 60238 59892
rect 61506 59836 61516 59892
rect 61572 59836 62076 59892
rect 62132 59836 72940 59892
rect 72996 59836 73006 59892
rect 76290 59836 76300 59892
rect 76356 59836 77308 59892
rect 77364 59836 77374 59892
rect 0 59780 800 59808
rect 79200 59780 80000 59808
rect 0 59724 2044 59780
rect 2100 59724 2110 59780
rect 2258 59724 2268 59780
rect 2324 59724 4172 59780
rect 4228 59724 4238 59780
rect 60274 59724 60284 59780
rect 60340 59724 61404 59780
rect 61460 59724 61470 59780
rect 74274 59724 74284 59780
rect 74340 59724 74508 59780
rect 74564 59724 80000 59780
rect 0 59696 800 59724
rect 79200 59696 80000 59724
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 59602 59500 59612 59556
rect 59668 59500 59948 59556
rect 60004 59500 60014 59556
rect 1922 59276 1932 59332
rect 1988 59276 3724 59332
rect 3780 59276 3790 59332
rect 58370 59164 58380 59220
rect 58436 59164 58940 59220
rect 58996 59164 74732 59220
rect 74788 59164 74798 59220
rect 0 59108 800 59136
rect 79200 59108 80000 59136
rect 0 59052 3948 59108
rect 4004 59052 4014 59108
rect 57362 59052 57372 59108
rect 57428 59052 61292 59108
rect 61348 59052 61852 59108
rect 61908 59052 62748 59108
rect 62804 59052 62814 59108
rect 77186 59052 77196 59108
rect 77252 59052 80000 59108
rect 0 59024 800 59052
rect 79200 59024 80000 59052
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 3490 58716 3500 58772
rect 3556 58716 4284 58772
rect 4340 58716 4350 58772
rect 3602 58604 3612 58660
rect 3668 58604 4956 58660
rect 5012 58604 5022 58660
rect 0 58436 800 58464
rect 79200 58436 80000 58464
rect 0 58380 2156 58436
rect 2212 58380 2222 58436
rect 57250 58380 57260 58436
rect 57316 58380 58156 58436
rect 58212 58380 58222 58436
rect 76962 58380 76972 58436
rect 77028 58380 80000 58436
rect 0 58352 800 58380
rect 79200 58352 80000 58380
rect 76290 58268 76300 58324
rect 76356 58268 77308 58324
rect 77364 58268 77374 58324
rect 2034 58156 2044 58212
rect 2100 58156 4172 58212
rect 4228 58156 4238 58212
rect 5282 58156 5292 58212
rect 5348 58156 56700 58212
rect 56756 58156 57148 58212
rect 57204 58156 57214 58212
rect 59266 58156 59276 58212
rect 59332 58156 59836 58212
rect 59892 58156 74844 58212
rect 74900 58156 74910 58212
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 0 57764 800 57792
rect 79200 57764 80000 57792
rect 0 57708 2268 57764
rect 2324 57708 2334 57764
rect 62850 57708 62860 57764
rect 62916 57708 63308 57764
rect 63364 57708 63374 57764
rect 76290 57708 76300 57764
rect 76356 57708 76860 57764
rect 76916 57708 76926 57764
rect 77410 57708 77420 57764
rect 77476 57708 80000 57764
rect 0 57680 800 57708
rect 79200 57680 80000 57708
rect 4274 57596 4284 57652
rect 4340 57596 54572 57652
rect 54628 57596 55132 57652
rect 55188 57596 55198 57652
rect 56130 57596 56140 57652
rect 56196 57596 58044 57652
rect 58100 57596 58110 57652
rect 58482 57596 58492 57652
rect 58548 57596 59164 57652
rect 59220 57596 59230 57652
rect 1922 57484 1932 57540
rect 1988 57484 3724 57540
rect 3780 57484 3790 57540
rect 4946 57484 4956 57540
rect 5012 57484 56028 57540
rect 56084 57484 56588 57540
rect 56644 57484 56654 57540
rect 58034 57372 58044 57428
rect 58100 57372 62748 57428
rect 62804 57372 62814 57428
rect 76738 57260 76748 57316
rect 76804 57260 77588 57316
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 0 57092 800 57120
rect 77532 57092 77588 57260
rect 79200 57092 80000 57120
rect 0 57036 1820 57092
rect 1876 57036 1886 57092
rect 3714 57036 3724 57092
rect 3780 57036 4620 57092
rect 4676 57036 4686 57092
rect 55906 57036 55916 57092
rect 55972 57036 67228 57092
rect 77532 57036 80000 57092
rect 0 57008 800 57036
rect 67172 56980 67228 57036
rect 79200 57008 80000 57036
rect 57810 56924 57820 56980
rect 57876 56924 58268 56980
rect 58324 56924 58334 56980
rect 67172 56924 74956 56980
rect 75012 56924 75022 56980
rect 58044 56868 58100 56924
rect 3826 56812 3836 56868
rect 3892 56812 8428 56868
rect 55234 56812 55244 56868
rect 55300 56812 57596 56868
rect 57652 56812 57662 56868
rect 58034 56812 58044 56868
rect 58100 56812 58110 56868
rect 8372 56756 8428 56812
rect 2258 56700 2268 56756
rect 2324 56700 3724 56756
rect 3780 56700 3790 56756
rect 8372 56700 56140 56756
rect 56196 56700 56588 56756
rect 56644 56700 56654 56756
rect 58930 56700 58940 56756
rect 58996 56700 59500 56756
rect 59556 56700 75180 56756
rect 75236 56700 75246 56756
rect 76290 56700 76300 56756
rect 76356 56700 77308 56756
rect 77364 56700 77374 56756
rect 0 56420 800 56448
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 79200 56420 80000 56448
rect 0 56364 2044 56420
rect 2100 56364 2110 56420
rect 77410 56364 77420 56420
rect 77476 56364 80000 56420
rect 0 56336 800 56364
rect 79200 56336 80000 56364
rect 56690 56252 56700 56308
rect 56756 56252 57820 56308
rect 57876 56252 57886 56308
rect 67172 56252 75068 56308
rect 75124 56252 75134 56308
rect 67172 56196 67228 56252
rect 1810 56140 1820 56196
rect 1876 56140 2268 56196
rect 2324 56140 3724 56196
rect 3780 56140 3790 56196
rect 57820 56140 67228 56196
rect 76290 56140 76300 56196
rect 76356 56140 76860 56196
rect 76916 56140 76926 56196
rect 57820 56084 57876 56140
rect 53218 56028 53228 56084
rect 53284 56028 55580 56084
rect 55636 56028 55646 56084
rect 56690 56028 56700 56084
rect 56756 56028 57820 56084
rect 57876 56028 57886 56084
rect 58258 56028 58268 56084
rect 58324 56028 58828 56084
rect 58884 56028 58894 56084
rect 4610 55916 4620 55972
rect 4676 55916 53116 55972
rect 53172 55916 53676 55972
rect 53732 55916 53742 55972
rect 57698 55916 57708 55972
rect 57764 55916 58604 55972
rect 58660 55916 58670 55972
rect 0 55748 800 55776
rect 79200 55748 80000 55776
rect 0 55692 1932 55748
rect 1988 55692 1998 55748
rect 76962 55692 76972 55748
rect 77028 55692 80000 55748
rect 0 55664 800 55692
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 79200 55664 80000 55692
rect 2044 55468 2156 55524
rect 2212 55468 2222 55524
rect 77298 55468 77308 55524
rect 77364 55468 79268 55524
rect 2044 55188 2100 55468
rect 79212 55412 79268 55468
rect 3266 55356 3276 55412
rect 3332 55356 3948 55412
rect 4004 55356 4014 55412
rect 54450 55356 54460 55412
rect 54516 55356 55020 55412
rect 55076 55356 55692 55412
rect 55748 55356 55758 55412
rect 78988 55356 79268 55412
rect 52322 55244 52332 55300
rect 52388 55244 54236 55300
rect 54292 55244 54572 55300
rect 54628 55244 55748 55300
rect 55906 55244 55916 55300
rect 55972 55244 56588 55300
rect 56644 55244 56654 55300
rect 55692 55188 55748 55244
rect 1036 55132 2100 55188
rect 3490 55132 3500 55188
rect 3556 55132 8428 55188
rect 50754 55132 50764 55188
rect 50820 55132 55468 55188
rect 55524 55132 55534 55188
rect 55692 55132 56364 55188
rect 56420 55132 56924 55188
rect 56980 55132 56990 55188
rect 57250 55132 57260 55188
rect 57316 55132 58044 55188
rect 58100 55132 58110 55188
rect 76290 55132 76300 55188
rect 76356 55132 77308 55188
rect 77364 55132 77374 55188
rect 0 55076 800 55104
rect 1036 55076 1092 55132
rect 8372 55076 8428 55132
rect 78988 55076 79044 55356
rect 79200 55076 80000 55104
rect 0 55020 1092 55076
rect 2034 55020 2044 55076
rect 2100 55020 3724 55076
rect 3780 55020 3790 55076
rect 8372 55020 50652 55076
rect 50708 55020 51212 55076
rect 51268 55020 51278 55076
rect 78988 55020 80000 55076
rect 0 54992 800 55020
rect 79200 54992 80000 55020
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 2146 54684 2156 54740
rect 2212 54684 3724 54740
rect 3780 54684 3790 54740
rect 53890 54684 53900 54740
rect 53956 54684 75068 54740
rect 75124 54684 75134 54740
rect 3378 54572 3388 54628
rect 3444 54572 3454 54628
rect 52210 54572 52220 54628
rect 52276 54572 54908 54628
rect 54964 54572 54974 54628
rect 56690 54572 56700 54628
rect 56756 54572 57372 54628
rect 57428 54572 74844 54628
rect 74900 54572 74910 54628
rect 76290 54572 76300 54628
rect 76356 54572 76860 54628
rect 76916 54572 76926 54628
rect 0 54404 800 54432
rect 3388 54404 3444 54572
rect 3602 54460 3612 54516
rect 3668 54460 51548 54516
rect 51604 54460 52108 54516
rect 52164 54460 52174 54516
rect 79200 54404 80000 54432
rect 0 54348 1820 54404
rect 1876 54348 1886 54404
rect 3388 54348 52780 54404
rect 52836 54348 53340 54404
rect 53396 54348 53406 54404
rect 54786 54348 54796 54404
rect 54852 54348 55244 54404
rect 55300 54348 55310 54404
rect 76962 54348 76972 54404
rect 77028 54348 80000 54404
rect 0 54320 800 54348
rect 79200 54320 80000 54348
rect 55346 54236 55356 54292
rect 55412 54236 55916 54292
rect 55972 54236 55982 54292
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 54674 53900 54684 53956
rect 54740 53900 54964 53956
rect 57586 53900 57596 53956
rect 57652 53900 58044 53956
rect 58100 53900 75068 53956
rect 75124 53900 75134 53956
rect 2034 53788 2044 53844
rect 2100 53788 2110 53844
rect 0 53732 800 53760
rect 2044 53732 2100 53788
rect 0 53676 2100 53732
rect 3378 53676 3388 53732
rect 3444 53676 48188 53732
rect 48244 53676 48254 53732
rect 52882 53676 52892 53732
rect 52948 53676 54684 53732
rect 54740 53676 54750 53732
rect 0 53648 800 53676
rect 54908 53508 54964 53900
rect 61394 53788 61404 53844
rect 61460 53788 74956 53844
rect 75012 53788 75022 53844
rect 77298 53788 77308 53844
rect 77364 53788 77374 53844
rect 77308 53732 77364 53788
rect 79200 53732 80000 53760
rect 77308 53676 80000 53732
rect 79200 53648 80000 53676
rect 76290 53564 76300 53620
rect 76356 53564 77308 53620
rect 77364 53564 77374 53620
rect 2034 53452 2044 53508
rect 2100 53452 3724 53508
rect 3780 53452 3790 53508
rect 54898 53452 54908 53508
rect 54964 53452 55580 53508
rect 55636 53452 55646 53508
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 76850 53228 76860 53284
rect 76916 53228 77140 53284
rect 0 53060 800 53088
rect 77084 53060 77140 53228
rect 79200 53060 80000 53088
rect 0 53004 2156 53060
rect 2212 53004 2222 53060
rect 76290 53004 76300 53060
rect 76356 53004 76860 53060
rect 76916 53004 76926 53060
rect 77084 53004 80000 53060
rect 0 52976 800 53004
rect 79200 52976 80000 53004
rect 3490 52892 3500 52948
rect 3556 52892 47740 52948
rect 47796 52892 48300 52948
rect 48356 52892 48366 52948
rect 50530 52892 50540 52948
rect 50596 52892 53116 52948
rect 53172 52892 53182 52948
rect 1922 52780 1932 52836
rect 1988 52780 3724 52836
rect 3780 52780 3790 52836
rect 3938 52780 3948 52836
rect 4004 52780 50428 52836
rect 50484 52780 50988 52836
rect 51044 52780 51054 52836
rect 52322 52780 52332 52836
rect 52388 52780 53340 52836
rect 53396 52780 53406 52836
rect 53666 52780 53676 52836
rect 53732 52780 54124 52836
rect 54180 52780 75180 52836
rect 75236 52780 75246 52836
rect 53340 52724 53396 52780
rect 3378 52668 3388 52724
rect 3444 52668 49532 52724
rect 49588 52668 49598 52724
rect 53340 52668 54012 52724
rect 54068 52668 54078 52724
rect 56476 52556 57484 52612
rect 57540 52556 57550 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 0 52388 800 52416
rect 56476 52388 56532 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 0 52332 2044 52388
rect 2100 52332 2110 52388
rect 54226 52332 54236 52388
rect 54292 52332 56532 52388
rect 57036 52444 60508 52500
rect 60564 52444 60574 52500
rect 0 52304 800 52332
rect 57036 52276 57092 52444
rect 79200 52388 80000 52416
rect 77298 52332 77308 52388
rect 77364 52332 80000 52388
rect 79200 52304 80000 52332
rect 48290 52220 48300 52276
rect 48356 52220 48860 52276
rect 48916 52220 48926 52276
rect 52658 52220 52668 52276
rect 52724 52220 57092 52276
rect 57372 52220 59276 52276
rect 59332 52220 59342 52276
rect 57372 52164 57428 52220
rect 52546 52108 52556 52164
rect 52612 52108 57428 52164
rect 59378 52108 59388 52164
rect 59444 52108 59948 52164
rect 60004 52108 75068 52164
rect 75124 52108 75134 52164
rect 3378 51996 3388 52052
rect 3444 51996 48972 52052
rect 49028 51996 49038 52052
rect 76290 51996 76300 52052
rect 76356 51996 77308 52052
rect 77364 51996 77374 52052
rect 2034 51884 2044 51940
rect 2100 51884 3724 51940
rect 3780 51884 3790 51940
rect 48402 51884 48412 51940
rect 48468 51884 52220 51940
rect 52276 51884 52286 51940
rect 52770 51884 52780 51940
rect 52836 51884 53676 51940
rect 53732 51884 53742 51940
rect 52098 51772 52108 51828
rect 52164 51772 52444 51828
rect 52500 51772 52510 51828
rect 0 51716 800 51744
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 79200 51716 80000 51744
rect 0 51660 1932 51716
rect 1988 51660 1998 51716
rect 76850 51660 76860 51716
rect 76916 51660 80000 51716
rect 0 51632 800 51660
rect 79200 51632 80000 51660
rect 51874 51548 51884 51604
rect 51940 51548 52892 51604
rect 52948 51548 53340 51604
rect 53396 51548 53406 51604
rect 53666 51548 53676 51604
rect 53732 51548 56252 51604
rect 56308 51548 57036 51604
rect 57092 51548 57102 51604
rect 56588 51492 56644 51548
rect 48514 51436 48524 51492
rect 48580 51436 53788 51492
rect 53844 51436 53854 51492
rect 56578 51436 56588 51492
rect 56644 51436 56654 51492
rect 76290 51436 76300 51492
rect 76356 51436 76860 51492
rect 76916 51436 76926 51492
rect 49634 51324 49644 51380
rect 49700 51324 52108 51380
rect 52164 51324 52174 51380
rect 55682 51324 55692 51380
rect 55748 51324 56252 51380
rect 56308 51324 56924 51380
rect 56980 51324 56990 51380
rect 2146 51212 2156 51268
rect 2212 51212 3724 51268
rect 3780 51212 3790 51268
rect 0 51044 800 51072
rect 79200 51044 80000 51072
rect 0 50988 2044 51044
rect 2100 50988 2110 51044
rect 77298 50988 77308 51044
rect 77364 50988 80000 51044
rect 0 50960 800 50988
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 79200 50960 80000 50988
rect 4946 50652 4956 50708
rect 5012 50652 72156 50708
rect 72212 50652 72604 50708
rect 72660 50652 72670 50708
rect 73490 50652 73500 50708
rect 73556 50652 74060 50708
rect 74116 50652 74126 50708
rect 1922 50540 1932 50596
rect 1988 50540 3724 50596
rect 3780 50540 3790 50596
rect 51762 50540 51772 50596
rect 51828 50540 52332 50596
rect 52388 50540 75180 50596
rect 75236 50540 75246 50596
rect 2146 50428 2156 50484
rect 2212 50428 2222 50484
rect 49522 50428 49532 50484
rect 49588 50428 50652 50484
rect 50708 50428 50718 50484
rect 76290 50428 76300 50484
rect 76356 50428 77308 50484
rect 77364 50428 77374 50484
rect 0 50372 800 50400
rect 2156 50372 2212 50428
rect 79200 50372 80000 50400
rect 0 50316 2212 50372
rect 50418 50316 50428 50372
rect 50484 50316 53452 50372
rect 53508 50316 53518 50372
rect 76850 50316 76860 50372
rect 76916 50316 80000 50372
rect 0 50288 800 50316
rect 79200 50288 80000 50316
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 72706 49980 72716 50036
rect 72772 49980 73836 50036
rect 73892 49980 73902 50036
rect 3602 49868 3612 49924
rect 3668 49868 20188 49924
rect 46722 49868 46732 49924
rect 46788 49868 50428 49924
rect 50484 49868 50494 49924
rect 76290 49868 76300 49924
rect 76356 49868 76860 49924
rect 76916 49868 76926 49924
rect 20132 49812 20188 49868
rect 1820 49756 1932 49812
rect 1988 49756 1998 49812
rect 3490 49756 3500 49812
rect 3556 49756 8428 49812
rect 20132 49756 46620 49812
rect 46676 49756 47180 49812
rect 47236 49756 47246 49812
rect 49410 49756 49420 49812
rect 49476 49756 50092 49812
rect 50148 49756 50652 49812
rect 50708 49756 50988 49812
rect 51044 49756 51054 49812
rect 72594 49756 72604 49812
rect 72660 49756 73612 49812
rect 73668 49756 73678 49812
rect 0 49700 800 49728
rect 1820 49700 1876 49756
rect 8372 49700 8428 49756
rect 79200 49700 80000 49728
rect 0 49644 1876 49700
rect 2034 49644 2044 49700
rect 2100 49644 3724 49700
rect 3780 49644 3790 49700
rect 8372 49644 48188 49700
rect 48244 49644 48748 49700
rect 48804 49644 48814 49700
rect 51538 49644 51548 49700
rect 51604 49644 51996 49700
rect 52052 49644 75068 49700
rect 75124 49644 75134 49700
rect 77298 49644 77308 49700
rect 77364 49644 80000 49700
rect 0 49616 800 49644
rect 79200 49616 80000 49644
rect 55458 49532 55468 49588
rect 55524 49532 56924 49588
rect 56980 49532 56990 49588
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 3378 49196 3388 49252
rect 3444 49196 48076 49252
rect 48132 49196 48412 49252
rect 48468 49196 48478 49252
rect 50642 49196 50652 49252
rect 50708 49196 51212 49252
rect 51268 49196 74844 49252
rect 74900 49196 74910 49252
rect 3266 49084 3276 49140
rect 3332 49084 66668 49140
rect 66724 49084 67116 49140
rect 67172 49084 67182 49140
rect 69458 49084 69468 49140
rect 69524 49084 74956 49140
rect 75012 49084 75022 49140
rect 0 49028 800 49056
rect 79200 49028 80000 49056
rect 0 48972 2044 49028
rect 2100 48972 2110 49028
rect 68562 48972 68572 49028
rect 68628 48972 69356 49028
rect 69412 48972 69422 49028
rect 76850 48972 76860 49028
rect 76916 48972 80000 49028
rect 0 48944 800 48972
rect 79200 48944 80000 48972
rect 68338 48860 68348 48916
rect 68404 48860 70028 48916
rect 70084 48860 72604 48916
rect 72660 48860 72670 48916
rect 76290 48860 76300 48916
rect 76356 48860 77308 48916
rect 77364 48860 77374 48916
rect 1922 48748 1932 48804
rect 1988 48748 4172 48804
rect 4228 48748 4238 48804
rect 48514 48748 48524 48804
rect 48580 48748 49644 48804
rect 49700 48748 49710 48804
rect 67218 48748 67228 48804
rect 67284 48748 68124 48804
rect 68180 48748 68190 48804
rect 67890 48636 67900 48692
rect 67956 48636 68908 48692
rect 68964 48636 73052 48692
rect 73108 48636 74060 48692
rect 74116 48636 74126 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 0 48356 800 48384
rect 79200 48356 80000 48384
rect 0 48300 1932 48356
rect 1988 48300 1998 48356
rect 77298 48300 77308 48356
rect 77364 48300 80000 48356
rect 0 48272 800 48300
rect 79200 48272 80000 48300
rect 48290 48188 48300 48244
rect 48356 48188 49868 48244
rect 49924 48188 49934 48244
rect 4834 48076 4844 48132
rect 4900 48076 5404 48132
rect 5460 48076 47068 48132
rect 47124 48076 47134 48132
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 0 47684 800 47712
rect 79200 47684 80000 47712
rect 0 47628 3724 47684
rect 3780 47628 3790 47684
rect 77858 47628 77868 47684
rect 77924 47628 80000 47684
rect 0 47600 800 47628
rect 79200 47600 80000 47628
rect 47394 47292 47404 47348
rect 47460 47292 47740 47348
rect 47796 47292 48076 47348
rect 48132 47292 48860 47348
rect 48916 47292 48926 47348
rect 49634 47292 49644 47348
rect 49700 47292 50204 47348
rect 50260 47292 75180 47348
rect 75236 47292 75246 47348
rect 48402 47180 48412 47236
rect 48468 47180 76748 47236
rect 76804 47180 77196 47236
rect 77252 47180 77262 47236
rect 75954 47068 75964 47124
rect 76020 47068 76030 47124
rect 0 47012 800 47040
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 75964 47012 76020 47068
rect 79200 47012 80000 47040
rect 0 46956 2044 47012
rect 2100 46956 2110 47012
rect 74274 46956 74284 47012
rect 74340 46956 74956 47012
rect 75012 46956 75022 47012
rect 75964 46956 80000 47012
rect 0 46928 800 46956
rect 79200 46928 80000 46956
rect 74498 46844 74508 46900
rect 74564 46844 74574 46900
rect 74508 46788 74564 46844
rect 3826 46732 3836 46788
rect 3892 46732 46396 46788
rect 46452 46732 46462 46788
rect 47730 46732 47740 46788
rect 47796 46732 74564 46788
rect 3042 46620 3052 46676
rect 3108 46620 3612 46676
rect 3668 46620 3678 46676
rect 45938 46620 45948 46676
rect 46004 46620 46732 46676
rect 46788 46620 47516 46676
rect 47572 46620 48188 46676
rect 48244 46620 48254 46676
rect 0 46340 800 46368
rect 79200 46340 80000 46368
rect 0 46284 1932 46340
rect 1988 46284 1998 46340
rect 76066 46284 76076 46340
rect 76132 46284 80000 46340
rect 0 46256 800 46284
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 79200 46256 80000 46284
rect 46050 45836 46060 45892
rect 46116 45836 46956 45892
rect 47012 45836 47740 45892
rect 47796 45836 47806 45892
rect 47170 45724 47180 45780
rect 47236 45724 74284 45780
rect 74340 45724 74350 45780
rect 0 45668 800 45696
rect 79200 45668 80000 45696
rect 0 45612 2044 45668
rect 2100 45612 2110 45668
rect 3714 45612 3724 45668
rect 3780 45612 45724 45668
rect 45780 45612 45790 45668
rect 46060 45612 74396 45668
rect 74452 45612 74956 45668
rect 75012 45612 75022 45668
rect 75954 45612 75964 45668
rect 76020 45612 80000 45668
rect 0 45584 800 45612
rect 46060 45556 46116 45612
rect 79200 45584 80000 45612
rect 45602 45500 45612 45556
rect 45668 45500 46116 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 3490 45276 3500 45332
rect 3556 45276 44380 45332
rect 44436 45276 44446 45332
rect 74498 45276 74508 45332
rect 74564 45276 74574 45332
rect 74508 45220 74564 45276
rect 3602 45164 3612 45220
rect 3668 45164 46172 45220
rect 46228 45164 46238 45220
rect 47394 45164 47404 45220
rect 47460 45164 74564 45220
rect 43922 45052 43932 45108
rect 43988 45052 44716 45108
rect 44772 45052 45388 45108
rect 45444 45052 45454 45108
rect 46498 45052 46508 45108
rect 46564 45052 47180 45108
rect 47236 45052 47852 45108
rect 47908 45052 47918 45108
rect 0 44996 800 45024
rect 79200 44996 80000 45024
rect 0 44940 1932 44996
rect 1988 44940 1998 44996
rect 3042 44940 3052 44996
rect 3108 44940 3612 44996
rect 3668 44940 43708 44996
rect 43764 44940 43774 44996
rect 76066 44940 76076 44996
rect 76132 44940 80000 44996
rect 0 44912 800 44940
rect 79200 44912 80000 44940
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 45378 44492 45388 44548
rect 45444 44492 46732 44548
rect 46788 44492 46798 44548
rect 0 44324 800 44352
rect 79200 44324 80000 44352
rect 0 44268 2044 44324
rect 2100 44268 2110 44324
rect 75954 44268 75964 44324
rect 76020 44268 80000 44324
rect 0 44240 800 44268
rect 79200 44240 80000 44268
rect 44034 44156 44044 44212
rect 44100 44156 44604 44212
rect 44660 44156 45500 44212
rect 45556 44156 46396 44212
rect 46452 44156 46462 44212
rect 3042 44044 3052 44100
rect 3108 44044 3500 44100
rect 3556 44044 43036 44100
rect 43092 44044 43102 44100
rect 45826 44044 45836 44100
rect 45892 44044 74508 44100
rect 74564 44044 74574 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 44482 43708 44492 43764
rect 44548 43708 74396 43764
rect 74452 43708 74956 43764
rect 75012 43708 75022 43764
rect 76066 43708 76076 43764
rect 76132 43708 76142 43764
rect 0 43652 800 43680
rect 76076 43652 76132 43708
rect 79200 43652 80000 43680
rect 0 43596 1932 43652
rect 1988 43596 1998 43652
rect 76076 43596 80000 43652
rect 0 43568 800 43596
rect 79200 43568 80000 43596
rect 42578 43484 42588 43540
rect 42644 43484 43372 43540
rect 43428 43484 44268 43540
rect 44324 43484 44940 43540
rect 44996 43484 45006 43540
rect 3042 43372 3052 43428
rect 3108 43372 3612 43428
rect 3668 43372 42364 43428
rect 42420 43372 42430 43428
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 0 42980 800 43008
rect 79200 42980 80000 43008
rect 0 42924 1932 42980
rect 1988 42924 1998 42980
rect 76066 42924 76076 42980
rect 76132 42924 80000 42980
rect 0 42896 800 42924
rect 79200 42896 80000 42924
rect 74386 42700 74396 42756
rect 74452 42700 74956 42756
rect 75012 42700 75022 42756
rect 3042 42588 3052 42644
rect 3108 42588 3500 42644
rect 3556 42588 41804 42644
rect 41860 42588 41870 42644
rect 42690 42588 42700 42644
rect 42756 42588 43484 42644
rect 43540 42588 44268 42644
rect 44324 42588 44334 42644
rect 42700 42532 42756 42588
rect 41906 42476 41916 42532
rect 41972 42476 42756 42532
rect 43698 42476 43708 42532
rect 43764 42476 74508 42532
rect 74564 42476 74574 42532
rect 0 42308 800 42336
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 79200 42308 80000 42336
rect 0 42252 1932 42308
rect 1988 42252 1998 42308
rect 76066 42252 76076 42308
rect 76132 42252 80000 42308
rect 0 42224 800 42252
rect 79200 42224 80000 42252
rect 43138 42028 43148 42084
rect 43204 42028 74396 42084
rect 74452 42028 74462 42084
rect 3042 41804 3052 41860
rect 3108 41804 3612 41860
rect 3668 41804 41020 41860
rect 41076 41804 41086 41860
rect 42130 41804 42140 41860
rect 42196 41804 42924 41860
rect 42980 41804 43596 41860
rect 43652 41804 43662 41860
rect 0 41636 800 41664
rect 79200 41636 80000 41664
rect 0 41580 1932 41636
rect 1988 41580 1998 41636
rect 76066 41580 76076 41636
rect 76132 41580 80000 41636
rect 0 41552 800 41580
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 79200 41552 80000 41580
rect 74386 41132 74396 41188
rect 74452 41132 74956 41188
rect 75012 41132 75022 41188
rect 0 40964 800 40992
rect 79200 40964 80000 40992
rect 0 40908 1932 40964
rect 1988 40908 1998 40964
rect 3042 40908 3052 40964
rect 3108 40908 3500 40964
rect 3556 40908 40348 40964
rect 40404 40908 40414 40964
rect 42466 40908 42476 40964
rect 42532 40908 74508 40964
rect 74564 40908 74574 40964
rect 76066 40908 76076 40964
rect 76132 40908 80000 40964
rect 0 40880 800 40908
rect 79200 40880 80000 40908
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 40562 40572 40572 40628
rect 40628 40572 41356 40628
rect 41412 40572 41804 40628
rect 41860 40572 42140 40628
rect 42196 40572 42364 40628
rect 42420 40572 42430 40628
rect 41906 40460 41916 40516
rect 41972 40460 74396 40516
rect 74452 40460 74462 40516
rect 3042 40348 3052 40404
rect 3108 40348 3612 40404
rect 3668 40348 39452 40404
rect 39508 40348 39518 40404
rect 40674 40348 40684 40404
rect 40740 40348 41580 40404
rect 41636 40348 42812 40404
rect 42868 40348 42878 40404
rect 76066 40348 76076 40404
rect 76132 40348 76142 40404
rect 0 40292 800 40320
rect 76076 40292 76132 40348
rect 79200 40292 80000 40320
rect 0 40236 1932 40292
rect 1988 40236 1998 40292
rect 76076 40236 80000 40292
rect 0 40208 800 40236
rect 79200 40208 80000 40236
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 39778 39900 39788 39956
rect 39844 39900 40124 39956
rect 40180 39900 40684 39956
rect 40740 39900 40750 39956
rect 0 39620 800 39648
rect 79200 39620 80000 39648
rect 0 39564 1932 39620
rect 1988 39564 1998 39620
rect 41010 39564 41020 39620
rect 41076 39564 74508 39620
rect 74564 39564 74574 39620
rect 76066 39564 76076 39620
rect 76132 39564 80000 39620
rect 0 39536 800 39564
rect 79200 39536 80000 39564
rect 3042 39452 3052 39508
rect 3108 39452 3612 39508
rect 3668 39452 38892 39508
rect 38948 39452 38958 39508
rect 39218 39452 39228 39508
rect 39284 39452 39788 39508
rect 39844 39452 39854 39508
rect 39228 39396 39284 39452
rect 38434 39340 38444 39396
rect 38500 39340 39004 39396
rect 39060 39340 39284 39396
rect 40114 39340 40124 39396
rect 40180 39340 74508 39396
rect 74564 39340 74956 39396
rect 75012 39340 75022 39396
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 0 38948 800 38976
rect 79200 38948 80000 38976
rect 0 38892 1932 38948
rect 1988 38892 1998 38948
rect 39666 38892 39676 38948
rect 39732 38892 74508 38948
rect 74564 38892 74956 38948
rect 75012 38892 75022 38948
rect 76066 38892 76076 38948
rect 76132 38892 80000 38948
rect 0 38864 800 38892
rect 79200 38864 80000 38892
rect 3042 38780 3052 38836
rect 3108 38780 3612 38836
rect 3668 38780 38332 38836
rect 38388 38780 38398 38836
rect 38658 38780 38668 38836
rect 38724 38780 39452 38836
rect 39508 38780 39518 38836
rect 38668 38724 38724 38780
rect 37874 38668 37884 38724
rect 37940 38668 38724 38724
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 0 38276 800 38304
rect 79200 38276 80000 38304
rect 0 38220 1932 38276
rect 1988 38220 1998 38276
rect 76066 38220 76076 38276
rect 76132 38220 80000 38276
rect 0 38192 800 38220
rect 79200 38192 80000 38220
rect 37986 37884 37996 37940
rect 38052 37884 38892 37940
rect 38948 37884 40012 37940
rect 40068 37884 40078 37940
rect 3042 37772 3052 37828
rect 3108 37772 3612 37828
rect 3668 37772 37660 37828
rect 37716 37772 37726 37828
rect 39106 37772 39116 37828
rect 39172 37772 74508 37828
rect 74564 37772 74956 37828
rect 75012 37772 75022 37828
rect 0 37604 800 37632
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 79200 37604 80000 37632
rect 0 37548 1932 37604
rect 1988 37548 1998 37604
rect 76066 37548 76076 37604
rect 76132 37548 80000 37604
rect 0 37520 800 37548
rect 79200 37520 80000 37548
rect 38434 37324 38444 37380
rect 38500 37324 74508 37380
rect 74564 37324 74956 37380
rect 75012 37324 75022 37380
rect 36530 37212 36540 37268
rect 36596 37212 37324 37268
rect 37380 37212 38108 37268
rect 38164 37212 39340 37268
rect 39396 37212 39406 37268
rect 3042 36988 3052 37044
rect 3108 36988 3612 37044
rect 3668 36988 36988 37044
rect 37044 36988 37054 37044
rect 0 36932 800 36960
rect 79200 36932 80000 36960
rect 0 36876 1932 36932
rect 1988 36876 1998 36932
rect 76066 36876 76076 36932
rect 76132 36876 80000 36932
rect 0 36848 800 36876
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 79200 36848 80000 36876
rect 35858 36316 35868 36372
rect 35924 36316 36540 36372
rect 36596 36316 36606 36372
rect 0 36260 800 36288
rect 79200 36260 80000 36288
rect 0 36204 1932 36260
rect 1988 36204 1998 36260
rect 3042 36204 3052 36260
rect 3108 36204 3612 36260
rect 3668 36204 36316 36260
rect 36372 36204 36382 36260
rect 37874 36204 37884 36260
rect 37940 36204 74508 36260
rect 74564 36204 74956 36260
rect 75012 36204 75022 36260
rect 76066 36204 76076 36260
rect 76132 36204 80000 36260
rect 0 36176 800 36204
rect 79200 36176 80000 36204
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 3042 35756 3052 35812
rect 3108 35756 3612 35812
rect 3668 35756 35644 35812
rect 35700 35756 35710 35812
rect 36978 35756 36988 35812
rect 37044 35756 74508 35812
rect 74564 35756 74956 35812
rect 75012 35756 75022 35812
rect 35970 35644 35980 35700
rect 36036 35644 36652 35700
rect 36708 35644 37884 35700
rect 37940 35644 38332 35700
rect 38388 35644 38398 35700
rect 0 35588 800 35616
rect 79200 35588 80000 35616
rect 0 35532 1932 35588
rect 1988 35532 1998 35588
rect 4834 35532 4844 35588
rect 4900 35532 5404 35588
rect 5460 35532 34300 35588
rect 34356 35532 34366 35588
rect 36530 35532 36540 35588
rect 36596 35532 37436 35588
rect 37492 35532 37502 35588
rect 76066 35532 76076 35588
rect 76132 35532 80000 35588
rect 0 35504 800 35532
rect 79200 35504 80000 35532
rect 35410 35420 35420 35476
rect 35476 35420 36092 35476
rect 36148 35420 37492 35476
rect 37436 35364 37492 35420
rect 37426 35308 37436 35364
rect 37492 35308 37502 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 0 34916 800 34944
rect 79200 34916 80000 34944
rect 0 34860 3724 34916
rect 3780 34860 3790 34916
rect 77858 34860 77868 34916
rect 77924 34860 80000 34916
rect 0 34832 800 34860
rect 79200 34832 80000 34860
rect 33842 34748 33852 34804
rect 33908 34748 34636 34804
rect 34692 34748 35308 34804
rect 35364 34748 35374 34804
rect 36418 34748 36428 34804
rect 36484 34748 74508 34804
rect 74564 34748 74956 34804
rect 75012 34748 75022 34804
rect 3042 34636 3052 34692
rect 3108 34636 4060 34692
rect 4116 34636 34748 34692
rect 34804 34636 34814 34692
rect 35522 34636 35532 34692
rect 35588 34636 76748 34692
rect 76804 34636 77196 34692
rect 77252 34636 77262 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 0 34244 800 34272
rect 79200 34244 80000 34272
rect 0 34188 1932 34244
rect 1988 34188 1998 34244
rect 35074 34188 35084 34244
rect 35140 34188 74508 34244
rect 74564 34188 74956 34244
rect 75012 34188 75022 34244
rect 76066 34188 76076 34244
rect 76132 34188 80000 34244
rect 0 34160 800 34188
rect 79200 34160 80000 34188
rect 34066 34076 34076 34132
rect 34132 34076 34860 34132
rect 34916 34076 36204 34132
rect 36260 34076 36270 34132
rect 3042 33964 3052 34020
rect 3108 33964 3612 34020
rect 3668 33964 33740 34020
rect 33796 33964 33806 34020
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 0 33572 800 33600
rect 79200 33572 80000 33600
rect 0 33516 1932 33572
rect 1988 33516 1998 33572
rect 76066 33516 76076 33572
rect 76132 33516 80000 33572
rect 0 33488 800 33516
rect 79200 33488 80000 33516
rect 32498 33292 32508 33348
rect 32564 33292 33180 33348
rect 33236 33292 34076 33348
rect 34132 33292 34142 33348
rect 3042 33180 3052 33236
rect 3108 33180 3612 33236
rect 3668 33180 32956 33236
rect 33012 33180 33022 33236
rect 34402 33068 34412 33124
rect 34468 33068 74508 33124
rect 74564 33068 74956 33124
rect 75012 33068 75022 33124
rect 0 32900 800 32928
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 79200 32900 80000 32928
rect 0 32844 1932 32900
rect 1988 32844 1998 32900
rect 76066 32844 76076 32900
rect 76132 32844 80000 32900
rect 0 32816 800 32844
rect 79200 32816 80000 32844
rect 33954 32620 33964 32676
rect 34020 32620 74508 32676
rect 74564 32620 74956 32676
rect 75012 32620 75022 32676
rect 31826 32508 31836 32564
rect 31892 32508 32508 32564
rect 32564 32508 33628 32564
rect 33684 32508 33694 32564
rect 3042 32284 3052 32340
rect 3108 32284 3612 32340
rect 3668 32284 32284 32340
rect 32340 32284 32350 32340
rect 0 32228 800 32256
rect 79200 32228 80000 32256
rect 0 32172 1932 32228
rect 1988 32172 1998 32228
rect 76524 32172 80000 32228
rect 0 32144 800 32172
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 76524 31892 76580 32172
rect 79200 32144 80000 32172
rect 76066 31836 76076 31892
rect 76132 31836 76580 31892
rect 31938 31724 31948 31780
rect 32004 31724 32844 31780
rect 32900 31724 33964 31780
rect 34020 31724 34030 31780
rect 31948 31668 32004 31724
rect 31154 31612 31164 31668
rect 31220 31612 32004 31668
rect 0 31556 800 31584
rect 79200 31556 80000 31584
rect 0 31500 1932 31556
rect 1988 31500 1998 31556
rect 3042 31500 3052 31556
rect 3108 31500 3612 31556
rect 3668 31500 31612 31556
rect 31668 31500 31678 31556
rect 33058 31500 33068 31556
rect 33124 31500 74508 31556
rect 74564 31500 74956 31556
rect 75012 31500 75022 31556
rect 76066 31500 76076 31556
rect 76132 31500 80000 31556
rect 0 31472 800 31500
rect 79200 31472 80000 31500
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 3042 31052 3052 31108
rect 3108 31052 3612 31108
rect 3668 31052 30940 31108
rect 30996 31052 31006 31108
rect 32274 31052 32284 31108
rect 32340 31052 74508 31108
rect 74564 31052 74956 31108
rect 75012 31052 75022 31108
rect 31266 30940 31276 30996
rect 31332 30940 32060 30996
rect 32116 30940 32732 30996
rect 32788 30940 32798 30996
rect 0 30884 800 30912
rect 79200 30884 80000 30912
rect 0 30828 1932 30884
rect 1988 30828 1998 30884
rect 4834 30828 4844 30884
rect 4900 30828 5404 30884
rect 5460 30828 29596 30884
rect 29652 30828 29662 30884
rect 76066 30828 76076 30884
rect 76132 30828 80000 30884
rect 0 30800 800 30828
rect 79200 30800 80000 30828
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 77858 30268 77868 30324
rect 77924 30268 77934 30324
rect 0 30212 800 30240
rect 77868 30212 77924 30268
rect 79200 30212 80000 30240
rect 0 30156 3724 30212
rect 3780 30156 3790 30212
rect 77868 30156 80000 30212
rect 0 30128 800 30156
rect 79200 30128 80000 30156
rect 28802 30044 28812 30100
rect 28868 30044 29372 30100
rect 29428 30044 29932 30100
rect 29988 30044 30492 30100
rect 30548 30044 30558 30100
rect 30930 30044 30940 30100
rect 30996 30044 31388 30100
rect 31444 30044 31454 30100
rect 31714 30044 31724 30100
rect 31780 30044 74508 30100
rect 74564 30044 74956 30100
rect 75012 30044 75022 30100
rect 3042 29932 3052 29988
rect 3108 29932 4060 29988
rect 4116 29932 30044 29988
rect 30100 29932 30110 29988
rect 30818 29932 30828 29988
rect 30884 29932 76748 29988
rect 76804 29932 77196 29988
rect 77252 29932 77262 29988
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 0 29540 800 29568
rect 79200 29540 80000 29568
rect 0 29484 1932 29540
rect 1988 29484 1998 29540
rect 30370 29484 30380 29540
rect 30436 29484 74508 29540
rect 74564 29484 74956 29540
rect 75012 29484 75022 29540
rect 76066 29484 76076 29540
rect 76132 29484 80000 29540
rect 0 29456 800 29484
rect 79200 29456 80000 29484
rect 28466 29372 28476 29428
rect 28532 29372 29260 29428
rect 29316 29372 30044 29428
rect 30100 29372 31556 29428
rect 31500 29316 31556 29372
rect 3042 29260 3052 29316
rect 3108 29260 3612 29316
rect 3668 29260 28924 29316
rect 28980 29260 28990 29316
rect 31490 29260 31500 29316
rect 31556 29260 31566 29316
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 0 28868 800 28896
rect 79200 28868 80000 28896
rect 0 28812 1932 28868
rect 1988 28812 1998 28868
rect 76066 28812 76076 28868
rect 76132 28812 80000 28868
rect 0 28784 800 28812
rect 79200 28784 80000 28812
rect 3042 28588 3052 28644
rect 3108 28588 3612 28644
rect 3668 28588 28252 28644
rect 28308 28588 28318 28644
rect 27682 28476 27692 28532
rect 27748 28476 28588 28532
rect 28644 28476 29372 28532
rect 29428 28476 29596 28532
rect 29652 28476 29662 28532
rect 29922 28364 29932 28420
rect 29988 28364 74508 28420
rect 74564 28364 74956 28420
rect 75012 28364 75022 28420
rect 0 28196 800 28224
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 79200 28196 80000 28224
rect 0 28140 1932 28196
rect 1988 28140 1998 28196
rect 76066 28140 76076 28196
rect 76132 28140 80000 28196
rect 0 28112 800 28140
rect 79200 28112 80000 28140
rect 28914 27916 28924 27972
rect 28980 27916 74508 27972
rect 74564 27916 74956 27972
rect 75012 27916 75022 27972
rect 27122 27804 27132 27860
rect 27188 27804 27804 27860
rect 27860 27804 28588 27860
rect 28644 27804 29820 27860
rect 29876 27804 29886 27860
rect 3042 27692 3052 27748
rect 3108 27692 3612 27748
rect 3668 27692 27580 27748
rect 27636 27692 27646 27748
rect 0 27524 800 27552
rect 79200 27524 80000 27552
rect 0 27468 1932 27524
rect 1988 27468 1998 27524
rect 76066 27468 76076 27524
rect 76132 27468 80000 27524
rect 0 27440 800 27468
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 79200 27440 80000 27468
rect 3042 27020 3052 27076
rect 3108 27020 3612 27076
rect 3668 27020 26908 27076
rect 26964 27020 26974 27076
rect 26450 26908 26460 26964
rect 26516 26908 27244 26964
rect 27300 26908 27916 26964
rect 27972 26908 28812 26964
rect 28868 26908 28878 26964
rect 0 26852 800 26880
rect 79200 26852 80000 26880
rect 0 26796 1932 26852
rect 1988 26796 1998 26852
rect 28242 26796 28252 26852
rect 28308 26796 74508 26852
rect 74564 26796 74956 26852
rect 75012 26796 75022 26852
rect 76066 26796 76076 26852
rect 76132 26796 80000 26852
rect 0 26768 800 26796
rect 79200 26768 80000 26796
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 27682 26348 27692 26404
rect 27748 26348 74508 26404
rect 74564 26348 74956 26404
rect 75012 26348 75022 26404
rect 25778 26236 25788 26292
rect 25844 26236 26572 26292
rect 26628 26236 27132 26292
rect 27188 26236 27356 26292
rect 27412 26236 27422 26292
rect 0 26180 800 26208
rect 79200 26180 80000 26208
rect 0 26124 1932 26180
rect 1988 26124 1998 26180
rect 4834 26124 4844 26180
rect 4900 26124 5404 26180
rect 5460 26124 24332 26180
rect 24388 26124 24398 26180
rect 76066 26124 76076 26180
rect 76132 26124 80000 26180
rect 0 26096 800 26124
rect 79200 26096 80000 26124
rect 27570 26012 27580 26068
rect 27636 26012 27646 26068
rect 27580 25956 27636 26012
rect 27346 25900 27356 25956
rect 27412 25900 27636 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 27010 25788 27020 25844
rect 27076 25788 27468 25844
rect 27524 25788 27534 25844
rect 0 25508 800 25536
rect 79200 25508 80000 25536
rect 0 25452 3724 25508
rect 3780 25452 3790 25508
rect 25554 25452 25564 25508
rect 25620 25452 26460 25508
rect 26516 25452 27580 25508
rect 27636 25452 27646 25508
rect 77858 25452 77868 25508
rect 77924 25452 80000 25508
rect 0 25424 800 25452
rect 79200 25424 80000 25452
rect 3042 25340 3052 25396
rect 3108 25340 4060 25396
rect 4116 25340 25228 25396
rect 25284 25340 25294 25396
rect 2930 25228 2940 25284
rect 2996 25228 3612 25284
rect 3668 25228 26236 25284
rect 26292 25228 26302 25284
rect 26674 25228 26684 25284
rect 26740 25228 74508 25284
rect 74564 25228 74956 25284
rect 75012 25228 75022 25284
rect 24658 25116 24668 25172
rect 24724 25116 25004 25172
rect 25060 25116 25900 25172
rect 25956 25116 25966 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 55412 24892 77196 24948
rect 77252 24892 77262 24948
rect 0 24836 800 24864
rect 55412 24836 55468 24892
rect 79200 24836 80000 24864
rect 0 24780 1932 24836
rect 1988 24780 1998 24836
rect 26114 24780 26124 24836
rect 26180 24780 55468 24836
rect 76066 24780 76076 24836
rect 76132 24780 80000 24836
rect 0 24752 800 24780
rect 79200 24752 80000 24780
rect 22754 24668 22764 24724
rect 22820 24668 23100 24724
rect 23156 24668 23996 24724
rect 24052 24668 24062 24724
rect 24882 24668 24892 24724
rect 24948 24668 74508 24724
rect 74564 24668 74956 24724
rect 75012 24668 75022 24724
rect 3042 24444 3052 24500
rect 3108 24444 3612 24500
rect 3668 24444 23660 24500
rect 23716 24444 23726 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 0 24164 800 24192
rect 79200 24164 80000 24192
rect 0 24108 1932 24164
rect 1988 24108 1998 24164
rect 76066 24108 76076 24164
rect 76132 24108 80000 24164
rect 0 24080 800 24108
rect 79200 24080 80000 24108
rect 3042 23660 3052 23716
rect 3108 23660 3612 23716
rect 3668 23660 23660 23716
rect 23716 23660 23726 23716
rect 25666 23660 25676 23716
rect 25732 23660 74508 23716
rect 74564 23660 74956 23716
rect 75012 23660 75022 23716
rect 0 23492 800 23520
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 79200 23492 80000 23520
rect 0 23436 1932 23492
rect 1988 23436 1998 23492
rect 76066 23436 76076 23492
rect 76132 23436 80000 23492
rect 0 23408 800 23436
rect 79200 23408 80000 23436
rect 23874 23212 23884 23268
rect 23940 23212 74508 23268
rect 74564 23212 74956 23268
rect 75012 23212 75022 23268
rect 22754 23100 22764 23156
rect 22820 23100 23100 23156
rect 23156 23100 23660 23156
rect 23716 23100 23726 23156
rect 3042 22988 3052 23044
rect 3108 22988 3612 23044
rect 3668 22988 22428 23044
rect 22484 22988 22494 23044
rect 24322 22876 24332 22932
rect 24388 22876 24398 22932
rect 0 22820 800 22848
rect 24332 22820 24388 22876
rect 79200 22820 80000 22848
rect 0 22764 1932 22820
rect 1988 22764 1998 22820
rect 24332 22764 24556 22820
rect 24612 22764 24622 22820
rect 76066 22764 76076 22820
rect 76132 22764 80000 22820
rect 0 22736 800 22764
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 79200 22736 80000 22764
rect 0 22148 800 22176
rect 79200 22148 80000 22176
rect 0 22092 1932 22148
rect 1988 22092 1998 22148
rect 3042 22092 3052 22148
rect 3108 22092 3612 22148
rect 3668 22092 22092 22148
rect 22148 22092 22158 22148
rect 23314 22092 23324 22148
rect 23380 22092 74508 22148
rect 74564 22092 74956 22148
rect 75012 22092 75022 22148
rect 76066 22092 76076 22148
rect 76132 22092 80000 22148
rect 0 22064 800 22092
rect 79200 22064 80000 22092
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 22642 21756 22652 21812
rect 22708 21756 23100 21812
rect 23156 21756 24220 21812
rect 24276 21756 24286 21812
rect 23986 21644 23996 21700
rect 24052 21644 74508 21700
rect 74564 21644 74956 21700
rect 75012 21644 75022 21700
rect 22082 21532 22092 21588
rect 22148 21532 23100 21588
rect 23156 21532 23660 21588
rect 23716 21532 23884 21588
rect 23940 21532 24444 21588
rect 24500 21532 24510 21588
rect 0 21476 800 21504
rect 79200 21476 80000 21504
rect 0 21420 1932 21476
rect 1988 21420 1998 21476
rect 4834 21420 4844 21476
rect 4900 21420 5404 21476
rect 5460 21420 19628 21476
rect 19684 21420 19694 21476
rect 76066 21420 76076 21476
rect 76132 21420 80000 21476
rect 0 21392 800 21420
rect 79200 21392 80000 21420
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 2930 20860 2940 20916
rect 2996 20860 3612 20916
rect 3668 20860 21756 20916
rect 21812 20860 21822 20916
rect 0 20804 800 20832
rect 79200 20804 80000 20832
rect 0 20748 3724 20804
rect 3780 20748 3790 20804
rect 20962 20748 20972 20804
rect 21028 20748 21868 20804
rect 21924 20748 22764 20804
rect 22820 20748 23212 20804
rect 23268 20748 23278 20804
rect 77858 20748 77868 20804
rect 77924 20748 80000 20804
rect 0 20720 800 20748
rect 79200 20720 80000 20748
rect 3042 20636 3052 20692
rect 3108 20636 4060 20692
rect 4116 20636 21644 20692
rect 21700 20636 21710 20692
rect 23538 20524 23548 20580
rect 23604 20524 74508 20580
rect 74564 20524 74956 20580
rect 75012 20524 75022 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 21186 20188 21196 20244
rect 21252 20188 77196 20244
rect 77252 20188 77262 20244
rect 0 20132 800 20160
rect 79200 20132 80000 20160
rect 0 20076 1932 20132
rect 1988 20076 1998 20132
rect 76066 20076 76076 20132
rect 76132 20076 80000 20132
rect 0 20048 800 20076
rect 79200 20048 80000 20076
rect 19506 19964 19516 20020
rect 19572 19964 20300 20020
rect 20356 19964 20860 20020
rect 20916 19964 21644 20020
rect 21700 19964 21710 20020
rect 3042 19852 3052 19908
rect 3108 19852 3612 19908
rect 3668 19852 19628 19908
rect 19684 19852 19694 19908
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 0 19460 800 19488
rect 79200 19460 80000 19488
rect 0 19404 1932 19460
rect 1988 19404 1998 19460
rect 76066 19404 76076 19460
rect 76132 19404 80000 19460
rect 0 19376 800 19404
rect 79200 19376 80000 19404
rect 21970 19068 21980 19124
rect 22036 19068 74508 19124
rect 74564 19068 74956 19124
rect 75012 19068 75022 19124
rect 18274 18956 18284 19012
rect 18340 18956 18956 19012
rect 19012 18956 19022 19012
rect 20850 18956 20860 19012
rect 20916 18956 74396 19012
rect 74452 18956 74462 19012
rect 3042 18844 3052 18900
rect 3108 18844 3612 18900
rect 3668 18844 18732 18900
rect 18788 18844 18798 18900
rect 0 18788 800 18816
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 79200 18788 80000 18816
rect 0 18732 1932 18788
rect 1988 18732 1998 18788
rect 76066 18732 76076 18788
rect 76132 18732 80000 18788
rect 0 18704 800 18732
rect 79200 18704 80000 18732
rect 20850 18620 20860 18676
rect 20916 18620 21532 18676
rect 21588 18620 21598 18676
rect 54898 18508 54908 18564
rect 54964 18508 55580 18564
rect 55636 18508 55646 18564
rect 20178 18396 20188 18452
rect 20244 18396 20524 18452
rect 20580 18396 20590 18452
rect 21074 18396 21084 18452
rect 21140 18396 74508 18452
rect 74564 18396 74956 18452
rect 75012 18396 75022 18452
rect 3042 18284 3052 18340
rect 3108 18284 3612 18340
rect 3668 18284 18620 18340
rect 18676 18284 18686 18340
rect 55122 18284 55132 18340
rect 55188 18284 55804 18340
rect 55860 18284 55870 18340
rect 0 18116 800 18144
rect 79200 18116 80000 18144
rect 0 18060 1932 18116
rect 1988 18060 1998 18116
rect 76066 18060 76076 18116
rect 76132 18060 80000 18116
rect 0 18032 800 18060
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 79200 18032 80000 18060
rect 20290 17612 20300 17668
rect 20356 17612 21532 17668
rect 21588 17612 21598 17668
rect 54114 17612 54124 17668
rect 54180 17612 55580 17668
rect 55636 17612 56140 17668
rect 56196 17612 56700 17668
rect 56756 17612 56766 17668
rect 18834 17500 18844 17556
rect 18900 17500 74508 17556
rect 74564 17500 74956 17556
rect 75012 17500 75022 17556
rect 0 17444 800 17472
rect 79200 17444 80000 17472
rect 0 17388 1932 17444
rect 1988 17388 1998 17444
rect 20850 17388 20860 17444
rect 20916 17388 26012 17444
rect 26068 17388 26078 17444
rect 55346 17388 55356 17444
rect 55412 17388 56028 17444
rect 56084 17388 56094 17444
rect 76066 17388 76076 17444
rect 76132 17388 80000 17444
rect 0 17360 800 17388
rect 79200 17360 80000 17388
rect 3042 17276 3052 17332
rect 3108 17276 3612 17332
rect 3668 17276 17612 17332
rect 17668 17276 17678 17332
rect 20178 17276 20188 17332
rect 20244 17276 20254 17332
rect 25218 17276 25228 17332
rect 25284 17276 26124 17332
rect 26180 17276 26572 17332
rect 26628 17276 26638 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 20188 17220 20244 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 20188 17164 20860 17220
rect 20916 17164 21980 17220
rect 22036 17164 22428 17220
rect 22484 17164 22494 17220
rect 23090 17164 23100 17220
rect 23156 17164 24444 17220
rect 24500 17164 25676 17220
rect 25732 17164 25742 17220
rect 18722 17052 18732 17108
rect 18788 17052 19292 17108
rect 19348 17052 21084 17108
rect 21140 17052 21150 17108
rect 23314 17052 23324 17108
rect 23380 17052 53676 17108
rect 53732 17052 55132 17108
rect 55188 17052 55198 17108
rect 3042 16940 3052 16996
rect 3108 16940 3612 16996
rect 3668 16940 16604 16996
rect 16660 16940 16670 16996
rect 18498 16940 18508 16996
rect 18564 16940 74508 16996
rect 74564 16940 74956 16996
rect 75012 16940 75022 16996
rect 4834 16828 4844 16884
rect 4900 16828 5404 16884
rect 5460 16828 15820 16884
rect 15876 16828 15886 16884
rect 16034 16828 16044 16884
rect 16100 16828 16380 16884
rect 16436 16828 16716 16884
rect 16772 16828 18732 16884
rect 18788 16828 19180 16884
rect 19236 16828 20412 16884
rect 20468 16828 20478 16884
rect 23650 16828 23660 16884
rect 23716 16828 24220 16884
rect 24276 16828 24286 16884
rect 24882 16828 24892 16884
rect 24948 16828 25900 16884
rect 25956 16828 25966 16884
rect 26674 16828 26684 16884
rect 26740 16828 54572 16884
rect 54628 16828 55356 16884
rect 55412 16828 55422 16884
rect 0 16772 800 16800
rect 79200 16772 80000 16800
rect 0 16716 1932 16772
rect 1988 16716 1998 16772
rect 20738 16716 20748 16772
rect 20804 16716 21196 16772
rect 21252 16716 22316 16772
rect 22372 16716 23212 16772
rect 23268 16716 23278 16772
rect 76066 16716 76076 16772
rect 76132 16716 80000 16772
rect 0 16688 800 16716
rect 79200 16688 80000 16716
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 19506 16156 19516 16212
rect 19572 16156 31948 16212
rect 0 16100 800 16128
rect 31892 16100 31948 16156
rect 79200 16100 80000 16128
rect 0 16044 3724 16100
rect 3780 16044 3790 16100
rect 18834 16044 18844 16100
rect 18900 16044 22652 16100
rect 22708 16044 22718 16100
rect 31892 16044 74508 16100
rect 74564 16044 74956 16100
rect 75012 16044 75022 16100
rect 77858 16044 77868 16100
rect 77924 16044 80000 16100
rect 0 16016 800 16044
rect 79200 16016 80000 16044
rect 19404 15932 20188 15988
rect 20244 15932 20254 15988
rect 19404 15876 19460 15932
rect 3042 15820 3052 15876
rect 3108 15820 4060 15876
rect 4116 15820 15708 15876
rect 15764 15820 15774 15876
rect 18498 15820 18508 15876
rect 18564 15820 19404 15876
rect 19460 15820 19470 15876
rect 19730 15820 19740 15876
rect 19796 15820 76748 15876
rect 76804 15820 77196 15876
rect 77252 15820 77262 15876
rect 22642 15708 22652 15764
rect 22708 15708 23436 15764
rect 23492 15708 24332 15764
rect 24388 15708 24398 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 0 15428 800 15456
rect 79200 15428 80000 15456
rect 0 15372 1932 15428
rect 1988 15372 1998 15428
rect 18274 15372 18284 15428
rect 18340 15372 19124 15428
rect 56354 15372 56364 15428
rect 56420 15372 74508 15428
rect 74564 15372 74956 15428
rect 75012 15372 75022 15428
rect 76066 15372 76076 15428
rect 76132 15372 80000 15428
rect 0 15344 800 15372
rect 19068 15316 19124 15372
rect 79200 15344 80000 15372
rect 16370 15260 16380 15316
rect 16436 15260 17052 15316
rect 17108 15260 18508 15316
rect 18564 15260 18574 15316
rect 19058 15260 19068 15316
rect 19124 15260 19134 15316
rect 55412 15260 56028 15316
rect 56084 15260 56094 15316
rect 3042 15148 3052 15204
rect 3108 15148 3612 15204
rect 3668 15148 14700 15204
rect 14756 15148 14766 15204
rect 15026 15148 15036 15204
rect 15092 15148 15484 15204
rect 15540 15148 19628 15204
rect 19684 15148 54124 15204
rect 54180 15148 55356 15204
rect 55412 15148 55468 15260
rect 17042 15036 17052 15092
rect 17108 15036 17724 15092
rect 17780 15036 17790 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 0 14756 800 14784
rect 79200 14756 80000 14784
rect 0 14700 1932 14756
rect 1988 14700 1998 14756
rect 76066 14700 76076 14756
rect 76132 14700 80000 14756
rect 0 14672 800 14700
rect 79200 14672 80000 14700
rect 55412 14476 56140 14532
rect 56196 14476 56812 14532
rect 56868 14476 56878 14532
rect 55412 14308 55468 14476
rect 3042 14252 3052 14308
rect 3108 14252 3612 14308
rect 3668 14252 14028 14308
rect 14084 14252 14094 14308
rect 14354 14252 14364 14308
rect 14420 14252 14812 14308
rect 14868 14252 16940 14308
rect 16996 14252 53676 14308
rect 53732 14252 55132 14308
rect 55188 14252 55468 14308
rect 56354 14252 56364 14308
rect 56420 14252 74508 14308
rect 74564 14252 74956 14308
rect 75012 14252 75022 14308
rect 0 14084 800 14112
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 79200 14084 80000 14112
rect 0 14028 1932 14084
rect 1988 14028 1998 14084
rect 76066 14028 76076 14084
rect 76132 14028 80000 14084
rect 0 14000 800 14028
rect 79200 14000 80000 14028
rect 55682 13804 55692 13860
rect 55748 13804 74508 13860
rect 74564 13804 74956 13860
rect 75012 13804 75022 13860
rect 13682 13692 13692 13748
rect 13748 13692 14140 13748
rect 14196 13692 16828 13748
rect 16884 13692 54572 13748
rect 54628 13692 55020 13748
rect 55076 13692 55356 13748
rect 55412 13692 55422 13748
rect 57810 13692 57820 13748
rect 57876 13692 74396 13748
rect 74452 13692 74462 13748
rect 3042 13580 3052 13636
rect 3108 13580 3612 13636
rect 3668 13580 13356 13636
rect 13412 13580 13422 13636
rect 12002 13468 12012 13524
rect 12068 13468 12796 13524
rect 12852 13468 14028 13524
rect 14084 13468 56700 13524
rect 56756 13468 57484 13524
rect 57540 13468 57550 13524
rect 0 13412 800 13440
rect 79200 13412 80000 13440
rect 0 13356 1932 13412
rect 1988 13356 1998 13412
rect 24322 13356 24332 13412
rect 24388 13356 25340 13412
rect 25396 13356 25406 13412
rect 76066 13356 76076 13412
rect 76132 13356 80000 13412
rect 0 13328 800 13356
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 79200 13328 80000 13356
rect 0 12740 800 12768
rect 79200 12740 80000 12768
rect 0 12684 1932 12740
rect 1988 12684 1998 12740
rect 3042 12684 3052 12740
rect 3108 12684 3612 12740
rect 3668 12684 12460 12740
rect 12516 12684 12526 12740
rect 76066 12684 76076 12740
rect 76132 12684 80000 12740
rect 0 12656 800 12684
rect 79200 12656 80000 12684
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 3042 12236 3052 12292
rect 3108 12236 3612 12292
rect 3668 12236 12236 12292
rect 12292 12236 12302 12292
rect 13458 12236 13468 12292
rect 13524 12236 74508 12292
rect 74564 12236 74956 12292
rect 75012 12236 75022 12292
rect 12562 12124 12572 12180
rect 12628 12124 12908 12180
rect 12964 12124 13244 12180
rect 13300 12124 13916 12180
rect 13972 12124 13982 12180
rect 0 12068 800 12096
rect 79200 12068 80000 12096
rect 0 12012 1932 12068
rect 1988 12012 1998 12068
rect 76066 12012 76076 12068
rect 76132 12012 80000 12068
rect 0 11984 800 12012
rect 79200 11984 80000 12012
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 3042 11452 3052 11508
rect 3108 11452 4060 11508
rect 4116 11452 11340 11508
rect 11396 11452 11406 11508
rect 0 11396 800 11424
rect 79200 11396 80000 11424
rect 0 11340 3724 11396
rect 3780 11340 3790 11396
rect 11778 11340 11788 11396
rect 11844 11340 12572 11396
rect 12628 11340 13580 11396
rect 13636 11340 13646 11396
rect 77858 11340 77868 11396
rect 77924 11340 80000 11396
rect 0 11312 800 11340
rect 79200 11312 80000 11340
rect 4834 11228 4844 11284
rect 4900 11228 10668 11284
rect 10724 11228 10734 11284
rect 12786 11228 12796 11284
rect 12852 11228 74508 11284
rect 74564 11228 74956 11284
rect 75012 11228 75022 11284
rect 11890 11116 11900 11172
rect 11956 11116 76748 11172
rect 76804 11116 77196 11172
rect 77252 11116 77262 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 0 10724 800 10752
rect 79200 10724 80000 10752
rect 0 10668 1932 10724
rect 1988 10668 1998 10724
rect 3042 10668 3052 10724
rect 3108 10668 10108 10724
rect 10164 10668 10174 10724
rect 11442 10668 11452 10724
rect 11508 10668 74508 10724
rect 74564 10668 74956 10724
rect 75012 10668 75022 10724
rect 76066 10668 76076 10724
rect 76132 10668 80000 10724
rect 0 10640 800 10668
rect 79200 10640 80000 10668
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 0 10052 800 10080
rect 79200 10052 80000 10080
rect 0 9996 1932 10052
rect 1988 9996 1998 10052
rect 76066 9996 76076 10052
rect 76132 9996 80000 10052
rect 0 9968 800 9996
rect 79200 9968 80000 9996
rect 3042 9660 3052 9716
rect 3108 9660 9436 9716
rect 9492 9660 9502 9716
rect 9650 9660 9660 9716
rect 9716 9660 10556 9716
rect 10612 9660 10622 9716
rect 10882 9548 10892 9604
rect 10948 9548 74508 9604
rect 74564 9548 74956 9604
rect 75012 9548 75022 9604
rect 0 9380 800 9408
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 79200 9380 80000 9408
rect 0 9324 1932 9380
rect 1988 9324 1998 9380
rect 76066 9324 76076 9380
rect 76132 9324 80000 9380
rect 0 9296 800 9324
rect 79200 9296 80000 9324
rect 3042 9100 3052 9156
rect 3108 9100 8652 9156
rect 8708 9100 8718 9156
rect 10210 9100 10220 9156
rect 10276 9100 74508 9156
rect 74564 9100 74956 9156
rect 75012 9100 75022 9156
rect 8978 8988 8988 9044
rect 9044 8988 9884 9044
rect 9940 8988 9950 9044
rect 0 8708 800 8736
rect 79200 8708 80000 8736
rect 0 8652 1932 8708
rect 1988 8652 1998 8708
rect 76524 8652 80000 8708
rect 0 8624 800 8652
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 76524 8372 76580 8652
rect 79200 8624 80000 8652
rect 76066 8316 76076 8372
rect 76132 8316 76580 8372
rect 3042 8092 3052 8148
rect 3108 8092 8092 8148
rect 8148 8092 8158 8148
rect 8418 8092 8428 8148
rect 8484 8092 8988 8148
rect 9044 8092 9054 8148
rect 0 8036 800 8064
rect 79200 8036 80000 8064
rect 0 7980 1932 8036
rect 1988 7980 1998 8036
rect 9426 7980 9436 8036
rect 9492 7980 74508 8036
rect 74564 7980 74956 8036
rect 75012 7980 75022 8036
rect 76066 7980 76076 8036
rect 76132 7980 80000 8036
rect 0 7952 800 7980
rect 79200 7952 80000 7980
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 3042 7532 3052 7588
rect 3108 7532 7420 7588
rect 7476 7532 7486 7588
rect 8754 7532 8764 7588
rect 8820 7532 74508 7588
rect 74564 7532 74956 7588
rect 75012 7532 75022 7588
rect 7634 7420 7644 7476
rect 7700 7420 8428 7476
rect 8484 7420 8494 7476
rect 0 7364 800 7392
rect 79200 7364 80000 7392
rect 0 7308 1932 7364
rect 1988 7308 1998 7364
rect 76066 7308 76076 7364
rect 76132 7308 80000 7364
rect 0 7280 800 7308
rect 79200 7280 80000 7308
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 3042 6748 3052 6804
rect 3108 6748 6524 6804
rect 6580 6748 6590 6804
rect 6850 6748 6860 6804
rect 6916 6748 7868 6804
rect 7924 6748 7934 6804
rect 77858 6748 77868 6804
rect 77924 6748 77934 6804
rect 0 6692 800 6720
rect 77868 6692 77924 6748
rect 79200 6692 80000 6720
rect 0 6636 3724 6692
rect 3780 6636 3790 6692
rect 5730 6636 5740 6692
rect 5796 6636 6300 6692
rect 6356 6636 6972 6692
rect 7028 6636 7038 6692
rect 7298 6636 7308 6692
rect 7364 6636 55468 6692
rect 57922 6636 57932 6692
rect 57988 6636 60284 6692
rect 60340 6636 60350 6692
rect 67666 6636 67676 6692
rect 67732 6636 68684 6692
rect 68740 6636 69356 6692
rect 69412 6636 69422 6692
rect 77868 6636 80000 6692
rect 0 6608 800 6636
rect 55412 6580 55468 6636
rect 79200 6608 80000 6636
rect 4834 6524 4844 6580
rect 4900 6524 6076 6580
rect 6132 6524 6142 6580
rect 26562 6524 26572 6580
rect 26628 6524 28028 6580
rect 28084 6524 28094 6580
rect 52434 6524 52444 6580
rect 52500 6524 54236 6580
rect 54292 6524 54302 6580
rect 55412 6524 76748 6580
rect 76804 6524 77196 6580
rect 77252 6524 77262 6580
rect 52994 6412 53004 6468
rect 53060 6412 55804 6468
rect 55860 6412 55870 6468
rect 58034 6412 58044 6468
rect 58100 6412 59164 6468
rect 59220 6412 59230 6468
rect 66770 6412 66780 6468
rect 66836 6412 67116 6468
rect 67172 6412 67182 6468
rect 52770 6300 52780 6356
rect 52836 6300 54460 6356
rect 54516 6300 55356 6356
rect 55412 6300 55422 6356
rect 56700 6300 57372 6356
rect 57428 6300 57438 6356
rect 57698 6300 57708 6356
rect 57764 6300 59612 6356
rect 59668 6300 59678 6356
rect 60050 6300 60060 6356
rect 60116 6300 62076 6356
rect 62132 6300 62142 6356
rect 63522 6300 63532 6356
rect 63588 6300 65772 6356
rect 65828 6300 65838 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 56700 6244 56756 6300
rect 51986 6188 51996 6244
rect 52052 6188 53004 6244
rect 53060 6188 53340 6244
rect 53396 6188 53406 6244
rect 54338 6188 54348 6244
rect 54404 6188 56756 6244
rect 56914 6188 56924 6244
rect 56980 6188 58156 6244
rect 58212 6188 58222 6244
rect 59714 6188 59724 6244
rect 59780 6188 61068 6244
rect 61124 6188 61516 6244
rect 61572 6188 61582 6244
rect 62850 6188 62860 6244
rect 62916 6188 64204 6244
rect 64260 6188 64270 6244
rect 65426 6188 65436 6244
rect 65492 6188 66332 6244
rect 66388 6188 66398 6244
rect 66770 6188 66780 6244
rect 66836 6188 67004 6244
rect 67060 6188 67340 6244
rect 67396 6188 67406 6244
rect 8194 6076 8204 6132
rect 8260 6076 74508 6132
rect 74564 6076 74956 6132
rect 75012 6076 75022 6132
rect 0 6020 800 6048
rect 79200 6020 80000 6048
rect 0 5964 1932 6020
rect 1988 5964 1998 6020
rect 3042 5964 3052 6020
rect 3108 5964 4620 6020
rect 4676 5964 4686 6020
rect 7298 5964 7308 6020
rect 7364 5964 8652 6020
rect 8708 5964 8718 6020
rect 19394 5964 19404 6020
rect 19460 5964 20300 6020
rect 20356 5964 20366 6020
rect 27682 5964 27692 6020
rect 27748 5964 28700 6020
rect 28756 5964 28766 6020
rect 29586 5964 29596 6020
rect 29652 5964 30380 6020
rect 30436 5964 31052 6020
rect 31108 5964 31118 6020
rect 34850 5964 34860 6020
rect 34916 5964 35196 6020
rect 35252 5964 35262 6020
rect 46722 5964 46732 6020
rect 46788 5964 47292 6020
rect 47348 5964 47358 6020
rect 53890 5964 53900 6020
rect 53956 5964 56364 6020
rect 56420 5964 56430 6020
rect 76066 5964 76076 6020
rect 76132 5964 80000 6020
rect 0 5936 800 5964
rect 28700 5908 28756 5964
rect 79200 5936 80000 5964
rect 16034 5852 16044 5908
rect 16100 5852 18396 5908
rect 18452 5852 18462 5908
rect 28700 5852 29484 5908
rect 29540 5852 29550 5908
rect 49970 5852 49980 5908
rect 50036 5852 50540 5908
rect 50596 5852 51212 5908
rect 51268 5852 51278 5908
rect 68786 5852 68796 5908
rect 68852 5852 70140 5908
rect 70196 5852 70812 5908
rect 70868 5852 70878 5908
rect 11218 5740 11228 5796
rect 11284 5740 11900 5796
rect 11956 5740 11966 5796
rect 12674 5740 12684 5796
rect 12740 5740 13916 5796
rect 13972 5740 13982 5796
rect 16706 5740 16716 5796
rect 16772 5740 17052 5796
rect 17108 5740 17118 5796
rect 38098 5740 38108 5796
rect 38164 5740 38780 5796
rect 38836 5740 38846 5796
rect 48962 5740 48972 5796
rect 49028 5740 49644 5796
rect 49700 5740 49710 5796
rect 67218 5740 67228 5796
rect 67284 5740 68012 5796
rect 68068 5740 68078 5796
rect 16594 5628 16604 5684
rect 16660 5628 17276 5684
rect 17332 5628 17948 5684
rect 18004 5628 18014 5684
rect 67778 5516 67788 5572
rect 67844 5516 69356 5572
rect 69412 5516 69422 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 31602 5404 31612 5460
rect 31668 5404 32396 5460
rect 32452 5404 33516 5460
rect 33572 5404 33582 5460
rect 67172 5404 68124 5460
rect 68180 5404 68190 5460
rect 0 5348 800 5376
rect 67172 5348 67228 5404
rect 79200 5348 80000 5376
rect 0 5292 1932 5348
rect 1988 5292 1998 5348
rect 50754 5292 50764 5348
rect 50820 5292 51660 5348
rect 51716 5292 67228 5348
rect 77858 5292 77868 5348
rect 77924 5292 80000 5348
rect 0 5264 800 5292
rect 79200 5264 80000 5292
rect 4610 5180 4620 5236
rect 4676 5180 5516 5236
rect 5572 5180 5582 5236
rect 16706 5180 16716 5236
rect 16772 5180 17164 5236
rect 17220 5180 17230 5236
rect 19506 5180 19516 5236
rect 19572 5180 21980 5236
rect 22036 5180 22046 5236
rect 38882 5180 38892 5236
rect 38948 5180 39676 5236
rect 39732 5180 39742 5236
rect 42914 5180 42924 5236
rect 42980 5180 43708 5236
rect 43764 5180 43774 5236
rect 47730 5180 47740 5236
rect 47796 5180 48748 5236
rect 48804 5180 48814 5236
rect 50978 5180 50988 5236
rect 51044 5180 51996 5236
rect 52052 5180 52062 5236
rect 55010 5180 55020 5236
rect 55076 5180 55916 5236
rect 55972 5180 55982 5236
rect 60946 5180 60956 5236
rect 61012 5180 62076 5236
rect 62132 5180 62142 5236
rect 66546 5180 66556 5236
rect 66612 5180 67788 5236
rect 67844 5180 67854 5236
rect 68002 5180 68012 5236
rect 68068 5180 70140 5236
rect 70196 5180 70206 5236
rect 20962 5068 20972 5124
rect 21028 5068 21644 5124
rect 21700 5068 21710 5124
rect 35634 5068 35644 5124
rect 35700 5068 36316 5124
rect 36372 5068 37436 5124
rect 37492 5068 37502 5124
rect 48290 5068 48300 5124
rect 48356 5068 49644 5124
rect 49700 5068 49710 5124
rect 68450 5068 68460 5124
rect 68516 5068 69244 5124
rect 69300 5068 69310 5124
rect 5058 4956 5068 5012
rect 5124 4956 6412 5012
rect 6468 4956 6478 5012
rect 10434 4956 10444 5012
rect 10500 4956 11116 5012
rect 11172 4956 11182 5012
rect 11330 4956 11340 5012
rect 11396 4956 12460 5012
rect 12516 4956 12526 5012
rect 13458 4956 13468 5012
rect 13524 4956 13692 5012
rect 13748 4956 13758 5012
rect 15810 4956 15820 5012
rect 15876 4956 17388 5012
rect 17444 4956 17454 5012
rect 17826 4956 17836 5012
rect 17892 4956 18732 5012
rect 18788 4956 18798 5012
rect 28354 4956 28364 5012
rect 28420 4956 29932 5012
rect 29988 4956 29998 5012
rect 41570 4956 41580 5012
rect 41636 4956 42812 5012
rect 42868 4956 42878 5012
rect 44818 4956 44828 5012
rect 44884 4956 45612 5012
rect 45668 4956 45678 5012
rect 52994 4956 53004 5012
rect 53060 4956 53564 5012
rect 53620 4956 53630 5012
rect 73490 4956 73500 5012
rect 73556 4956 75068 5012
rect 75124 4956 75134 5012
rect 4946 4844 4956 4900
rect 5012 4844 76524 4900
rect 76580 4844 76590 4900
rect 4162 4732 4172 4788
rect 4228 4732 5292 4788
rect 5348 4732 6860 4788
rect 6916 4732 6926 4788
rect 12450 4732 12460 4788
rect 12516 4732 14476 4788
rect 14532 4732 14542 4788
rect 37986 4732 37996 4788
rect 38052 4732 38220 4788
rect 38276 4732 38668 4788
rect 38724 4732 38734 4788
rect 40226 4732 40236 4788
rect 40292 4732 41468 4788
rect 41524 4732 41534 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 6738 4620 6748 4676
rect 6804 4620 8428 4676
rect 8372 4564 8428 4620
rect 3042 4508 3052 4564
rect 3108 4508 4620 4564
rect 4676 4508 4686 4564
rect 8372 4508 74508 4564
rect 74564 4508 74574 4564
rect 19842 4396 19852 4452
rect 19908 4396 21308 4452
rect 21364 4396 21374 4452
rect 29810 4396 29820 4452
rect 29876 4396 30828 4452
rect 30884 4396 30894 4452
rect 63746 4396 63756 4452
rect 63812 4396 67452 4452
rect 67508 4396 67518 4452
rect 72482 4396 72492 4452
rect 72548 4396 73388 4452
rect 73444 4396 74396 4452
rect 74452 4396 74462 4452
rect 8372 4284 9660 4340
rect 9716 4284 9726 4340
rect 24770 4284 24780 4340
rect 24836 4284 26012 4340
rect 26068 4284 26078 4340
rect 32274 4284 32284 4340
rect 32340 4284 33516 4340
rect 33572 4284 33582 4340
rect 49858 4284 49868 4340
rect 49924 4284 51548 4340
rect 51604 4284 51614 4340
rect 63186 4284 63196 4340
rect 63252 4284 63868 4340
rect 63924 4284 64540 4340
rect 64596 4284 64606 4340
rect 66882 4284 66892 4340
rect 66948 4284 68236 4340
rect 68292 4284 68908 4340
rect 68964 4284 68974 4340
rect 8082 4172 8092 4228
rect 8148 4172 8316 4228
rect 8372 4172 8428 4284
rect 24098 4172 24108 4228
rect 24164 4172 25564 4228
rect 25620 4172 25630 4228
rect 26114 4172 26124 4228
rect 26180 4172 26796 4228
rect 26852 4172 26862 4228
rect 32834 4172 32844 4228
rect 32900 4172 33964 4228
rect 34020 4172 34030 4228
rect 44370 4172 44380 4228
rect 44436 4172 45388 4228
rect 45444 4172 45724 4228
rect 45780 4172 45790 4228
rect 46274 4172 46284 4228
rect 46340 4172 47516 4228
rect 47572 4172 47582 4228
rect 49634 4172 49644 4228
rect 49700 4172 52220 4228
rect 52276 4172 52286 4228
rect 53666 4172 53676 4228
rect 53732 4172 55468 4228
rect 55524 4172 55534 4228
rect 57698 4172 57708 4228
rect 57764 4172 59948 4228
rect 60004 4172 60014 4228
rect 61842 4172 61852 4228
rect 61908 4172 62972 4228
rect 63028 4172 63038 4228
rect 65762 4172 65772 4228
rect 65828 4172 67340 4228
rect 67396 4172 67406 4228
rect 70914 4172 70924 4228
rect 70980 4172 71932 4228
rect 71988 4172 71998 4228
rect 47618 4060 47628 4116
rect 47684 4060 48748 4116
rect 48804 4060 50540 4116
rect 50596 4060 50606 4116
rect 63746 4060 63756 4116
rect 63812 4060 66108 4116
rect 66164 4060 66174 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 50194 3724 50204 3780
rect 50260 3724 52108 3780
rect 52164 3724 52780 3780
rect 52836 3724 52846 3780
rect 59714 3724 59724 3780
rect 59780 3724 61740 3780
rect 61796 3724 61806 3780
rect 69122 3724 69132 3780
rect 69188 3724 70028 3780
rect 70084 3724 70094 3780
rect 74162 3724 74172 3780
rect 74228 3724 75628 3780
rect 75684 3724 76300 3780
rect 76356 3724 76366 3780
rect 7970 3612 7980 3668
rect 8036 3612 8652 3668
rect 8708 3612 9548 3668
rect 9604 3612 9614 3668
rect 37874 3612 37884 3668
rect 37940 3612 38892 3668
rect 38948 3612 40124 3668
rect 40180 3612 40190 3668
rect 43586 3612 43596 3668
rect 43652 3612 45948 3668
rect 46004 3612 46844 3668
rect 46900 3612 46910 3668
rect 47842 3612 47852 3668
rect 47908 3612 48860 3668
rect 48916 3612 48926 3668
rect 50306 3612 50316 3668
rect 50372 3612 53564 3668
rect 53620 3612 53630 3668
rect 54338 3612 54348 3668
rect 54404 3612 57372 3668
rect 57428 3612 57438 3668
rect 60386 3612 60396 3668
rect 60452 3612 63084 3668
rect 63140 3612 63150 3668
rect 67442 3612 67452 3668
rect 67508 3612 68348 3668
rect 68404 3612 68414 3668
rect 69906 3612 69916 3668
rect 69972 3612 71260 3668
rect 71316 3612 71326 3668
rect 73826 3612 73836 3668
rect 73892 3612 76972 3668
rect 77028 3612 77038 3668
rect 21858 3500 21868 3556
rect 21924 3500 22540 3556
rect 22596 3500 23324 3556
rect 23380 3500 23390 3556
rect 35522 3500 35532 3556
rect 35588 3500 36204 3556
rect 36260 3500 36988 3556
rect 37044 3500 37054 3556
rect 42914 3500 42924 3556
rect 42980 3500 44268 3556
rect 44324 3500 44334 3556
rect 51650 3500 51660 3556
rect 51716 3500 54012 3556
rect 54068 3500 54078 3556
rect 55794 3500 55804 3556
rect 55860 3500 58156 3556
rect 58212 3500 58222 3556
rect 58370 3500 58380 3556
rect 58436 3500 61292 3556
rect 61348 3500 61358 3556
rect 62514 3500 62524 3556
rect 62580 3500 65212 3556
rect 65268 3500 65278 3556
rect 3938 3388 3948 3444
rect 4004 3388 5740 3444
rect 5796 3388 5806 3444
rect 7858 3388 7868 3444
rect 7924 3388 9324 3444
rect 9380 3388 9996 3444
rect 10052 3388 10062 3444
rect 10882 3388 10892 3444
rect 10948 3388 11676 3444
rect 11732 3388 11742 3444
rect 13794 3388 13804 3444
rect 13860 3388 14700 3444
rect 14756 3388 14766 3444
rect 15362 3388 15372 3444
rect 15428 3388 17612 3444
rect 17668 3388 18060 3444
rect 18116 3388 18126 3444
rect 23426 3388 23436 3444
rect 23492 3388 25340 3444
rect 25396 3388 25406 3444
rect 27458 3388 27468 3444
rect 27524 3388 29708 3444
rect 29764 3388 29774 3444
rect 31378 3388 31388 3444
rect 31444 3388 33180 3444
rect 33236 3388 33246 3444
rect 34402 3388 34412 3444
rect 34468 3388 35196 3444
rect 35252 3388 36876 3444
rect 36932 3388 36942 3444
rect 38322 3388 38332 3444
rect 38388 3388 39564 3444
rect 39620 3388 39630 3444
rect 41570 3388 41580 3444
rect 41636 3388 42812 3444
rect 42868 3388 43708 3444
rect 43764 3388 43774 3444
rect 45602 3388 45612 3444
rect 45668 3388 48188 3444
rect 48244 3388 49868 3444
rect 49924 3388 49934 3444
rect 52322 3388 52332 3444
rect 52388 3388 55692 3444
rect 55748 3388 55758 3444
rect 56354 3388 56364 3444
rect 56420 3388 59164 3444
rect 59220 3388 59230 3444
rect 64418 3388 64428 3444
rect 64484 3388 66444 3444
rect 66500 3388 66510 3444
rect 71138 3388 71148 3444
rect 71204 3388 72716 3444
rect 72772 3388 73388 3444
rect 73444 3388 73454 3444
rect 74498 3388 74508 3444
rect 74564 3388 75068 3444
rect 75124 3388 76412 3444
rect 76468 3388 76478 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 76076 4768 76892
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 76860 20128 76892
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 76076 35488 76892
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 76860 50848 76892
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 76076 66208 76892
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__I dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 72240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A1
timestamp 1669390400
transform 1 0 21056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A2
timestamp 1669390400
transform 1 0 19936 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A3
timestamp 1669390400
transform 1 0 21504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A4
timestamp 1669390400
transform 1 0 21952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__A1
timestamp 1669390400
transform -1 0 25088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__A2
timestamp 1669390400
transform 1 0 25312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__A1
timestamp 1669390400
transform 1 0 24416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__A2
timestamp 1669390400
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__A1
timestamp 1669390400
transform 1 0 16688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__A2
timestamp 1669390400
transform 1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__A3
timestamp 1669390400
transform 1 0 19040 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__A4
timestamp 1669390400
transform 1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__A1
timestamp 1669390400
transform 1 0 23856 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__A2
timestamp 1669390400
transform 1 0 22288 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__A3
timestamp 1669390400
transform 1 0 24304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__A4
timestamp 1669390400
transform 1 0 24080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__A1
timestamp 1669390400
transform 1 0 54096 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__A2
timestamp 1669390400
transform 1 0 53648 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__A3
timestamp 1669390400
transform 1 0 54544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__A1
timestamp 1669390400
transform 1 0 54096 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__A2
timestamp 1669390400
transform 1 0 54544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__A3
timestamp 1669390400
transform 1 0 53648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__I
timestamp 1669390400
transform -1 0 56784 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__I
timestamp 1669390400
transform 1 0 66976 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__I
timestamp 1669390400
transform 1 0 56672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__A2
timestamp 1669390400
transform 1 0 54544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__A3
timestamp 1669390400
transform 1 0 54992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__I
timestamp 1669390400
transform -1 0 56448 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__I
timestamp 1669390400
transform -1 0 66864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__I
timestamp 1669390400
transform -1 0 74144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__A2
timestamp 1669390400
transform 1 0 73024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__B1
timestamp 1669390400
transform 1 0 72576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I
timestamp 1669390400
transform -1 0 66752 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__A2
timestamp 1669390400
transform -1 0 68992 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__B1
timestamp 1669390400
transform -1 0 70112 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__I
timestamp 1669390400
transform 1 0 48048 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I
timestamp 1669390400
transform 1 0 55664 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__I
timestamp 1669390400
transform -1 0 55664 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__I
timestamp 1669390400
transform 1 0 51296 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1669390400
transform -1 0 50288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__I
timestamp 1669390400
transform 1 0 48720 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__I
timestamp 1669390400
transform -1 0 51296 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I
timestamp 1669390400
transform 1 0 47152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__I
timestamp 1669390400
transform 1 0 51968 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__I
timestamp 1669390400
transform -1 0 49056 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__I
timestamp 1669390400
transform -1 0 52416 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__I
timestamp 1669390400
transform -1 0 49616 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__I
timestamp 1669390400
transform 1 0 52192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__I
timestamp 1669390400
transform -1 0 60032 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__I
timestamp 1669390400
transform 1 0 48832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__I
timestamp 1669390400
transform -1 0 61488 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__146__I
timestamp 1669390400
transform 1 0 47712 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__I
timestamp 1669390400
transform 1 0 58016 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__I
timestamp 1669390400
transform 1 0 50960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__I
timestamp 1669390400
transform -1 0 54208 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__I
timestamp 1669390400
transform 1 0 53312 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I
timestamp 1669390400
transform -1 0 54880 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__155__I
timestamp 1669390400
transform -1 0 53760 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__I
timestamp 1669390400
transform 1 0 51520 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__I
timestamp 1669390400
transform -1 0 56560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__I
timestamp 1669390400
transform 1 0 51184 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__I
timestamp 1669390400
transform 1 0 57344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__I
timestamp 1669390400
transform 1 0 53648 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__I
timestamp 1669390400
transform -1 0 57904 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__I
timestamp 1669390400
transform -1 0 56224 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__I
timestamp 1669390400
transform 1 0 56336 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__I
timestamp 1669390400
transform -1 0 59584 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__I
timestamp 1669390400
transform 1 0 54544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I
timestamp 1669390400
transform 1 0 63280 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__I
timestamp 1669390400
transform 1 0 56560 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I
timestamp 1669390400
transform -1 0 59920 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__I
timestamp 1669390400
transform -1 0 56784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1669390400
transform 1 0 58912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I
timestamp 1669390400
transform 1 0 58464 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1669390400
transform 1 0 61824 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I
timestamp 1669390400
transform 1 0 59024 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I
timestamp 1669390400
transform -1 0 62160 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I
timestamp 1669390400
transform -1 0 57904 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1669390400
transform -1 0 67200 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__I
timestamp 1669390400
transform 1 0 58016 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I
timestamp 1669390400
transform 1 0 65296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__I
timestamp 1669390400
transform -1 0 59920 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__I
timestamp 1669390400
transform -1 0 62272 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__I
timestamp 1669390400
transform 1 0 61936 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__I
timestamp 1669390400
transform 1 0 62720 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__I
timestamp 1669390400
transform 1 0 62272 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I
timestamp 1669390400
transform -1 0 61264 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__I
timestamp 1669390400
transform 1 0 60144 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__I
timestamp 1669390400
transform 1 0 68656 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__I
timestamp 1669390400
transform 1 0 59808 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I
timestamp 1669390400
transform -1 0 63840 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__I
timestamp 1669390400
transform 1 0 61600 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I
timestamp 1669390400
transform -1 0 65072 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__I
timestamp 1669390400
transform -1 0 60816 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I
timestamp 1669390400
transform 1 0 65968 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__I
timestamp 1669390400
transform 1 0 65296 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__I
timestamp 1669390400
transform 1 0 67088 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__I
timestamp 1669390400
transform 1 0 62496 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__I
timestamp 1669390400
transform 1 0 64848 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__I
timestamp 1669390400
transform 1 0 63840 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__I
timestamp 1669390400
transform 1 0 67424 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__I
timestamp 1669390400
transform 1 0 63952 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__I
timestamp 1669390400
transform -1 0 66864 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__I
timestamp 1669390400
transform -1 0 66416 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__I
timestamp 1669390400
transform 1 0 68432 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__I
timestamp 1669390400
transform 1 0 67088 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__I
timestamp 1669390400
transform 1 0 73696 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__A2
timestamp 1669390400
transform 1 0 74368 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__I
timestamp 1669390400
transform 1 0 74368 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__A2
timestamp 1669390400
transform -1 0 74144 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__A2
timestamp 1669390400
transform 1 0 70112 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__A2
timestamp 1669390400
transform -1 0 69776 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__I
timestamp 1669390400
transform 1 0 13552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__I
timestamp 1669390400
transform 1 0 13888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__I
timestamp 1669390400
transform 1 0 56672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__I
timestamp 1669390400
transform 1 0 54992 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__I
timestamp 1669390400
transform 1 0 56784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__I
timestamp 1669390400
transform 1 0 55440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__I
timestamp 1669390400
transform 1 0 20160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__I
timestamp 1669390400
transform 1 0 20384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__I
timestamp 1669390400
transform 1 0 17584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__I
timestamp 1669390400
transform -1 0 17248 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__I
timestamp 1669390400
transform 1 0 19712 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__I
timestamp 1669390400
transform 1 0 21504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__I
timestamp 1669390400
transform 1 0 22400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__I
timestamp 1669390400
transform 1 0 21616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__I
timestamp 1669390400
transform -1 0 22848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__I
timestamp 1669390400
transform 1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__I
timestamp 1669390400
transform -1 0 24416 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__I
timestamp 1669390400
transform 1 0 23744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__I
timestamp 1669390400
transform -1 0 24976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__I
timestamp 1669390400
transform 1 0 23072 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__I
timestamp 1669390400
transform 1 0 26096 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__I
timestamp 1669390400
transform 1 0 26544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__I
timestamp 1669390400
transform -1 0 12096 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__280__I
timestamp 1669390400
transform -1 0 12992 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__I
timestamp 1669390400
transform -1 0 12096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__I
timestamp 1669390400
transform 1 0 14112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__283__I
timestamp 1669390400
transform 1 0 14784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__I
timestamp 1669390400
transform 1 0 15456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__I
timestamp 1669390400
transform 1 0 16352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__I
timestamp 1669390400
transform -1 0 16464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__I
timestamp 1669390400
transform 1 0 17136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__288__I
timestamp 1669390400
transform -1 0 18256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__I
timestamp 1669390400
transform 1 0 19264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__I
timestamp 1669390400
transform -1 0 18368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__291__I
timestamp 1669390400
transform 1 0 20160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__I
timestamp 1669390400
transform -1 0 19600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__I
timestamp 1669390400
transform -1 0 21056 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__I
timestamp 1669390400
transform 1 0 23072 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__I
timestamp 1669390400
transform 1 0 22624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__I
timestamp 1669390400
transform -1 0 23184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__I
timestamp 1669390400
transform 1 0 24304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__I
timestamp 1669390400
transform -1 0 22848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__I
timestamp 1669390400
transform -1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__I
timestamp 1669390400
transform 1 0 27552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__I
timestamp 1669390400
transform 1 0 27104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__I
timestamp 1669390400
transform -1 0 28896 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__I
timestamp 1669390400
transform 1 0 29792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__I
timestamp 1669390400
transform 1 0 29344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__I
timestamp 1669390400
transform 1 0 31472 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__I
timestamp 1669390400
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__I
timestamp 1669390400
transform 1 0 31024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__I
timestamp 1669390400
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__I
timestamp 1669390400
transform 1 0 33936 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__I
timestamp 1669390400
transform 1 0 33488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__I
timestamp 1669390400
transform 1 0 34384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__I
timestamp 1669390400
transform 1 0 36176 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__I
timestamp 1669390400
transform 1 0 35728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__314__I
timestamp 1669390400
transform 1 0 37408 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__I
timestamp 1669390400
transform 1 0 37856 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__I
timestamp 1669390400
transform 1 0 37408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__I
timestamp 1669390400
transform 1 0 39312 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__318__I
timestamp 1669390400
transform 1 0 38864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__I
timestamp 1669390400
transform 1 0 39536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__I
timestamp 1669390400
transform -1 0 38528 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__321__I
timestamp 1669390400
transform 1 0 40320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__I
timestamp 1669390400
transform 1 0 42784 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__323__I
timestamp 1669390400
transform 1 0 42336 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__I
timestamp 1669390400
transform 1 0 42896 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__I
timestamp 1669390400
transform -1 0 44352 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__I
timestamp 1669390400
transform 1 0 44912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__I
timestamp 1669390400
transform -1 0 46480 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__I
timestamp 1669390400
transform 1 0 46704 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__I
timestamp 1669390400
transform 1 0 48272 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__I
timestamp 1669390400
transform -1 0 48272 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__I
timestamp 1669390400
transform 1 0 48160 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__332__I
timestamp 1669390400
transform 1 0 48832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__I
timestamp 1669390400
transform -1 0 25872 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__I
timestamp 1669390400
transform -1 0 26544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__I
timestamp 1669390400
transform -1 0 27216 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__I
timestamp 1669390400
transform -1 0 27888 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__I
timestamp 1669390400
transform -1 0 28560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__I
timestamp 1669390400
transform -1 0 29456 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__I
timestamp 1669390400
transform -1 0 30800 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__I
timestamp 1669390400
transform 1 0 32144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__I
timestamp 1669390400
transform -1 0 31248 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__I
timestamp 1669390400
transform -1 0 31920 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__I
timestamp 1669390400
transform -1 0 32592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__I
timestamp 1669390400
transform 1 0 34832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__I
timestamp 1669390400
transform -1 0 33936 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__I
timestamp 1669390400
transform -1 0 35504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__I
timestamp 1669390400
transform 1 0 38304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__I
timestamp 1669390400
transform -1 0 35952 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__I
timestamp 1669390400
transform -1 0 36624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__I
timestamp 1669390400
transform 1 0 39984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__I
timestamp 1669390400
transform -1 0 37968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__I
timestamp 1669390400
transform -1 0 39088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__I
timestamp 1669390400
transform -1 0 40208 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__I
timestamp 1669390400
transform 1 0 41440 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__I
timestamp 1669390400
transform -1 0 40656 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__I
timestamp 1669390400
transform 1 0 43568 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__I
timestamp 1669390400
transform -1 0 42000 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__I
timestamp 1669390400
transform -1 0 42672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__I
timestamp 1669390400
transform -1 0 44688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__I
timestamp 1669390400
transform -1 0 44016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__I
timestamp 1669390400
transform 1 0 47824 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__I
timestamp 1669390400
transform -1 0 47824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__I
timestamp 1669390400
transform -1 0 46032 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__I
timestamp 1669390400
transform -1 0 47824 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__I
timestamp 1669390400
transform 1 0 71680 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__I
timestamp 1669390400
transform -1 0 72576 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__I
timestamp 1669390400
transform 1 0 72800 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__I
timestamp 1669390400
transform -1 0 73696 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__I
timestamp 1669390400
transform -1 0 69552 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__I
timestamp 1669390400
transform -1 0 70224 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__I
timestamp 1669390400
transform -1 0 70896 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__372__I
timestamp 1669390400
transform 1 0 72352 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__I
timestamp 1669390400
transform 1 0 69888 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__374__I
timestamp 1669390400
transform -1 0 71232 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 77392 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform 1 0 4144 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 4256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform -1 0 10976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform 1 0 13888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform -1 0 13552 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform -1 0 14560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform -1 0 13888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform 1 0 18032 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform 1 0 18368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform 1 0 17920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1669390400
transform 1 0 17584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1669390400
transform -1 0 18144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1669390400
transform -1 0 5824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1669390400
transform 1 0 18816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1669390400
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1669390400
transform 1 0 21952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1669390400
transform -1 0 21728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1669390400
transform 1 0 21280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1669390400
transform -1 0 21952 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1669390400
transform -1 0 22848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1669390400
transform 1 0 22512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1669390400
transform 1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1669390400
transform 1 0 25984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1669390400
transform 1 0 6832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1669390400
transform -1 0 25424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1669390400
transform 1 0 26768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1669390400
transform 1 0 8624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1669390400
transform 1 0 9632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1669390400
transform 1 0 9520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1669390400
transform 1 0 9968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1669390400
transform 1 0 11088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1669390400
transform 1 0 11872 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1669390400
transform 1 0 14448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1669390400
transform 1 0 75040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1669390400
transform -1 0 77392 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1669390400
transform -1 0 77392 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1669390400
transform 1 0 76832 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1669390400
transform -1 0 77392 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1669390400
transform 1 0 76832 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1669390400
transform -1 0 77392 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1669390400
transform 1 0 76832 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1669390400
transform -1 0 77392 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1669390400
transform -1 0 74592 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1669390400
transform 1 0 76832 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1669390400
transform -1 0 77392 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1669390400
transform 1 0 76832 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1669390400
transform 1 0 76832 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1669390400
transform -1 0 77392 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1669390400
transform 1 0 76832 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1669390400
transform -1 0 77392 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1669390400
transform -1 0 74592 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1669390400
transform 1 0 76832 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1669390400
transform -1 0 77392 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1669390400
transform 1 0 76832 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1669390400
transform -1 0 77392 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1669390400
transform 1 0 76832 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1669390400
transform -1 0 77392 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1669390400
transform -1 0 77392 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1669390400
transform -1 0 74592 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1669390400
transform 1 0 76832 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1669390400
transform -1 0 77392 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1669390400
transform 1 0 76832 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1669390400
transform -1 0 77392 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1669390400
transform 1 0 76832 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1669390400
transform -1 0 77392 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1669390400
transform 1 0 76832 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1669390400
transform 1 0 4144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1669390400
transform 1 0 3696 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1669390400
transform 1 0 3696 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1669390400
transform 1 0 4144 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1669390400
transform 1 0 3696 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1669390400
transform 1 0 4144 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1669390400
transform 1 0 3696 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1669390400
transform -1 0 3920 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1669390400
transform 1 0 3696 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1669390400
transform 1 0 3696 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1669390400
transform 1 0 4144 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1669390400
transform 1 0 3696 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1669390400
transform 1 0 3696 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1669390400
transform 1 0 4144 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1669390400
transform 1 0 3696 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1669390400
transform -1 0 3920 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input84_I
timestamp 1669390400
transform 1 0 3696 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input85_I
timestamp 1669390400
transform 1 0 3696 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input86_I
timestamp 1669390400
transform 1 0 4144 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input87_I
timestamp 1669390400
transform 1 0 3696 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input88_I
timestamp 1669390400
transform 1 0 4144 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input89_I
timestamp 1669390400
transform 1 0 3696 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input90_I
timestamp 1669390400
transform 1 0 3696 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input91_I
timestamp 1669390400
transform -1 0 3920 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input92_I
timestamp 1669390400
transform 1 0 3696 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input93_I
timestamp 1669390400
transform 1 0 3696 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input94_I
timestamp 1669390400
transform 1 0 3696 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input95_I
timestamp 1669390400
transform 1 0 3696 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input96_I
timestamp 1669390400
transform 1 0 3696 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input97_I
timestamp 1669390400
transform 1 0 3696 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input98_I
timestamp 1669390400
transform 1 0 3696 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input99_I
timestamp 1669390400
transform 1 0 3696 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input100_I
timestamp 1669390400
transform -1 0 26656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input101_I
timestamp 1669390400
transform -1 0 33264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input102_I
timestamp 1669390400
transform 1 0 34496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input103_I
timestamp 1669390400
transform -1 0 34720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input104_I
timestamp 1669390400
transform 1 0 37408 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input105_I
timestamp 1669390400
transform 1 0 36960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input106_I
timestamp 1669390400
transform -1 0 34496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input107_I
timestamp 1669390400
transform 1 0 38752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input108_I
timestamp 1669390400
transform -1 0 38080 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input109_I
timestamp 1669390400
transform -1 0 37968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input110_I
timestamp 1669390400
transform -1 0 38416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input111_I
timestamp 1669390400
transform 1 0 29456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input112_I
timestamp 1669390400
transform -1 0 40320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input113_I
timestamp 1669390400
transform 1 0 41216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input114_I
timestamp 1669390400
transform 1 0 43680 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input115_I
timestamp 1669390400
transform -1 0 42336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input116_I
timestamp 1669390400
transform -1 0 44352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input117_I
timestamp 1669390400
transform 1 0 46816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input118_I
timestamp 1669390400
transform -1 0 45472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input119_I
timestamp 1669390400
transform -1 0 44912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input120_I
timestamp 1669390400
transform -1 0 48272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input121_I
timestamp 1669390400
transform 1 0 47488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input122_I
timestamp 1669390400
transform 1 0 29904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input123_I
timestamp 1669390400
transform -1 0 46816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input124_I
timestamp 1669390400
transform 1 0 48720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input125_I
timestamp 1669390400
transform 1 0 29120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input126_I
timestamp 1669390400
transform 1 0 31024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input127_I
timestamp 1669390400
transform -1 0 29792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input128_I
timestamp 1669390400
transform -1 0 30912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input129_I
timestamp 1669390400
transform 1 0 33488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input130_I
timestamp 1669390400
transform 1 0 33488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input131_I
timestamp 1669390400
transform 1 0 33936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input132_I
timestamp 1669390400
transform -1 0 70336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input133_I
timestamp 1669390400
transform -1 0 72800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input134_I
timestamp 1669390400
transform -1 0 71680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input135_I
timestamp 1669390400
transform -1 0 73472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input136_I
timestamp 1669390400
transform -1 0 73920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input137_I
timestamp 1669390400
transform -1 0 69664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output138_I
timestamp 1669390400
transform -1 0 75712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output139_I
timestamp 1669390400
transform -1 0 76608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output140_I
timestamp 1669390400
transform -1 0 74592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output141_I
timestamp 1669390400
transform -1 0 74592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output142_I
timestamp 1669390400
transform -1 0 74592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output143_I
timestamp 1669390400
transform -1 0 74592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output144_I
timestamp 1669390400
transform -1 0 74592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output145_I
timestamp 1669390400
transform -1 0 74592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output146_I
timestamp 1669390400
transform 1 0 77168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output147_I
timestamp 1669390400
transform -1 0 74592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output148_I
timestamp 1669390400
transform -1 0 74592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output149_I
timestamp 1669390400
transform -1 0 74592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output150_I
timestamp 1669390400
transform -1 0 74592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output151_I
timestamp 1669390400
transform -1 0 74592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output152_I
timestamp 1669390400
transform -1 0 74592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output153_I
timestamp 1669390400
transform -1 0 74592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output154_I
timestamp 1669390400
transform 1 0 77168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output155_I
timestamp 1669390400
transform -1 0 74592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output156_I
timestamp 1669390400
transform -1 0 74592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output157_I
timestamp 1669390400
transform -1 0 74592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output158_I
timestamp 1669390400
transform -1 0 74592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output159_I
timestamp 1669390400
transform -1 0 74592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output160_I
timestamp 1669390400
transform -1 0 74592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output161_I
timestamp 1669390400
transform 1 0 77168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output162_I
timestamp 1669390400
transform 1 0 77168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output163_I
timestamp 1669390400
transform -1 0 74592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output164_I
timestamp 1669390400
transform -1 0 74592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output165_I
timestamp 1669390400
transform -1 0 74592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output166_I
timestamp 1669390400
transform -1 0 74592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output167_I
timestamp 1669390400
transform -1 0 74592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output168_I
timestamp 1669390400
transform -1 0 74592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output169_I
timestamp 1669390400
transform -1 0 74592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output170_I
timestamp 1669390400
transform 1 0 77168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output172_I
timestamp 1669390400
transform -1 0 4144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output173_I
timestamp 1669390400
transform -1 0 3696 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output174_I
timestamp 1669390400
transform -1 0 3696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output175_I
timestamp 1669390400
transform -1 0 3696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output176_I
timestamp 1669390400
transform -1 0 3696 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output177_I
timestamp 1669390400
transform -1 0 3696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output178_I
timestamp 1669390400
transform -1 0 5488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output179_I
timestamp 1669390400
transform -1 0 4144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output180_I
timestamp 1669390400
transform -1 0 3696 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output181_I
timestamp 1669390400
transform -1 0 3696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output183_I
timestamp 1669390400
transform -1 0 3696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output184_I
timestamp 1669390400
transform -1 0 3696 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output185_I
timestamp 1669390400
transform -1 0 3696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output186_I
timestamp 1669390400
transform -1 0 5488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output187_I
timestamp 1669390400
transform -1 0 4144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output188_I
timestamp 1669390400
transform -1 0 3696 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output189_I
timestamp 1669390400
transform -1 0 3696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output190_I
timestamp 1669390400
transform -1 0 3696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output191_I
timestamp 1669390400
transform -1 0 3696 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output192_I
timestamp 1669390400
transform -1 0 3696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output194_I
timestamp 1669390400
transform -1 0 5488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output195_I
timestamp 1669390400
transform -1 0 4144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output204_I
timestamp 1669390400
transform 1 0 3472 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output205_I
timestamp 1669390400
transform 1 0 51632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output206_I
timestamp 1669390400
transform -1 0 55104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output207_I
timestamp 1669390400
transform 1 0 57344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output208_I
timestamp 1669390400
transform 1 0 58128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output209_I
timestamp 1669390400
transform 1 0 58688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output210_I
timestamp 1669390400
transform 1 0 59584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output211_I
timestamp 1669390400
transform 1 0 60256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output212_I
timestamp 1669390400
transform 1 0 59136 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output213_I
timestamp 1669390400
transform 1 0 61488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output214_I
timestamp 1669390400
transform 1 0 62048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output215_I
timestamp 1669390400
transform -1 0 61264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output216_I
timestamp 1669390400
transform 1 0 51184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output217_I
timestamp 1669390400
transform 1 0 64512 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output218_I
timestamp 1669390400
transform 1 0 64176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output219_I
timestamp 1669390400
transform 1 0 65296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output220_I
timestamp 1669390400
transform 1 0 65744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output221_I
timestamp 1669390400
transform 1 0 68320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output222_I
timestamp 1669390400
transform 1 0 66304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output223_I
timestamp 1669390400
transform 1 0 68880 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output224_I
timestamp 1669390400
transform 1 0 66752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output225_I
timestamp 1669390400
transform 1 0 66752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output226_I
timestamp 1669390400
transform -1 0 69552 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output227_I
timestamp 1669390400
transform -1 0 51632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output228_I
timestamp 1669390400
transform 1 0 70784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output229_I
timestamp 1669390400
transform -1 0 68768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output230_I
timestamp 1669390400
transform -1 0 52192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output231_I
timestamp 1669390400
transform -1 0 51184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output232_I
timestamp 1669390400
transform 1 0 52976 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output233_I
timestamp 1669390400
transform 1 0 54208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output234_I
timestamp 1669390400
transform 1 0 55328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output235_I
timestamp 1669390400
transform 1 0 55776 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output236_I
timestamp 1669390400
transform 1 0 56336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output237_I
timestamp 1669390400
transform -1 0 74592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output238_I
timestamp 1669390400
transform -1 0 74592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output239_I
timestamp 1669390400
transform -1 0 74592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output240_I
timestamp 1669390400
transform 1 0 77168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output241_I
timestamp 1669390400
transform -1 0 74592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output242_I
timestamp 1669390400
transform -1 0 74592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output243_I
timestamp 1669390400
transform -1 0 74592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output244_I
timestamp 1669390400
transform -1 0 74592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output245_I
timestamp 1669390400
transform -1 0 74592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output246_I
timestamp 1669390400
transform -1 0 74592 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output247_I
timestamp 1669390400
transform -1 0 74592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output248_I
timestamp 1669390400
transform -1 0 74592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output249_I
timestamp 1669390400
transform -1 0 74592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output250_I
timestamp 1669390400
transform 1 0 74368 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output251_I
timestamp 1669390400
transform -1 0 74592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output252_I
timestamp 1669390400
transform 1 0 74368 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output253_I
timestamp 1669390400
transform -1 0 74592 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output254_I
timestamp 1669390400
transform 1 0 74368 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output255_I
timestamp 1669390400
transform -1 0 74592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output256_I
timestamp 1669390400
transform 1 0 74368 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output257_I
timestamp 1669390400
transform -1 0 74592 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output258_I
timestamp 1669390400
transform 1 0 74368 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output259_I
timestamp 1669390400
transform -1 0 74592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output260_I
timestamp 1669390400
transform -1 0 74592 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output261_I
timestamp 1669390400
transform 1 0 77168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output262_I
timestamp 1669390400
transform -1 0 74592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output263_I
timestamp 1669390400
transform -1 0 74592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output264_I
timestamp 1669390400
transform 1 0 77168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output265_I
timestamp 1669390400
transform -1 0 74592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output266_I
timestamp 1669390400
transform -1 0 74592 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output267_I
timestamp 1669390400
transform -1 0 74592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output268_I
timestamp 1669390400
transform -1 0 74592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output269_I
timestamp 1669390400
transform -1 0 3696 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output270_I
timestamp 1669390400
transform -1 0 3696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output271_I
timestamp 1669390400
transform -1 0 3696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output272_I
timestamp 1669390400
transform -1 0 5488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output273_I
timestamp 1669390400
transform -1 0 4144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output274_I
timestamp 1669390400
transform -1 0 3696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output275_I
timestamp 1669390400
transform -1 0 3696 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output276_I
timestamp 1669390400
transform -1 0 3696 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output277_I
timestamp 1669390400
transform -1 0 3696 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output278_I
timestamp 1669390400
transform -1 0 3696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output279_I
timestamp 1669390400
transform -1 0 3696 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output280_I
timestamp 1669390400
transform -1 0 3696 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output281_I
timestamp 1669390400
transform -1 0 3696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output282_I
timestamp 1669390400
transform 1 0 3472 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output283_I
timestamp 1669390400
transform -1 0 3696 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output284_I
timestamp 1669390400
transform 1 0 3472 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output285_I
timestamp 1669390400
transform -1 0 3696 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output286_I
timestamp 1669390400
transform 1 0 3472 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output287_I
timestamp 1669390400
transform -1 0 3696 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output288_I
timestamp 1669390400
transform 1 0 3472 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output289_I
timestamp 1669390400
transform -1 0 3696 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output290_I
timestamp 1669390400
transform 1 0 3472 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output291_I
timestamp 1669390400
transform -1 0 3696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output292_I
timestamp 1669390400
transform -1 0 3920 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output293_I
timestamp 1669390400
transform -1 0 5488 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output294_I
timestamp 1669390400
transform -1 0 3696 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output295_I
timestamp 1669390400
transform -1 0 3696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output296_I
timestamp 1669390400
transform -1 0 5488 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output297_I
timestamp 1669390400
transform -1 0 4144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output298_I
timestamp 1669390400
transform -1 0 3696 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output299_I
timestamp 1669390400
transform -1 0 3696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output300_I
timestamp 1669390400
transform -1 0 3696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output305_I
timestamp 1669390400
transform 1 0 3920 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output306_I
timestamp 1669390400
transform -1 0 5488 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output307_I
timestamp 1669390400
transform -1 0 3920 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output308_I
timestamp 1669390400
transform -1 0 5488 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output310_I
timestamp 1669390400
transform -1 0 3696 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output312_I
timestamp 1669390400
transform -1 0 3696 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48
timestamp 1669390400
transform 1 0 6720 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75
timestamp 1669390400
transform 1 0 9744 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10192 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83
timestamp 1669390400
transform 1 0 10640 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86
timestamp 1669390400
transform 1 0 10976 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109
timestamp 1669390400
transform 1 0 13552 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112
timestamp 1669390400
transform 1 0 13888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_168
timestamp 1669390400
transform 1 0 20160 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_172
timestamp 1669390400
transform 1 0 20608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1669390400
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_180
timestamp 1669390400
transform 1 0 21504 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_188
timestamp 1669390400
transform 1 0 22400 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_191
timestamp 1669390400
transform 1 0 22736 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_215
timestamp 1669390400
transform 1 0 25424 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_223
timestamp 1669390400
transform 1 0 26320 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_227
timestamp 1669390400
transform 1 0 26768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_250
timestamp 1669390400
transform 1 0 29344 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_254
timestamp 1669390400
transform 1 0 29792 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_262
timestamp 1669390400
transform 1 0 30688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1669390400
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_285
timestamp 1669390400
transform 1 0 33264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_293
timestamp 1669390400
transform 1 0 34160 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_296
timestamp 1669390400
transform 1 0 34496 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1669390400
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_320
timestamp 1669390400
transform 1 0 37184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_324
timestamp 1669390400
transform 1 0 37632 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_327
timestamp 1669390400
transform 1 0 37968 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_331
timestamp 1669390400
transform 1 0 38416 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_358
timestamp 1669390400
transform 1 0 41440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_376
timestamp 1669390400
transform 1 0 43456 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_380
timestamp 1669390400
transform 1 0 43904 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1669390400
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_404
timestamp 1669390400
transform 1 0 46592 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_408
timestamp 1669390400
transform 1 0 47040 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_416
timestamp 1669390400
transform 1 0 47936 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1669390400
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_439
timestamp 1669390400
transform 1 0 50512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_445
timestamp 1669390400
transform 1 0 51184 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_449
timestamp 1669390400
transform 1 0 51632 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_451
timestamp 1669390400
transform 1 0 51856 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1669390400
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_472
timestamp 1669390400
transform 1 0 54208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_488
timestamp 1669390400
transform 1 0 56000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_507
timestamp 1669390400
transform 1 0 58128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_523
timestamp 1669390400
transform 1 0 59920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_527
timestamp 1669390400
transform 1 0 60368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_542
timestamp 1669390400
transform 1 0 62048 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_558
timestamp 1669390400
transform 1 0 63840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_562
timestamp 1669390400
transform 1 0 64288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_577
timestamp 1669390400
transform 1 0 65968 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_593
timestamp 1669390400
transform 1 0 67760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1669390400
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_600
timestamp 1669390400
transform 1 0 68544 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_610
timestamp 1669390400
transform 1 0 69664 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_628
timestamp 1669390400
transform 1 0 71680 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_632
timestamp 1669390400
transform 1 0 72128 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_649
timestamp 1669390400
transform 1 0 74032 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_657
timestamp 1669390400
transform 1 0 74928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_660
timestamp 1669390400
transform 1 0 75264 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1669390400
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1669390400
transform 1 0 76048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_682
timestamp 1669390400
transform 1 0 77728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_686
timestamp 1669390400
transform 1 0 78176 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_18
timestamp 1669390400
transform 1 0 3360 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_26
timestamp 1669390400
transform 1 0 4256 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_34
timestamp 1669390400
transform 1 0 5152 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_52
timestamp 1669390400
transform 1 0 7168 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_76
timestamp 1669390400
transform 1 0 9856 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_94
timestamp 1669390400
transform 1 0 11872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_112
timestamp 1669390400
transform 1 0 13888 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_139
timestamp 1669390400
transform 1 0 16912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_147
timestamp 1669390400
transform 1 0 17808 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_151
timestamp 1669390400
transform 1 0 18256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_155
timestamp 1669390400
transform 1 0 18704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_158
timestamp 1669390400
transform 1 0 19040 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_176
timestamp 1669390400
transform 1 0 21056 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_194
timestamp 1669390400
transform 1 0 23072 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_218
timestamp 1669390400
transform 1 0 25760 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_222
timestamp 1669390400
transform 1 0 26208 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_226
timestamp 1669390400
transform 1 0 26656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_229
timestamp 1669390400
transform 1 0 26992 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_247
timestamp 1669390400
transform 1 0 29008 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_265
timestamp 1669390400
transform 1 0 31024 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_289
timestamp 1669390400
transform 1 0 33712 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_293
timestamp 1669390400
transform 1 0 34160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_295
timestamp 1669390400
transform 1 0 34384 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_298
timestamp 1669390400
transform 1 0 34720 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_316
timestamp 1669390400
transform 1 0 36736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_334
timestamp 1669390400
transform 1 0 38752 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_352
timestamp 1669390400
transform 1 0 40768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_374
timestamp 1669390400
transform 1 0 43232 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_392
timestamp 1669390400
transform 1 0 45248 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_410
timestamp 1669390400
transform 1 0 47264 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_414
timestamp 1669390400
transform 1 0 47712 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_422
timestamp 1669390400
transform 1 0 48608 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_445
timestamp 1669390400
transform 1 0 51184 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_461
timestamp 1669390400
transform 1 0 52976 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_477
timestamp 1669390400
transform 1 0 54768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_493
timestamp 1669390400
transform 1 0 56560 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_514
timestamp 1669390400
transform 1 0 58912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_530
timestamp 1669390400
transform 1 0 60704 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_546
timestamp 1669390400
transform 1 0 62496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_562
timestamp 1669390400
transform 1 0 64288 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_566
timestamp 1669390400
transform 1 0 64736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1669390400
transform 1 0 65184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_585
timestamp 1669390400
transform 1 0 66864 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_601
timestamp 1669390400
transform 1 0 68656 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_605
timestamp 1669390400
transform 1 0 69104 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_609
timestamp 1669390400
transform 1 0 69552 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_613
timestamp 1669390400
transform 1 0 70000 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_616
timestamp 1669390400
transform 1 0 70336 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_634
timestamp 1669390400
transform 1 0 72352 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_638
timestamp 1669390400
transform 1 0 72800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1669390400
transform 1 0 73136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_658
timestamp 1669390400
transform 1 0 75040 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_676
timestamp 1669390400
transform 1 0 77056 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_684
timestamp 1669390400
transform 1 0 77952 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_17
timestamp 1669390400
transform 1 0 3248 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_25
timestamp 1669390400
transform 1 0 4144 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_27
timestamp 1669390400
transform 1 0 4368 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_41
timestamp 1669390400
transform 1 0 5936 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_43
timestamp 1669390400
transform 1 0 6160 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_50
timestamp 1669390400
transform 1 0 6944 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_52
timestamp 1669390400
transform 1 0 7168 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_69
timestamp 1669390400
transform 1 0 9072 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_87
timestamp 1669390400
transform 1 0 11088 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_115
timestamp 1669390400
transform 1 0 14224 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_119
timestamp 1669390400
transform 1 0 14672 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_123
timestamp 1669390400
transform 1 0 15120 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_140
timestamp 1669390400
transform 1 0 17024 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_158
timestamp 1669390400
transform 1 0 19040 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_182
timestamp 1669390400
transform 1 0 21728 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_186
timestamp 1669390400
transform 1 0 22176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_192
timestamp 1669390400
transform 1 0 22848 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_194
timestamp 1669390400
transform 1 0 23072 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_211
timestamp 1669390400
transform 1 0 24976 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_229
timestamp 1669390400
transform 1 0 26992 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_253
timestamp 1669390400
transform 1 0 29680 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_257
timestamp 1669390400
transform 1 0 30128 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_261
timestamp 1669390400
transform 1 0 30576 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_264
timestamp 1669390400
transform 1 0 30912 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_282
timestamp 1669390400
transform 1 0 32928 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_300
timestamp 1669390400
transform 1 0 34944 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_324
timestamp 1669390400
transform 1 0 37632 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_328
timestamp 1669390400
transform 1 0 38080 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_346
timestamp 1669390400
transform 1 0 40096 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_364
timestamp 1669390400
transform 1 0 42112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_382
timestamp 1669390400
transform 1 0 44128 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_386
timestamp 1669390400
transform 1 0 44576 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_409
timestamp 1669390400
transform 1 0 47152 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_427
timestamp 1669390400
transform 1 0 49168 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_443
timestamp 1669390400
transform 1 0 50960 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_459
timestamp 1669390400
transform 1 0 52752 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_478
timestamp 1669390400
transform 1 0 54880 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_494
timestamp 1669390400
transform 1 0 56672 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_512
timestamp 1669390400
transform 1 0 58688 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_530
timestamp 1669390400
transform 1 0 60704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_534
timestamp 1669390400
transform 1 0 61152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_549
timestamp 1669390400
transform 1 0 62832 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_551
timestamp 1669390400
transform 1 0 63056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_566
timestamp 1669390400
transform 1 0 64736 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_584
timestamp 1669390400
transform 1 0 66752 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_600
timestamp 1669390400
transform 1 0 68544 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_602
timestamp 1669390400
transform 1 0 68768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1669390400
transform 1 0 69104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_620
timestamp 1669390400
transform 1 0 70784 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_624
timestamp 1669390400
transform 1 0 71232 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_628
timestamp 1669390400
transform 1 0 71680 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_646
timestamp 1669390400
transform 1 0 73696 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_664
timestamp 1669390400
transform 1 0 75712 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_668
timestamp 1669390400
transform 1 0 76160 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_672
timestamp 1669390400
transform 1 0 76608 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_676
timestamp 1669390400
transform 1 0 77056 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_684
timestamp 1669390400
transform 1 0 77952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_17
timestamp 1669390400
transform 1 0 3248 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_21
timestamp 1669390400
transform 1 0 3696 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_23
timestamp 1669390400
transform 1 0 3920 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_26
timestamp 1669390400
transform 1 0 4256 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_34
timestamp 1669390400
transform 1 0 5152 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_52
timestamp 1669390400
transform 1 0 7168 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_81
timestamp 1669390400
transform 1 0 10416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_85
timestamp 1669390400
transform 1 0 10864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_89
timestamp 1669390400
transform 1 0 11312 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_93
timestamp 1669390400
transform 1 0 11760 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_96
timestamp 1669390400
transform 1 0 12096 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_104
timestamp 1669390400
transform 1 0 12992 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_106
timestamp 1669390400
transform 1 0 13216 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_109
timestamp 1669390400
transform 1 0 13552 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_111
timestamp 1669390400
transform 1 0 13776 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_114
timestamp 1669390400
transform 1 0 14112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_118
timestamp 1669390400
transform 1 0 14560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_122
timestamp 1669390400
transform 1 0 15008 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_124
timestamp 1669390400
transform 1 0 15232 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_150
timestamp 1669390400
transform 1 0 18144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_154
timestamp 1669390400
transform 1 0 18592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_172
timestamp 1669390400
transform 1 0 20608 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_190
timestamp 1669390400
transform 1 0 22624 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1669390400
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_247
timestamp 1669390400
transform 1 0 29008 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_265
timestamp 1669390400
transform 1 0 31024 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_289
timestamp 1669390400
transform 1 0 33712 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_293
timestamp 1669390400
transform 1 0 34160 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_295
timestamp 1669390400
transform 1 0 34384 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_298
timestamp 1669390400
transform 1 0 34720 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_316
timestamp 1669390400
transform 1 0 36736 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_332
timestamp 1669390400
transform 1 0 38528 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_336
timestamp 1669390400
transform 1 0 38976 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_344
timestamp 1669390400
transform 1 0 39872 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_348
timestamp 1669390400
transform 1 0 40320 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_352
timestamp 1669390400
transform 1 0 40768 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_361
timestamp 1669390400
transform 1 0 41776 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_363
timestamp 1669390400
transform 1 0 42000 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_366
timestamp 1669390400
transform 1 0 42336 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_382
timestamp 1669390400
transform 1 0 44128 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_390
timestamp 1669390400
transform 1 0 45024 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_394
timestamp 1669390400
transform 1 0 45472 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_402
timestamp 1669390400
transform 1 0 46368 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_406
timestamp 1669390400
transform 1 0 46816 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_424
timestamp 1669390400
transform 1 0 48832 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_443
timestamp 1669390400
transform 1 0 50960 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_447
timestamp 1669390400
transform 1 0 51408 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_451
timestamp 1669390400
transform 1 0 51856 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_459
timestamp 1669390400
transform 1 0 52752 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_463
timestamp 1669390400
transform 1 0 53200 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_471
timestamp 1669390400
transform 1 0 54096 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_474
timestamp 1669390400
transform 1 0 54432 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_480
timestamp 1669390400
transform 1 0 55104 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_484
timestamp 1669390400
transform 1 0 55552 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_488
timestamp 1669390400
transform 1 0 56000 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_490
timestamp 1669390400
transform 1 0 56224 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_493
timestamp 1669390400
transform 1 0 56560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_502
timestamp 1669390400
transform 1 0 57568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_506
timestamp 1669390400
transform 1 0 58016 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_509
timestamp 1669390400
transform 1 0 58352 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_511
timestamp 1669390400
transform 1 0 58576 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_514
timestamp 1669390400
transform 1 0 58912 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_518
timestamp 1669390400
transform 1 0 59360 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_522
timestamp 1669390400
transform 1 0 59808 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_528
timestamp 1669390400
transform 1 0 60480 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_532
timestamp 1669390400
transform 1 0 60928 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_535
timestamp 1669390400
transform 1 0 61264 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_539
timestamp 1669390400
transform 1 0 61712 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_541
timestamp 1669390400
transform 1 0 61936 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_544
timestamp 1669390400
transform 1 0 62272 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_560
timestamp 1669390400
transform 1 0 64064 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_563
timestamp 1669390400
transform 1 0 64400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1669390400
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_570
timestamp 1669390400
transform 1 0 65184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_573
timestamp 1669390400
transform 1 0 65520 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_577
timestamp 1669390400
transform 1 0 65968 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_579
timestamp 1669390400
transform 1 0 66192 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_582
timestamp 1669390400
transform 1 0 66528 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_586
timestamp 1669390400
transform 1 0 66976 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_602
timestamp 1669390400
transform 1 0 68768 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_618
timestamp 1669390400
transform 1 0 70560 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_622
timestamp 1669390400
transform 1 0 71008 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1669390400
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_641
timestamp 1669390400
transform 1 0 73136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_644
timestamp 1669390400
transform 1 0 73472 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_648
timestamp 1669390400
transform 1 0 73920 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_654
timestamp 1669390400
transform 1 0 74592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_670
timestamp 1669390400
transform 1 0 76384 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_686
timestamp 1669390400
transform 1 0 78176 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_17
timestamp 1669390400
transform 1 0 3248 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_33
timestamp 1669390400
transform 1 0 5040 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_47
timestamp 1669390400
transform 1 0 6608 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_55
timestamp 1669390400
transform 1 0 7504 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_63
timestamp 1669390400
transform 1 0 8400 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_67 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 8848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_99
timestamp 1669390400
transform 1 0 12432 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_103
timestamp 1669390400
transform 1 0 12880 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_124
timestamp 1669390400
transform 1 0 15232 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_148
timestamp 1669390400
transform 1 0 17920 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_166
timestamp 1669390400
transform 1 0 19936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_170
timestamp 1669390400
transform 1 0 20384 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_174
timestamp 1669390400
transform 1 0 20832 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_181
timestamp 1669390400
transform 1 0 21616 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_184
timestamp 1669390400
transform 1 0 21952 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_202
timestamp 1669390400
transform 1 0 23968 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_218
timestamp 1669390400
transform 1 0 25760 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_222
timestamp 1669390400
transform 1 0 26208 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_226
timestamp 1669390400
transform 1 0 26656 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_244
timestamp 1669390400
transform 1 0 28672 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_258
timestamp 1669390400
transform 1 0 30240 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_262
timestamp 1669390400
transform 1 0 30688 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_264
timestamp 1669390400
transform 1 0 30912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_267
timestamp 1669390400
transform 1 0 31248 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_299
timestamp 1669390400
transform 1 0 34832 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_315
timestamp 1669390400
transform 1 0 36624 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1669390400
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1669390400
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1669390400
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1669390400
transform 1 0 60368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1669390400
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_534
timestamp 1669390400
transform 1 0 61152 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_566
timestamp 1669390400
transform 1 0 64736 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_582
timestamp 1669390400
transform 1 0 66528 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_586
timestamp 1669390400
transform 1 0 66976 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_594
timestamp 1669390400
transform 1 0 67872 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_598
timestamp 1669390400
transform 1 0 68320 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1669390400
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_605
timestamp 1669390400
transform 1 0 69104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_620
timestamp 1669390400
transform 1 0 70784 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_654
timestamp 1669390400
transform 1 0 74592 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_670
timestamp 1669390400
transform 1 0 76384 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_676
timestamp 1669390400
transform 1 0 77056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_679
timestamp 1669390400
transform 1 0 77392 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_687
timestamp 1669390400
transform 1 0 78288 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_17
timestamp 1669390400
transform 1 0 3248 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_33
timestamp 1669390400
transform 1 0 5040 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_41
timestamp 1669390400
transform 1 0 5936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_51
timestamp 1669390400
transform 1 0 7056 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_59
timestamp 1669390400
transform 1 0 7952 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_61
timestamp 1669390400
transform 1 0 8176 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_68
timestamp 1669390400
transform 1 0 8960 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1669390400
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_150
timestamp 1669390400
transform 1 0 18144 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_182
timestamp 1669390400
transform 1 0 21728 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_198
timestamp 1669390400
transform 1 0 23520 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_206
timestamp 1669390400
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_210
timestamp 1669390400
transform 1 0 24864 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1669390400
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1669390400
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1669390400
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1669390400
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1669390400
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_563
timestamp 1669390400
transform 1 0 64400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1669390400
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_570
timestamp 1669390400
transform 1 0 65184 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_634
timestamp 1669390400
transform 1 0 72352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1669390400
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_641
timestamp 1669390400
transform 1 0 73136 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_649
timestamp 1669390400
transform 1 0 74032 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_651
timestamp 1669390400
transform 1 0 74256 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_654
timestamp 1669390400
transform 1 0 74592 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_670
timestamp 1669390400
transform 1 0 76384 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_686
timestamp 1669390400
transform 1 0 78176 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_17
timestamp 1669390400
transform 1 0 3248 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_33
timestamp 1669390400
transform 1 0 5040 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_53
timestamp 1669390400
transform 1 0 7280 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_57
timestamp 1669390400
transform 1 0 7728 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_65
timestamp 1669390400
transform 1 0 8624 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_67
timestamp 1669390400
transform 1 0 8848 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_74
timestamp 1669390400
transform 1 0 9632 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1669390400
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1669390400
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1669390400
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1669390400
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1669390400
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1669390400
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_534
timestamp 1669390400
transform 1 0 61152 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_598
timestamp 1669390400
transform 1 0 68320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1669390400
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_605
timestamp 1669390400
transform 1 0 69104 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_637
timestamp 1669390400
transform 1 0 72688 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_645
timestamp 1669390400
transform 1 0 73584 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_649
timestamp 1669390400
transform 1 0 74032 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_651
timestamp 1669390400
transform 1 0 74256 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_654
timestamp 1669390400
transform 1 0 74592 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_670
timestamp 1669390400
transform 1 0 76384 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_676
timestamp 1669390400
transform 1 0 77056 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_684
timestamp 1669390400
transform 1 0 77952 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_17
timestamp 1669390400
transform 1 0 3248 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_49
timestamp 1669390400
transform 1 0 6832 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_57
timestamp 1669390400
transform 1 0 7728 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_61
timestamp 1669390400
transform 1 0 8176 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_63
timestamp 1669390400
transform 1 0 8400 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_81
timestamp 1669390400
transform 1 0 10416 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_113
timestamp 1669390400
transform 1 0 14000 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_129
timestamp 1669390400
transform 1 0 15792 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1669390400
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1669390400
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1669390400
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1669390400
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1669390400
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1669390400
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_563
timestamp 1669390400
transform 1 0 64400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1669390400
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_570
timestamp 1669390400
transform 1 0 65184 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_634
timestamp 1669390400
transform 1 0 72352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1669390400
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_641
timestamp 1669390400
transform 1 0 73136 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_649
timestamp 1669390400
transform 1 0 74032 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_651
timestamp 1669390400
transform 1 0 74256 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_654
timestamp 1669390400
transform 1 0 74592 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_670
timestamp 1669390400
transform 1 0 76384 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_686
timestamp 1669390400
transform 1 0 78176 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_17
timestamp 1669390400
transform 1 0 3248 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_33
timestamp 1669390400
transform 1 0 5040 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_69
timestamp 1669390400
transform 1 0 9072 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_77
timestamp 1669390400
transform 1 0 9968 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_87
timestamp 1669390400
transform 1 0 11088 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_103
timestamp 1669390400
transform 1 0 12880 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1669390400
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1669390400
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1669390400
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1669390400
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1669390400
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1669390400
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1669390400
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_598
timestamp 1669390400
transform 1 0 68320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1669390400
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_605
timestamp 1669390400
transform 1 0 69104 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_637
timestamp 1669390400
transform 1 0 72688 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_645
timestamp 1669390400
transform 1 0 73584 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_649
timestamp 1669390400
transform 1 0 74032 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_651
timestamp 1669390400
transform 1 0 74256 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_654
timestamp 1669390400
transform 1 0 74592 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_670
timestamp 1669390400
transform 1 0 76384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_676
timestamp 1669390400
transform 1 0 77056 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_684
timestamp 1669390400
transform 1 0 77952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_17
timestamp 1669390400
transform 1 0 3248 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_49
timestamp 1669390400
transform 1 0 6832 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_65
timestamp 1669390400
transform 1 0 8624 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_69
timestamp 1669390400
transform 1 0 9072 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_83
timestamp 1669390400
transform 1 0 10640 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_85
timestamp 1669390400
transform 1 0 10864 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_92
timestamp 1669390400
transform 1 0 11648 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_124
timestamp 1669390400
transform 1 0 15232 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_140
timestamp 1669390400
transform 1 0 17024 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1669390400
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1669390400
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1669390400
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1669390400
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_563
timestamp 1669390400
transform 1 0 64400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1669390400
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1669390400
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1669390400
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1669390400
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_641
timestamp 1669390400
transform 1 0 73136 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_649
timestamp 1669390400
transform 1 0 74032 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_651
timestamp 1669390400
transform 1 0 74256 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_654
timestamp 1669390400
transform 1 0 74592 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_670
timestamp 1669390400
transform 1 0 76384 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_686
timestamp 1669390400
transform 1 0 78176 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_17
timestamp 1669390400
transform 1 0 3248 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_21
timestamp 1669390400
transform 1 0 3696 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_25
timestamp 1669390400
transform 1 0 4144 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_33
timestamp 1669390400
transform 1 0 5040 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_69
timestamp 1669390400
transform 1 0 9072 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_77
timestamp 1669390400
transform 1 0 9968 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_81
timestamp 1669390400
transform 1 0 10416 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_88
timestamp 1669390400
transform 1 0 11200 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_96
timestamp 1669390400
transform 1 0 12096 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_104
timestamp 1669390400
transform 1 0 12992 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_111
timestamp 1669390400
transform 1 0 13776 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_175
timestamp 1669390400
transform 1 0 20944 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1669390400
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1669390400
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1669390400
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1669390400
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1669390400
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1669390400
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_598
timestamp 1669390400
transform 1 0 68320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1669390400
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_605
timestamp 1669390400
transform 1 0 69104 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_637
timestamp 1669390400
transform 1 0 72688 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_645
timestamp 1669390400
transform 1 0 73584 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_649
timestamp 1669390400
transform 1 0 74032 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_651
timestamp 1669390400
transform 1 0 74256 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_654
timestamp 1669390400
transform 1 0 74592 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_670
timestamp 1669390400
transform 1 0 76384 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_676
timestamp 1669390400
transform 1 0 77056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_679
timestamp 1669390400
transform 1 0 77392 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_687
timestamp 1669390400
transform 1 0 78288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_17
timestamp 1669390400
transform 1 0 3248 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_33
timestamp 1669390400
transform 1 0 5040 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_65
timestamp 1669390400
transform 1 0 8624 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_69
timestamp 1669390400
transform 1 0 9072 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_81
timestamp 1669390400
transform 1 0 10416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_85
timestamp 1669390400
transform 1 0 10864 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_87
timestamp 1669390400
transform 1 0 11088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_94
timestamp 1669390400
transform 1 0 11872 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_102
timestamp 1669390400
transform 1 0 12768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_110
timestamp 1669390400
transform 1 0 13664 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_114
timestamp 1669390400
transform 1 0 14112 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_130
timestamp 1669390400
transform 1 0 15904 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_138
timestamp 1669390400
transform 1 0 16800 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1669390400
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1669390400
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1669390400
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1669390400
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_563
timestamp 1669390400
transform 1 0 64400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1669390400
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1669390400
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1669390400
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1669390400
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_641
timestamp 1669390400
transform 1 0 73136 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_649
timestamp 1669390400
transform 1 0 74032 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_651
timestamp 1669390400
transform 1 0 74256 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_654
timestamp 1669390400
transform 1 0 74592 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_670
timestamp 1669390400
transform 1 0 76384 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_686
timestamp 1669390400
transform 1 0 78176 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_17
timestamp 1669390400
transform 1 0 3248 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_21
timestamp 1669390400
transform 1 0 3696 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_29
timestamp 1669390400
transform 1 0 4592 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_33
timestamp 1669390400
transform 1 0 5040 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_69
timestamp 1669390400
transform 1 0 9072 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_85
timestamp 1669390400
transform 1 0 10864 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_93
timestamp 1669390400
transform 1 0 11760 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_96
timestamp 1669390400
transform 1 0 12096 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_100
timestamp 1669390400
transform 1 0 12544 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_104
timestamp 1669390400
transform 1 0 12992 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1669390400
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1669390400
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_481
timestamp 1669390400
transform 1 0 55216 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_513
timestamp 1669390400
transform 1 0 58800 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_529
timestamp 1669390400
transform 1 0 60592 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1669390400
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1669390400
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_598
timestamp 1669390400
transform 1 0 68320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1669390400
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_605
timestamp 1669390400
transform 1 0 69104 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_637
timestamp 1669390400
transform 1 0 72688 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_645
timestamp 1669390400
transform 1 0 73584 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_649
timestamp 1669390400
transform 1 0 74032 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_651
timestamp 1669390400
transform 1 0 74256 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_654
timestamp 1669390400
transform 1 0 74592 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_670
timestamp 1669390400
transform 1 0 76384 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_676
timestamp 1669390400
transform 1 0 77056 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_684
timestamp 1669390400
transform 1 0 77952 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_17
timestamp 1669390400
transform 1 0 3248 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_21
timestamp 1669390400
transform 1 0 3696 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_53
timestamp 1669390400
transform 1 0 7280 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_69
timestamp 1669390400
transform 1 0 9072 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_89
timestamp 1669390400
transform 1 0 11312 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_93
timestamp 1669390400
transform 1 0 11760 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_96
timestamp 1669390400
transform 1 0 12096 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_104
timestamp 1669390400
transform 1 0 12992 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_112
timestamp 1669390400
transform 1 0 13888 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_116
timestamp 1669390400
transform 1 0 14336 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_132
timestamp 1669390400
transform 1 0 16128 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_140
timestamp 1669390400
transform 1 0 17024 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1669390400
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1669390400
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1669390400
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1669390400
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_460
timestamp 1669390400
transform 1 0 52864 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_468
timestamp 1669390400
transform 1 0 53760 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_472
timestamp 1669390400
transform 1 0 54208 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_474
timestamp 1669390400
transform 1 0 54432 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_477
timestamp 1669390400
transform 1 0 54768 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_487
timestamp 1669390400
transform 1 0 55888 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_491
timestamp 1669390400
transform 1 0 56336 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_493
timestamp 1669390400
transform 1 0 56560 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1669390400
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_506
timestamp 1669390400
transform 1 0 58016 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_538
timestamp 1669390400
transform 1 0 61600 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_554
timestamp 1669390400
transform 1 0 63392 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_562
timestamp 1669390400
transform 1 0 64288 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_566
timestamp 1669390400
transform 1 0 64736 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1669390400
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1669390400
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1669390400
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_641
timestamp 1669390400
transform 1 0 73136 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_649
timestamp 1669390400
transform 1 0 74032 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_651
timestamp 1669390400
transform 1 0 74256 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_654
timestamp 1669390400
transform 1 0 74592 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_670
timestamp 1669390400
transform 1 0 76384 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_686
timestamp 1669390400
transform 1 0 78176 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_17
timestamp 1669390400
transform 1 0 3248 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_21
timestamp 1669390400
transform 1 0 3696 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_29
timestamp 1669390400
transform 1 0 4592 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_33
timestamp 1669390400
transform 1 0 5040 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_118
timestamp 1669390400
transform 1 0 14560 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_122
timestamp 1669390400
transform 1 0 15008 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_154
timestamp 1669390400
transform 1 0 18592 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_170
timestamp 1669390400
transform 1 0 20384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_174
timestamp 1669390400
transform 1 0 20832 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1669390400
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1669390400
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1669390400
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1669390400
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_469
timestamp 1669390400
transform 1 0 53872 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_473
timestamp 1669390400
transform 1 0 54320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_485
timestamp 1669390400
transform 1 0 55664 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_493
timestamp 1669390400
transform 1 0 56560 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_497
timestamp 1669390400
transform 1 0 57008 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_529
timestamp 1669390400
transform 1 0 60592 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1669390400
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1669390400
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1669390400
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1669390400
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_605
timestamp 1669390400
transform 1 0 69104 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_637
timestamp 1669390400
transform 1 0 72688 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_645
timestamp 1669390400
transform 1 0 73584 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_649
timestamp 1669390400
transform 1 0 74032 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_651
timestamp 1669390400
transform 1 0 74256 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_654
timestamp 1669390400
transform 1 0 74592 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_670
timestamp 1669390400
transform 1 0 76384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_676
timestamp 1669390400
transform 1 0 77056 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_684
timestamp 1669390400
transform 1 0 77952 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_17
timestamp 1669390400
transform 1 0 3248 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_21
timestamp 1669390400
transform 1 0 3696 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_53
timestamp 1669390400
transform 1 0 7280 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_69
timestamp 1669390400
transform 1 0 9072 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_105
timestamp 1669390400
transform 1 0 13104 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_113
timestamp 1669390400
transform 1 0 14000 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_117
timestamp 1669390400
transform 1 0 14448 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_124
timestamp 1669390400
transform 1 0 15232 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_128
timestamp 1669390400
transform 1 0 15680 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_132
timestamp 1669390400
transform 1 0 16128 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_136
timestamp 1669390400
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_140
timestamp 1669390400
transform 1 0 17024 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_148
timestamp 1669390400
transform 1 0 17920 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_152
timestamp 1669390400
transform 1 0 18368 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_156
timestamp 1669390400
transform 1 0 18816 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_160
timestamp 1669390400
transform 1 0 19264 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_192
timestamp 1669390400
transform 1 0 22848 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1669390400
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_460
timestamp 1669390400
transform 1 0 52864 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_476
timestamp 1669390400
transform 1 0 54656 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_480
timestamp 1669390400
transform 1 0 55104 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_482
timestamp 1669390400
transform 1 0 55328 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_485
timestamp 1669390400
transform 1 0 55664 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_493
timestamp 1669390400
transform 1 0 56560 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1669390400
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1669390400
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1669390400
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1669390400
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1669390400
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_641
timestamp 1669390400
transform 1 0 73136 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_649
timestamp 1669390400
transform 1 0 74032 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_651
timestamp 1669390400
transform 1 0 74256 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_654
timestamp 1669390400
transform 1 0 74592 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_670
timestamp 1669390400
transform 1 0 76384 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_686
timestamp 1669390400
transform 1 0 78176 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_17
timestamp 1669390400
transform 1 0 3248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_21
timestamp 1669390400
transform 1 0 3696 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_25
timestamp 1669390400
transform 1 0 4144 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_33
timestamp 1669390400
transform 1 0 5040 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_124
timestamp 1669390400
transform 1 0 15232 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_134
timestamp 1669390400
transform 1 0 16352 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_136
timestamp 1669390400
transform 1 0 16576 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_139
timestamp 1669390400
transform 1 0 16912 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_143
timestamp 1669390400
transform 1 0 17360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_147
timestamp 1669390400
transform 1 0 17808 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_158
timestamp 1669390400
transform 1 0 19040 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_166
timestamp 1669390400
transform 1 0 19936 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_170
timestamp 1669390400
transform 1 0 20384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_174
timestamp 1669390400
transform 1 0 20832 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_187
timestamp 1669390400
transform 1 0 22288 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_197
timestamp 1669390400
transform 1 0 23408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_203
timestamp 1669390400
transform 1 0 24080 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_207
timestamp 1669390400
transform 1 0 24528 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_239
timestamp 1669390400
transform 1 0 28112 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1669390400
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1669390400
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1669390400
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1669390400
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1669390400
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1669390400
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_598
timestamp 1669390400
transform 1 0 68320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1669390400
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_605
timestamp 1669390400
transform 1 0 69104 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_637
timestamp 1669390400
transform 1 0 72688 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_645
timestamp 1669390400
transform 1 0 73584 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_649
timestamp 1669390400
transform 1 0 74032 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_651
timestamp 1669390400
transform 1 0 74256 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_654
timestamp 1669390400
transform 1 0 74592 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_670
timestamp 1669390400
transform 1 0 76384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_676
timestamp 1669390400
transform 1 0 77056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_679
timestamp 1669390400
transform 1 0 77392 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_687
timestamp 1669390400
transform 1 0 78288 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_17
timestamp 1669390400
transform 1 0 3248 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_33
timestamp 1669390400
transform 1 0 5040 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_37
timestamp 1669390400
transform 1 0 5488 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_69
timestamp 1669390400
transform 1 0 9072 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_105
timestamp 1669390400
transform 1 0 13104 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_121
timestamp 1669390400
transform 1 0 14896 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_125
timestamp 1669390400
transform 1 0 15344 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_133
timestamp 1669390400
transform 1 0 16240 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_147
timestamp 1669390400
transform 1 0 17808 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_155
timestamp 1669390400
transform 1 0 18704 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_157
timestamp 1669390400
transform 1 0 18928 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_164
timestamp 1669390400
transform 1 0 19712 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_168
timestamp 1669390400
transform 1 0 20160 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_172
timestamp 1669390400
transform 1 0 20608 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_178
timestamp 1669390400
transform 1 0 21280 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_186
timestamp 1669390400
transform 1 0 22176 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_189
timestamp 1669390400
transform 1 0 22512 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_201
timestamp 1669390400
transform 1 0 23856 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_205
timestamp 1669390400
transform 1 0 24304 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_208
timestamp 1669390400
transform 1 0 24640 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_227
timestamp 1669390400
transform 1 0 26768 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_259
timestamp 1669390400
transform 1 0 30352 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_275
timestamp 1669390400
transform 1 0 32144 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1669390400
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1669390400
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_460
timestamp 1669390400
transform 1 0 52864 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_468
timestamp 1669390400
transform 1 0 53760 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_472
timestamp 1669390400
transform 1 0 54208 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_474
timestamp 1669390400
transform 1 0 54432 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_477
timestamp 1669390400
transform 1 0 54768 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_493
timestamp 1669390400
transform 1 0 56560 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_563
timestamp 1669390400
transform 1 0 64400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1669390400
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1669390400
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_634
timestamp 1669390400
transform 1 0 72352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1669390400
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_641
timestamp 1669390400
transform 1 0 73136 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_649
timestamp 1669390400
transform 1 0 74032 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_651
timestamp 1669390400
transform 1 0 74256 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_654
timestamp 1669390400
transform 1 0 74592 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_670
timestamp 1669390400
transform 1 0 76384 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_686
timestamp 1669390400
transform 1 0 78176 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_17
timestamp 1669390400
transform 1 0 3248 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_21
timestamp 1669390400
transform 1 0 3696 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_29
timestamp 1669390400
transform 1 0 4592 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_33
timestamp 1669390400
transform 1 0 5040 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_124
timestamp 1669390400
transform 1 0 15232 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_132
timestamp 1669390400
transform 1 0 16128 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_135
timestamp 1669390400
transform 1 0 16464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_139
timestamp 1669390400
transform 1 0 16912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_142
timestamp 1669390400
transform 1 0 17248 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_150
timestamp 1669390400
transform 1 0 18144 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_158
timestamp 1669390400
transform 1 0 19040 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_162
timestamp 1669390400
transform 1 0 19488 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_182
timestamp 1669390400
transform 1 0 21728 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_186
timestamp 1669390400
transform 1 0 22176 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_202
timestamp 1669390400
transform 1 0 23968 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_205
timestamp 1669390400
transform 1 0 24304 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_209
timestamp 1669390400
transform 1 0 24752 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_212
timestamp 1669390400
transform 1 0 25088 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_216
timestamp 1669390400
transform 1 0 25536 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_224
timestamp 1669390400
transform 1 0 26432 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_240
timestamp 1669390400
transform 1 0 28224 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1669390400
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1669390400
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_469
timestamp 1669390400
transform 1 0 53872 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_473
timestamp 1669390400
transform 1 0 54320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_486
timestamp 1669390400
transform 1 0 55776 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_492
timestamp 1669390400
transform 1 0 56448 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_496
timestamp 1669390400
transform 1 0 56896 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_528
timestamp 1669390400
transform 1 0 60480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1669390400
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_598
timestamp 1669390400
transform 1 0 68320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1669390400
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_605
timestamp 1669390400
transform 1 0 69104 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_637
timestamp 1669390400
transform 1 0 72688 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_645
timestamp 1669390400
transform 1 0 73584 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_649
timestamp 1669390400
transform 1 0 74032 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_651
timestamp 1669390400
transform 1 0 74256 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_654
timestamp 1669390400
transform 1 0 74592 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_670
timestamp 1669390400
transform 1 0 76384 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_676
timestamp 1669390400
transform 1 0 77056 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_684
timestamp 1669390400
transform 1 0 77952 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_17
timestamp 1669390400
transform 1 0 3248 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_21
timestamp 1669390400
transform 1 0 3696 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_53
timestamp 1669390400
transform 1 0 7280 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_69
timestamp 1669390400
transform 1 0 9072 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1669390400
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_148
timestamp 1669390400
transform 1 0 17920 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_151
timestamp 1669390400
transform 1 0 18256 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_159
timestamp 1669390400
transform 1 0 19152 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_163
timestamp 1669390400
transform 1 0 19600 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_166
timestamp 1669390400
transform 1 0 19936 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_170
timestamp 1669390400
transform 1 0 20384 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_178
timestamp 1669390400
transform 1 0 21280 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_182
timestamp 1669390400
transform 1 0 21728 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_198
timestamp 1669390400
transform 1 0 23520 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_206
timestamp 1669390400
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_210
timestamp 1669390400
transform 1 0 24864 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1669390400
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_460
timestamp 1669390400
transform 1 0 52864 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_468
timestamp 1669390400
transform 1 0 53760 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_472
timestamp 1669390400
transform 1 0 54208 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_474
timestamp 1669390400
transform 1 0 54432 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_477
timestamp 1669390400
transform 1 0 54768 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_481
timestamp 1669390400
transform 1 0 55216 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1669390400
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_563
timestamp 1669390400
transform 1 0 64400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1669390400
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1669390400
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1669390400
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1669390400
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_641
timestamp 1669390400
transform 1 0 73136 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_649
timestamp 1669390400
transform 1 0 74032 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_651
timestamp 1669390400
transform 1 0 74256 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_654
timestamp 1669390400
transform 1 0 74592 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_670
timestamp 1669390400
transform 1 0 76384 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_686
timestamp 1669390400
transform 1 0 78176 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_17
timestamp 1669390400
transform 1 0 3248 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_21
timestamp 1669390400
transform 1 0 3696 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_29
timestamp 1669390400
transform 1 0 4592 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_33
timestamp 1669390400
transform 1 0 5040 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_140
timestamp 1669390400
transform 1 0 17024 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_148
timestamp 1669390400
transform 1 0 17920 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_152
timestamp 1669390400
transform 1 0 18368 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_160
timestamp 1669390400
transform 1 0 19264 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_168
timestamp 1669390400
transform 1 0 20160 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_186
timestamp 1669390400
transform 1 0 22176 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_190
timestamp 1669390400
transform 1 0 22624 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_222
timestamp 1669390400
transform 1 0 26208 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_238
timestamp 1669390400
transform 1 0 28000 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_246
timestamp 1669390400
transform 1 0 28896 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1669390400
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1669390400
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_527
timestamp 1669390400
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1669390400
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1669390400
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_598
timestamp 1669390400
transform 1 0 68320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1669390400
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_605
timestamp 1669390400
transform 1 0 69104 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_637
timestamp 1669390400
transform 1 0 72688 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_645
timestamp 1669390400
transform 1 0 73584 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_649
timestamp 1669390400
transform 1 0 74032 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_651
timestamp 1669390400
transform 1 0 74256 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_654
timestamp 1669390400
transform 1 0 74592 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_670
timestamp 1669390400
transform 1 0 76384 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_676
timestamp 1669390400
transform 1 0 77056 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_684
timestamp 1669390400
transform 1 0 77952 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_17
timestamp 1669390400
transform 1 0 3248 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_21
timestamp 1669390400
transform 1 0 3696 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_53
timestamp 1669390400
transform 1 0 7280 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_69
timestamp 1669390400
transform 1 0 9072 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_160
timestamp 1669390400
transform 1 0 19264 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_163
timestamp 1669390400
transform 1 0 19600 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_171
timestamp 1669390400
transform 1 0 20496 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_179
timestamp 1669390400
transform 1 0 21392 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_183
timestamp 1669390400
transform 1 0 21840 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_199
timestamp 1669390400
transform 1 0 23632 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_207
timestamp 1669390400
transform 1 0 24528 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_211
timestamp 1669390400
transform 1 0 24976 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1669390400
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1669390400
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1669390400
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1669390400
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_563
timestamp 1669390400
transform 1 0 64400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1669390400
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1669390400
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_634
timestamp 1669390400
transform 1 0 72352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1669390400
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_641
timestamp 1669390400
transform 1 0 73136 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_649
timestamp 1669390400
transform 1 0 74032 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_651
timestamp 1669390400
transform 1 0 74256 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_654
timestamp 1669390400
transform 1 0 74592 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_670
timestamp 1669390400
transform 1 0 76384 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_686
timestamp 1669390400
transform 1 0 78176 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_17
timestamp 1669390400
transform 1 0 3248 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_21
timestamp 1669390400
transform 1 0 3696 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_25
timestamp 1669390400
transform 1 0 4144 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_33
timestamp 1669390400
transform 1 0 5040 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_186
timestamp 1669390400
transform 1 0 22176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_192
timestamp 1669390400
transform 1 0 22848 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_200
timestamp 1669390400
transform 1 0 23744 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_232
timestamp 1669390400
transform 1 0 27328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1669390400
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1669390400
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_527
timestamp 1669390400
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1669390400
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1669390400
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_598
timestamp 1669390400
transform 1 0 68320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1669390400
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_605
timestamp 1669390400
transform 1 0 69104 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_637
timestamp 1669390400
transform 1 0 72688 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_645
timestamp 1669390400
transform 1 0 73584 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_649
timestamp 1669390400
transform 1 0 74032 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_651
timestamp 1669390400
transform 1 0 74256 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_654
timestamp 1669390400
transform 1 0 74592 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_670
timestamp 1669390400
transform 1 0 76384 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_676
timestamp 1669390400
transform 1 0 77056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_679
timestamp 1669390400
transform 1 0 77392 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_687
timestamp 1669390400
transform 1 0 78288 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_17
timestamp 1669390400
transform 1 0 3248 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_33
timestamp 1669390400
transform 1 0 5040 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_37
timestamp 1669390400
transform 1 0 5488 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_69
timestamp 1669390400
transform 1 0 9072 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_176
timestamp 1669390400
transform 1 0 21056 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_180
timestamp 1669390400
transform 1 0 21504 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_187
timestamp 1669390400
transform 1 0 22288 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_189
timestamp 1669390400
transform 1 0 22512 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_192
timestamp 1669390400
transform 1 0 22848 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_196
timestamp 1669390400
transform 1 0 23296 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_204
timestamp 1669390400
transform 1 0 24192 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1669390400
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1669390400
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1669390400
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_563
timestamp 1669390400
transform 1 0 64400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1669390400
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1669390400
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_634
timestamp 1669390400
transform 1 0 72352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1669390400
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_641
timestamp 1669390400
transform 1 0 73136 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_649
timestamp 1669390400
transform 1 0 74032 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_651
timestamp 1669390400
transform 1 0 74256 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_654
timestamp 1669390400
transform 1 0 74592 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_670
timestamp 1669390400
transform 1 0 76384 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_686
timestamp 1669390400
transform 1 0 78176 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_17
timestamp 1669390400
transform 1 0 3248 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_21
timestamp 1669390400
transform 1 0 3696 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_29
timestamp 1669390400
transform 1 0 4592 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_33
timestamp 1669390400
transform 1 0 5040 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1669390400
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_183
timestamp 1669390400
transform 1 0 21840 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_190
timestamp 1669390400
transform 1 0 22624 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_198
timestamp 1669390400
transform 1 0 23520 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_202
timestamp 1669390400
transform 1 0 23968 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_206
timestamp 1669390400
transform 1 0 24416 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_238
timestamp 1669390400
transform 1 0 28000 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_246
timestamp 1669390400
transform 1 0 28896 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1669390400
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1669390400
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1669390400
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_527
timestamp 1669390400
transform 1 0 60368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1669390400
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1669390400
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_598
timestamp 1669390400
transform 1 0 68320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1669390400
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_605
timestamp 1669390400
transform 1 0 69104 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_637
timestamp 1669390400
transform 1 0 72688 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_645
timestamp 1669390400
transform 1 0 73584 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_649
timestamp 1669390400
transform 1 0 74032 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_651
timestamp 1669390400
transform 1 0 74256 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_654
timestamp 1669390400
transform 1 0 74592 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_670
timestamp 1669390400
transform 1 0 76384 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_676
timestamp 1669390400
transform 1 0 77056 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_684
timestamp 1669390400
transform 1 0 77952 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_17
timestamp 1669390400
transform 1 0 3248 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_21
timestamp 1669390400
transform 1 0 3696 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_53
timestamp 1669390400
transform 1 0 7280 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_69
timestamp 1669390400
transform 1 0 9072 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_176
timestamp 1669390400
transform 1 0 21056 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_184
timestamp 1669390400
transform 1 0 21952 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_186
timestamp 1669390400
transform 1 0 22176 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_193
timestamp 1669390400
transform 1 0 22960 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_203
timestamp 1669390400
transform 1 0 24080 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_207
timestamp 1669390400
transform 1 0 24528 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_211
timestamp 1669390400
transform 1 0 24976 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1669390400
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1669390400
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1669390400
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_563
timestamp 1669390400
transform 1 0 64400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1669390400
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1669390400
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1669390400
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1669390400
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_641
timestamp 1669390400
transform 1 0 73136 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_649
timestamp 1669390400
transform 1 0 74032 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_651
timestamp 1669390400
transform 1 0 74256 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_654
timestamp 1669390400
transform 1 0 74592 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_670
timestamp 1669390400
transform 1 0 76384 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_686
timestamp 1669390400
transform 1 0 78176 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_17
timestamp 1669390400
transform 1 0 3248 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_21
timestamp 1669390400
transform 1 0 3696 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_29
timestamp 1669390400
transform 1 0 4592 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_33
timestamp 1669390400
transform 1 0 5040 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1669390400
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_187
timestamp 1669390400
transform 1 0 22288 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_191
timestamp 1669390400
transform 1 0 22736 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_195
timestamp 1669390400
transform 1 0 23184 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_197
timestamp 1669390400
transform 1 0 23408 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_204
timestamp 1669390400
transform 1 0 24192 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_208
timestamp 1669390400
transform 1 0 24640 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_211
timestamp 1669390400
transform 1 0 24976 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_219
timestamp 1669390400
transform 1 0 25872 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_223
timestamp 1669390400
transform 1 0 26320 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_239
timestamp 1669390400
transform 1 0 28112 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1669390400
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1669390400
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_527
timestamp 1669390400
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1669390400
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1669390400
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_598
timestamp 1669390400
transform 1 0 68320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1669390400
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_605
timestamp 1669390400
transform 1 0 69104 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_637
timestamp 1669390400
transform 1 0 72688 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_645
timestamp 1669390400
transform 1 0 73584 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_649
timestamp 1669390400
transform 1 0 74032 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_651
timestamp 1669390400
transform 1 0 74256 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_654
timestamp 1669390400
transform 1 0 74592 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_670
timestamp 1669390400
transform 1 0 76384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_676
timestamp 1669390400
transform 1 0 77056 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_684
timestamp 1669390400
transform 1 0 77952 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_17
timestamp 1669390400
transform 1 0 3248 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_21
timestamp 1669390400
transform 1 0 3696 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_53
timestamp 1669390400
transform 1 0 7280 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_69
timestamp 1669390400
transform 1 0 9072 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_176
timestamp 1669390400
transform 1 0 21056 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_184
timestamp 1669390400
transform 1 0 21952 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_188
timestamp 1669390400
transform 1 0 22400 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_192
timestamp 1669390400
transform 1 0 22848 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_196
timestamp 1669390400
transform 1 0 23296 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_204
timestamp 1669390400
transform 1 0 24192 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_223
timestamp 1669390400
transform 1 0 26320 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_227
timestamp 1669390400
transform 1 0 26768 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_259
timestamp 1669390400
transform 1 0 30352 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_275
timestamp 1669390400
transform 1 0 32144 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1669390400
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1669390400
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_563
timestamp 1669390400
transform 1 0 64400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1669390400
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1669390400
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1669390400
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1669390400
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_641
timestamp 1669390400
transform 1 0 73136 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_649
timestamp 1669390400
transform 1 0 74032 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_651
timestamp 1669390400
transform 1 0 74256 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_654
timestamp 1669390400
transform 1 0 74592 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_670
timestamp 1669390400
transform 1 0 76384 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_686
timestamp 1669390400
transform 1 0 78176 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_17
timestamp 1669390400
transform 1 0 3248 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_21
timestamp 1669390400
transform 1 0 3696 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_25
timestamp 1669390400
transform 1 0 4144 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_33
timestamp 1669390400
transform 1 0 5040 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_195
timestamp 1669390400
transform 1 0 23184 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_203
timestamp 1669390400
transform 1 0 24080 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_210
timestamp 1669390400
transform 1 0 24864 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_218
timestamp 1669390400
transform 1 0 25760 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_228
timestamp 1669390400
transform 1 0 26880 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_232
timestamp 1669390400
transform 1 0 27328 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_236
timestamp 1669390400
transform 1 0 27776 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_244
timestamp 1669390400
transform 1 0 28672 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1669390400
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1669390400
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_527
timestamp 1669390400
transform 1 0 60368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1669390400
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1669390400
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1669390400
transform 1 0 68320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1669390400
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_605
timestamp 1669390400
transform 1 0 69104 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_637
timestamp 1669390400
transform 1 0 72688 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_645
timestamp 1669390400
transform 1 0 73584 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_649
timestamp 1669390400
transform 1 0 74032 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_651
timestamp 1669390400
transform 1 0 74256 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_654
timestamp 1669390400
transform 1 0 74592 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_670
timestamp 1669390400
transform 1 0 76384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_676
timestamp 1669390400
transform 1 0 77056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_679
timestamp 1669390400
transform 1 0 77392 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_687
timestamp 1669390400
transform 1 0 78288 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_17
timestamp 1669390400
transform 1 0 3248 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_33
timestamp 1669390400
transform 1 0 5040 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_37
timestamp 1669390400
transform 1 0 5488 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_69
timestamp 1669390400
transform 1 0 9072 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_219
timestamp 1669390400
transform 1 0 25872 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_227
timestamp 1669390400
transform 1 0 26768 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_237
timestamp 1669390400
transform 1 0 27888 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_269
timestamp 1669390400
transform 1 0 31472 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_277
timestamp 1669390400
transform 1 0 32368 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_281
timestamp 1669390400
transform 1 0 32816 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1669390400
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1669390400
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1669390400
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_563
timestamp 1669390400
transform 1 0 64400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1669390400
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1669390400
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1669390400
transform 1 0 72352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1669390400
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_641
timestamp 1669390400
transform 1 0 73136 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_649
timestamp 1669390400
transform 1 0 74032 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_651
timestamp 1669390400
transform 1 0 74256 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_654
timestamp 1669390400
transform 1 0 74592 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_670
timestamp 1669390400
transform 1 0 76384 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_686
timestamp 1669390400
transform 1 0 78176 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_17
timestamp 1669390400
transform 1 0 3248 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_21
timestamp 1669390400
transform 1 0 3696 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_29
timestamp 1669390400
transform 1 0 4592 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_33
timestamp 1669390400
transform 1 0 5040 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_211
timestamp 1669390400
transform 1 0 24976 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_219
timestamp 1669390400
transform 1 0 25872 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_225
timestamp 1669390400
transform 1 0 26544 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_233
timestamp 1669390400
transform 1 0 27440 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_235
timestamp 1669390400
transform 1 0 27664 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_242
timestamp 1669390400
transform 1 0 28448 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_246
timestamp 1669390400
transform 1 0 28896 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1669390400
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1669390400
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1669390400
transform 1 0 60368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1669390400
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1669390400
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1669390400
transform 1 0 68320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1669390400
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_605
timestamp 1669390400
transform 1 0 69104 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_637
timestamp 1669390400
transform 1 0 72688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_645
timestamp 1669390400
transform 1 0 73584 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_649
timestamp 1669390400
transform 1 0 74032 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_651
timestamp 1669390400
transform 1 0 74256 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_654
timestamp 1669390400
transform 1 0 74592 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_670
timestamp 1669390400
transform 1 0 76384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_676
timestamp 1669390400
transform 1 0 77056 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_684
timestamp 1669390400
transform 1 0 77952 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_17
timestamp 1669390400
transform 1 0 3248 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_21
timestamp 1669390400
transform 1 0 3696 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_53
timestamp 1669390400
transform 1 0 7280 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_69
timestamp 1669390400
transform 1 0 9072 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_223
timestamp 1669390400
transform 1 0 26320 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_227
timestamp 1669390400
transform 1 0 26768 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_231
timestamp 1669390400
transform 1 0 27216 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_239
timestamp 1669390400
transform 1 0 28112 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_241
timestamp 1669390400
transform 1 0 28336 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_248
timestamp 1669390400
transform 1 0 29120 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_252
timestamp 1669390400
transform 1 0 29568 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_256
timestamp 1669390400
transform 1 0 30016 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_272
timestamp 1669390400
transform 1 0 31808 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_280
timestamp 1669390400
transform 1 0 32704 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1669390400
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1669390400
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1669390400
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1669390400
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1669390400
transform 1 0 64400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1669390400
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1669390400
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1669390400
transform 1 0 72352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1669390400
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_641
timestamp 1669390400
transform 1 0 73136 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_649
timestamp 1669390400
transform 1 0 74032 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_651
timestamp 1669390400
transform 1 0 74256 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_654
timestamp 1669390400
transform 1 0 74592 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_670
timestamp 1669390400
transform 1 0 76384 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_686
timestamp 1669390400
transform 1 0 78176 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_17
timestamp 1669390400
transform 1 0 3248 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_21
timestamp 1669390400
transform 1 0 3696 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_29
timestamp 1669390400
transform 1 0 4592 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_33
timestamp 1669390400
transform 1 0 5040 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_211
timestamp 1669390400
transform 1 0 24976 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_227
timestamp 1669390400
transform 1 0 26768 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_237
timestamp 1669390400
transform 1 0 27888 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_245
timestamp 1669390400
transform 1 0 28784 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_257
timestamp 1669390400
transform 1 0 30128 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_289
timestamp 1669390400
transform 1 0 33712 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_305
timestamp 1669390400
transform 1 0 35504 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_313
timestamp 1669390400
transform 1 0 36400 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_317
timestamp 1669390400
transform 1 0 36848 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1669390400
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1669390400
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1669390400
transform 1 0 60368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1669390400
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1669390400
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1669390400
transform 1 0 68320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1669390400
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_605
timestamp 1669390400
transform 1 0 69104 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_637
timestamp 1669390400
transform 1 0 72688 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_645
timestamp 1669390400
transform 1 0 73584 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_649
timestamp 1669390400
transform 1 0 74032 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_651
timestamp 1669390400
transform 1 0 74256 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_654
timestamp 1669390400
transform 1 0 74592 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_670
timestamp 1669390400
transform 1 0 76384 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_676
timestamp 1669390400
transform 1 0 77056 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_684
timestamp 1669390400
transform 1 0 77952 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_17
timestamp 1669390400
transform 1 0 3248 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_21
timestamp 1669390400
transform 1 0 3696 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_53
timestamp 1669390400
transform 1 0 7280 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_69
timestamp 1669390400
transform 1 0 9072 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_231
timestamp 1669390400
transform 1 0 27216 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_239
timestamp 1669390400
transform 1 0 28112 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_243
timestamp 1669390400
transform 1 0 28560 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_251
timestamp 1669390400
transform 1 0 29456 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_261
timestamp 1669390400
transform 1 0 30576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_267
timestamp 1669390400
transform 1 0 31248 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_271
timestamp 1669390400
transform 1 0 31696 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1669390400
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1669390400
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1669390400
transform 1 0 64400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1669390400
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1669390400
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1669390400
transform 1 0 72352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1669390400
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_641
timestamp 1669390400
transform 1 0 73136 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_649
timestamp 1669390400
transform 1 0 74032 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_651
timestamp 1669390400
transform 1 0 74256 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_654
timestamp 1669390400
transform 1 0 74592 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_670
timestamp 1669390400
transform 1 0 76384 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_686
timestamp 1669390400
transform 1 0 78176 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_17
timestamp 1669390400
transform 1 0 3248 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_21
timestamp 1669390400
transform 1 0 3696 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_25
timestamp 1669390400
transform 1 0 4144 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_33
timestamp 1669390400
transform 1 0 5040 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_257
timestamp 1669390400
transform 1 0 30128 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_265
timestamp 1669390400
transform 1 0 31024 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_273
timestamp 1669390400
transform 1 0 31920 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_277
timestamp 1669390400
transform 1 0 32368 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_309
timestamp 1669390400
transform 1 0 35952 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_317
timestamp 1669390400
transform 1 0 36848 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1669390400
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1669390400
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1669390400
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1669390400
transform 1 0 60368 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1669390400
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1669390400
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1669390400
transform 1 0 68320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1669390400
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_605
timestamp 1669390400
transform 1 0 69104 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_637
timestamp 1669390400
transform 1 0 72688 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_645
timestamp 1669390400
transform 1 0 73584 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_649
timestamp 1669390400
transform 1 0 74032 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_651
timestamp 1669390400
transform 1 0 74256 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_654
timestamp 1669390400
transform 1 0 74592 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_670
timestamp 1669390400
transform 1 0 76384 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_676
timestamp 1669390400
transform 1 0 77056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_679
timestamp 1669390400
transform 1 0 77392 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_687
timestamp 1669390400
transform 1 0 78288 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_17
timestamp 1669390400
transform 1 0 3248 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_33
timestamp 1669390400
transform 1 0 5040 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_37
timestamp 1669390400
transform 1 0 5488 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_69
timestamp 1669390400
transform 1 0 9072 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_247
timestamp 1669390400
transform 1 0 29008 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_251
timestamp 1669390400
transform 1 0 29456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_261
timestamp 1669390400
transform 1 0 30576 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_269
timestamp 1669390400
transform 1 0 31472 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_271
timestamp 1669390400
transform 1 0 31696 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_278
timestamp 1669390400
transform 1 0 32480 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_282
timestamp 1669390400
transform 1 0 32928 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1669390400
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1669390400
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1669390400
transform 1 0 64400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1669390400
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1669390400
transform 1 0 65184 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1669390400
transform 1 0 72352 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1669390400
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_641
timestamp 1669390400
transform 1 0 73136 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_649
timestamp 1669390400
transform 1 0 74032 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_651
timestamp 1669390400
transform 1 0 74256 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_654
timestamp 1669390400
transform 1 0 74592 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_670
timestamp 1669390400
transform 1 0 76384 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_686
timestamp 1669390400
transform 1 0 78176 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_17
timestamp 1669390400
transform 1 0 3248 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_21
timestamp 1669390400
transform 1 0 3696 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_29
timestamp 1669390400
transform 1 0 4592 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_33
timestamp 1669390400
transform 1 0 5040 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_258
timestamp 1669390400
transform 1 0 30240 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_260
timestamp 1669390400
transform 1 0 30464 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_263
timestamp 1669390400
transform 1 0 30800 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_267
timestamp 1669390400
transform 1 0 31248 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_275
timestamp 1669390400
transform 1 0 32144 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_285
timestamp 1669390400
transform 1 0 33264 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_289
timestamp 1669390400
transform 1 0 33712 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_293
timestamp 1669390400
transform 1 0 34160 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_309
timestamp 1669390400
transform 1 0 35952 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_317
timestamp 1669390400
transform 1 0 36848 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1669390400
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1669390400
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1669390400
transform 1 0 60368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1669390400
transform 1 0 60816 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1669390400
transform 1 0 61152 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_598
timestamp 1669390400
transform 1 0 68320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1669390400
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_605
timestamp 1669390400
transform 1 0 69104 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_637
timestamp 1669390400
transform 1 0 72688 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_645
timestamp 1669390400
transform 1 0 73584 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_649
timestamp 1669390400
transform 1 0 74032 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_651
timestamp 1669390400
transform 1 0 74256 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_654
timestamp 1669390400
transform 1 0 74592 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_670
timestamp 1669390400
transform 1 0 76384 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_676
timestamp 1669390400
transform 1 0 77056 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_684
timestamp 1669390400
transform 1 0 77952 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_17
timestamp 1669390400
transform 1 0 3248 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_21
timestamp 1669390400
transform 1 0 3696 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_53
timestamp 1669390400
transform 1 0 7280 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_69
timestamp 1669390400
transform 1 0 9072 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_247
timestamp 1669390400
transform 1 0 29008 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_263
timestamp 1669390400
transform 1 0 30800 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_273
timestamp 1669390400
transform 1 0 31920 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_281
timestamp 1669390400
transform 1 0 32816 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_293
timestamp 1669390400
transform 1 0 34160 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_297
timestamp 1669390400
transform 1 0 34608 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_329
timestamp 1669390400
transform 1 0 38192 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_345
timestamp 1669390400
transform 1 0 39984 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_353
timestamp 1669390400
transform 1 0 40880 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1669390400
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1669390400
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1669390400
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1669390400
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_563
timestamp 1669390400
transform 1 0 64400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1669390400
transform 1 0 64848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1669390400
transform 1 0 65184 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_634
timestamp 1669390400
transform 1 0 72352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1669390400
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_641
timestamp 1669390400
transform 1 0 73136 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_649
timestamp 1669390400
transform 1 0 74032 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_651
timestamp 1669390400
transform 1 0 74256 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_654
timestamp 1669390400
transform 1 0 74592 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_670
timestamp 1669390400
transform 1 0 76384 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_686
timestamp 1669390400
transform 1 0 78176 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_17
timestamp 1669390400
transform 1 0 3248 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_21
timestamp 1669390400
transform 1 0 3696 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_29
timestamp 1669390400
transform 1 0 4592 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_33
timestamp 1669390400
transform 1 0 5040 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1669390400
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_266
timestamp 1669390400
transform 1 0 31136 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_274
timestamp 1669390400
transform 1 0 32032 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_276
timestamp 1669390400
transform 1 0 32256 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_279
timestamp 1669390400
transform 1 0 32592 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_287
timestamp 1669390400
transform 1 0 33488 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_297
timestamp 1669390400
transform 1 0 34608 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_301
timestamp 1669390400
transform 1 0 35056 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_317
timestamp 1669390400
transform 1 0 36848 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1669390400
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1669390400
transform 1 0 52416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_527
timestamp 1669390400
transform 1 0 60368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1669390400
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_534
timestamp 1669390400
transform 1 0 61152 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_598
timestamp 1669390400
transform 1 0 68320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1669390400
transform 1 0 68768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_605
timestamp 1669390400
transform 1 0 69104 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_637
timestamp 1669390400
transform 1 0 72688 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_645
timestamp 1669390400
transform 1 0 73584 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_649
timestamp 1669390400
transform 1 0 74032 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_651
timestamp 1669390400
transform 1 0 74256 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_654
timestamp 1669390400
transform 1 0 74592 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_670
timestamp 1669390400
transform 1 0 76384 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_676
timestamp 1669390400
transform 1 0 77056 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_684
timestamp 1669390400
transform 1 0 77952 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_17
timestamp 1669390400
transform 1 0 3248 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_21
timestamp 1669390400
transform 1 0 3696 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_53
timestamp 1669390400
transform 1 0 7280 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_69
timestamp 1669390400
transform 1 0 9072 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_294
timestamp 1669390400
transform 1 0 34272 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_296
timestamp 1669390400
transform 1 0 34496 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_303
timestamp 1669390400
transform 1 0 35280 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_309
timestamp 1669390400
transform 1 0 35952 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_313
timestamp 1669390400
transform 1 0 36400 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_345
timestamp 1669390400
transform 1 0 39984 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_353
timestamp 1669390400
transform 1 0 40880 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1669390400
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1669390400
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1669390400
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_563
timestamp 1669390400
transform 1 0 64400 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1669390400
transform 1 0 64848 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_570
timestamp 1669390400
transform 1 0 65184 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_634
timestamp 1669390400
transform 1 0 72352 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1669390400
transform 1 0 72800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_641
timestamp 1669390400
transform 1 0 73136 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_649
timestamp 1669390400
transform 1 0 74032 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_651
timestamp 1669390400
transform 1 0 74256 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_654
timestamp 1669390400
transform 1 0 74592 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_670
timestamp 1669390400
transform 1 0 76384 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_686
timestamp 1669390400
transform 1 0 78176 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_17
timestamp 1669390400
transform 1 0 3248 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_21
timestamp 1669390400
transform 1 0 3696 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_25
timestamp 1669390400
transform 1 0 4144 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_33
timestamp 1669390400
transform 1 0 5040 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_282
timestamp 1669390400
transform 1 0 32928 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_286
timestamp 1669390400
transform 1 0 33376 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_288
timestamp 1669390400
transform 1 0 33600 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_291
timestamp 1669390400
transform 1 0 33936 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_299
timestamp 1669390400
transform 1 0 34832 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_307
timestamp 1669390400
transform 1 0 35728 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_315
timestamp 1669390400
transform 1 0 36624 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_324
timestamp 1669390400
transform 1 0 37632 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_388
timestamp 1669390400
transform 1 0 44800 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1669390400
transform 1 0 52416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1669390400
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_527
timestamp 1669390400
transform 1 0 60368 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1669390400
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_534
timestamp 1669390400
transform 1 0 61152 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_598
timestamp 1669390400
transform 1 0 68320 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1669390400
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_605
timestamp 1669390400
transform 1 0 69104 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_637
timestamp 1669390400
transform 1 0 72688 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_645
timestamp 1669390400
transform 1 0 73584 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_649
timestamp 1669390400
transform 1 0 74032 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_651
timestamp 1669390400
transform 1 0 74256 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_654
timestamp 1669390400
transform 1 0 74592 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_670
timestamp 1669390400
transform 1 0 76384 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_676
timestamp 1669390400
transform 1 0 77056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_679
timestamp 1669390400
transform 1 0 77392 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_687
timestamp 1669390400
transform 1 0 78288 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_17
timestamp 1669390400
transform 1 0 3248 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_33
timestamp 1669390400
transform 1 0 5040 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_37
timestamp 1669390400
transform 1 0 5488 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_69
timestamp 1669390400
transform 1 0 9072 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1669390400
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1669390400
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_294
timestamp 1669390400
transform 1 0 34272 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_296
timestamp 1669390400
transform 1 0 34496 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_303
timestamp 1669390400
transform 1 0 35280 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_311
timestamp 1669390400
transform 1 0 36176 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_313
timestamp 1669390400
transform 1 0 36400 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_320
timestamp 1669390400
transform 1 0 37184 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_324
timestamp 1669390400
transform 1 0 37632 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_328
timestamp 1669390400
transform 1 0 38080 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_332
timestamp 1669390400
transform 1 0 38528 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_348
timestamp 1669390400
transform 1 0 40320 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_352
timestamp 1669390400
transform 1 0 40768 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1669390400
transform 1 0 48496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1669390400
transform 1 0 56448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1669390400
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_563
timestamp 1669390400
transform 1 0 64400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1669390400
transform 1 0 64848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_570
timestamp 1669390400
transform 1 0 65184 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_634
timestamp 1669390400
transform 1 0 72352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1669390400
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_641
timestamp 1669390400
transform 1 0 73136 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_649
timestamp 1669390400
transform 1 0 74032 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_651
timestamp 1669390400
transform 1 0 74256 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_654
timestamp 1669390400
transform 1 0 74592 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_670
timestamp 1669390400
transform 1 0 76384 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_686
timestamp 1669390400
transform 1 0 78176 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_17
timestamp 1669390400
transform 1 0 3248 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_21
timestamp 1669390400
transform 1 0 3696 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_29
timestamp 1669390400
transform 1 0 4592 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_33
timestamp 1669390400
transform 1 0 5040 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1669390400
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_282
timestamp 1669390400
transform 1 0 32928 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_298
timestamp 1669390400
transform 1 0 34720 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_302
timestamp 1669390400
transform 1 0 35168 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_305
timestamp 1669390400
transform 1 0 35504 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_309
timestamp 1669390400
transform 1 0 35952 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_317
timestamp 1669390400
transform 1 0 36848 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_328
timestamp 1669390400
transform 1 0 38080 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_360
timestamp 1669390400
transform 1 0 41664 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_376
timestamp 1669390400
transform 1 0 43456 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_384
timestamp 1669390400
transform 1 0 44352 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_388
timestamp 1669390400
transform 1 0 44800 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_456
timestamp 1669390400
transform 1 0 52416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1669390400
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_527
timestamp 1669390400
transform 1 0 60368 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_531
timestamp 1669390400
transform 1 0 60816 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_534
timestamp 1669390400
transform 1 0 61152 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_598
timestamp 1669390400
transform 1 0 68320 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_602
timestamp 1669390400
transform 1 0 68768 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_605
timestamp 1669390400
transform 1 0 69104 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_637
timestamp 1669390400
transform 1 0 72688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_645
timestamp 1669390400
transform 1 0 73584 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_649
timestamp 1669390400
transform 1 0 74032 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_651
timestamp 1669390400
transform 1 0 74256 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_654
timestamp 1669390400
transform 1 0 74592 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_670
timestamp 1669390400
transform 1 0 76384 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_676
timestamp 1669390400
transform 1 0 77056 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_684
timestamp 1669390400
transform 1 0 77952 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_17
timestamp 1669390400
transform 1 0 3248 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_21
timestamp 1669390400
transform 1 0 3696 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_53
timestamp 1669390400
transform 1 0 7280 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_69
timestamp 1669390400
transform 1 0 9072 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1669390400
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1669390400
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_302
timestamp 1669390400
transform 1 0 35168 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_310
timestamp 1669390400
transform 1 0 36064 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_312
timestamp 1669390400
transform 1 0 36288 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_315
timestamp 1669390400
transform 1 0 36624 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_323
timestamp 1669390400
transform 1 0 37520 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_333
timestamp 1669390400
transform 1 0 38640 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_337
timestamp 1669390400
transform 1 0 39088 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_341
timestamp 1669390400
transform 1 0 39536 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_349
timestamp 1669390400
transform 1 0 40432 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_353
timestamp 1669390400
transform 1 0 40880 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_421
timestamp 1669390400
transform 1 0 48496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1669390400
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_428
timestamp 1669390400
transform 1 0 49280 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_492
timestamp 1669390400
transform 1 0 56448 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_496
timestamp 1669390400
transform 1 0 56896 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_499
timestamp 1669390400
transform 1 0 57232 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_563
timestamp 1669390400
transform 1 0 64400 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_567
timestamp 1669390400
transform 1 0 64848 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_570
timestamp 1669390400
transform 1 0 65184 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_634
timestamp 1669390400
transform 1 0 72352 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_638
timestamp 1669390400
transform 1 0 72800 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_641
timestamp 1669390400
transform 1 0 73136 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_649
timestamp 1669390400
transform 1 0 74032 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_651
timestamp 1669390400
transform 1 0 74256 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_654
timestamp 1669390400
transform 1 0 74592 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_670
timestamp 1669390400
transform 1 0 76384 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_686
timestamp 1669390400
transform 1 0 78176 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_17
timestamp 1669390400
transform 1 0 3248 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_21
timestamp 1669390400
transform 1 0 3696 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_29
timestamp 1669390400
transform 1 0 4592 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_33
timestamp 1669390400
transform 1 0 5040 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1669390400
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1669390400
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1669390400
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1669390400
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_329
timestamp 1669390400
transform 1 0 38192 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_339
timestamp 1669390400
transform 1 0 39312 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_343
timestamp 1669390400
transform 1 0 39760 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_347
timestamp 1669390400
transform 1 0 40208 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_379
timestamp 1669390400
transform 1 0 43792 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_387
timestamp 1669390400
transform 1 0 44688 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1669390400
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_456
timestamp 1669390400
transform 1 0 52416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1669390400
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_463
timestamp 1669390400
transform 1 0 53200 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_527
timestamp 1669390400
transform 1 0 60368 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_531
timestamp 1669390400
transform 1 0 60816 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_534
timestamp 1669390400
transform 1 0 61152 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_598
timestamp 1669390400
transform 1 0 68320 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_602
timestamp 1669390400
transform 1 0 68768 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_605
timestamp 1669390400
transform 1 0 69104 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_637
timestamp 1669390400
transform 1 0 72688 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_645
timestamp 1669390400
transform 1 0 73584 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_649
timestamp 1669390400
transform 1 0 74032 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_651
timestamp 1669390400
transform 1 0 74256 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_654
timestamp 1669390400
transform 1 0 74592 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_670
timestamp 1669390400
transform 1 0 76384 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_676
timestamp 1669390400
transform 1 0 77056 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_684
timestamp 1669390400
transform 1 0 77952 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_17
timestamp 1669390400
transform 1 0 3248 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_21
timestamp 1669390400
transform 1 0 3696 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_53
timestamp 1669390400
transform 1 0 7280 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_69
timestamp 1669390400
transform 1 0 9072 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1669390400
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_318
timestamp 1669390400
transform 1 0 36960 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_322
timestamp 1669390400
transform 1 0 37408 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_324
timestamp 1669390400
transform 1 0 37632 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_327
timestamp 1669390400
transform 1 0 37968 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_335
timestamp 1669390400
transform 1 0 38864 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_337
timestamp 1669390400
transform 1 0 39088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_344
timestamp 1669390400
transform 1 0 39872 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1669390400
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_421
timestamp 1669390400
transform 1 0 48496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1669390400
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_428
timestamp 1669390400
transform 1 0 49280 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_492
timestamp 1669390400
transform 1 0 56448 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1669390400
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_499
timestamp 1669390400
transform 1 0 57232 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_563
timestamp 1669390400
transform 1 0 64400 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_567
timestamp 1669390400
transform 1 0 64848 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_570
timestamp 1669390400
transform 1 0 65184 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_634
timestamp 1669390400
transform 1 0 72352 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_638
timestamp 1669390400
transform 1 0 72800 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_641
timestamp 1669390400
transform 1 0 73136 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_649
timestamp 1669390400
transform 1 0 74032 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_651
timestamp 1669390400
transform 1 0 74256 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_654
timestamp 1669390400
transform 1 0 74592 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_670
timestamp 1669390400
transform 1 0 76384 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_686
timestamp 1669390400
transform 1 0 78176 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_17
timestamp 1669390400
transform 1 0 3248 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_21
timestamp 1669390400
transform 1 0 3696 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_29
timestamp 1669390400
transform 1 0 4592 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_33
timestamp 1669390400
transform 1 0 5040 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1669390400
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1669390400
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1669390400
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_329
timestamp 1669390400
transform 1 0 38192 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_332
timestamp 1669390400
transform 1 0 38528 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_340
timestamp 1669390400
transform 1 0 39424 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_348
timestamp 1669390400
transform 1 0 40320 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_356
timestamp 1669390400
transform 1 0 41216 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_360
timestamp 1669390400
transform 1 0 41664 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_376
timestamp 1669390400
transform 1 0 43456 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_384
timestamp 1669390400
transform 1 0 44352 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_388
timestamp 1669390400
transform 1 0 44800 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_456
timestamp 1669390400
transform 1 0 52416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_460
timestamp 1669390400
transform 1 0 52864 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_463
timestamp 1669390400
transform 1 0 53200 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_527
timestamp 1669390400
transform 1 0 60368 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_531
timestamp 1669390400
transform 1 0 60816 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_534
timestamp 1669390400
transform 1 0 61152 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_598
timestamp 1669390400
transform 1 0 68320 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_602
timestamp 1669390400
transform 1 0 68768 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_605
timestamp 1669390400
transform 1 0 69104 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_637
timestamp 1669390400
transform 1 0 72688 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_645
timestamp 1669390400
transform 1 0 73584 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_649
timestamp 1669390400
transform 1 0 74032 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_651
timestamp 1669390400
transform 1 0 74256 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_654
timestamp 1669390400
transform 1 0 74592 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_670
timestamp 1669390400
transform 1 0 76384 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_676
timestamp 1669390400
transform 1 0 77056 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_684
timestamp 1669390400
transform 1 0 77952 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_17
timestamp 1669390400
transform 1 0 3248 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_21
timestamp 1669390400
transform 1 0 3696 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_53
timestamp 1669390400
transform 1 0 7280 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_69
timestamp 1669390400
transform 1 0 9072 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1669390400
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1669390400
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1669390400
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1669390400
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1669390400
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_318
timestamp 1669390400
transform 1 0 36960 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_334
timestamp 1669390400
transform 1 0 38752 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_337
timestamp 1669390400
transform 1 0 39088 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_345
timestamp 1669390400
transform 1 0 39984 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_353
timestamp 1669390400
transform 1 0 40880 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_364
timestamp 1669390400
transform 1 0 42112 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_368
timestamp 1669390400
transform 1 0 42560 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_372
timestamp 1669390400
transform 1 0 43008 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_404
timestamp 1669390400
transform 1 0 46592 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_420
timestamp 1669390400
transform 1 0 48384 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_424
timestamp 1669390400
transform 1 0 48832 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_428
timestamp 1669390400
transform 1 0 49280 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_492
timestamp 1669390400
transform 1 0 56448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1669390400
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_499
timestamp 1669390400
transform 1 0 57232 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_563
timestamp 1669390400
transform 1 0 64400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_567
timestamp 1669390400
transform 1 0 64848 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_570
timestamp 1669390400
transform 1 0 65184 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_634
timestamp 1669390400
transform 1 0 72352 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_638
timestamp 1669390400
transform 1 0 72800 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_641
timestamp 1669390400
transform 1 0 73136 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_649
timestamp 1669390400
transform 1 0 74032 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_651
timestamp 1669390400
transform 1 0 74256 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_654
timestamp 1669390400
transform 1 0 74592 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_670
timestamp 1669390400
transform 1 0 76384 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_686
timestamp 1669390400
transform 1 0 78176 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_17
timestamp 1669390400
transform 1 0 3248 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_21
timestamp 1669390400
transform 1 0 3696 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_29
timestamp 1669390400
transform 1 0 4592 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_33
timestamp 1669390400
transform 1 0 5040 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1669390400
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1669390400
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1669390400
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1669390400
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1669390400
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1669390400
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_337
timestamp 1669390400
transform 1 0 39088 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_347
timestamp 1669390400
transform 1 0 40208 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_351
timestamp 1669390400
transform 1 0 40656 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_359
timestamp 1669390400
transform 1 0 41552 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_369
timestamp 1669390400
transform 1 0 42672 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_373
timestamp 1669390400
transform 1 0 43120 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1669390400
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_456
timestamp 1669390400
transform 1 0 52416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1669390400
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_463
timestamp 1669390400
transform 1 0 53200 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_527
timestamp 1669390400
transform 1 0 60368 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_531
timestamp 1669390400
transform 1 0 60816 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_534
timestamp 1669390400
transform 1 0 61152 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_598
timestamp 1669390400
transform 1 0 68320 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_602
timestamp 1669390400
transform 1 0 68768 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_605
timestamp 1669390400
transform 1 0 69104 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_637
timestamp 1669390400
transform 1 0 72688 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_645
timestamp 1669390400
transform 1 0 73584 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_649
timestamp 1669390400
transform 1 0 74032 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_651
timestamp 1669390400
transform 1 0 74256 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_654
timestamp 1669390400
transform 1 0 74592 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_670
timestamp 1669390400
transform 1 0 76384 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_676
timestamp 1669390400
transform 1 0 77056 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_684
timestamp 1669390400
transform 1 0 77952 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_17
timestamp 1669390400
transform 1 0 3248 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_21
timestamp 1669390400
transform 1 0 3696 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_53
timestamp 1669390400
transform 1 0 7280 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_69
timestamp 1669390400
transform 1 0 9072 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1669390400
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1669390400
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1669390400
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1669390400
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1669390400
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1669390400
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1669390400
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_359
timestamp 1669390400
transform 1 0 41552 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_366
timestamp 1669390400
transform 1 0 42336 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_368
timestamp 1669390400
transform 1 0 42560 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_375
timestamp 1669390400
transform 1 0 43344 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_379
timestamp 1669390400
transform 1 0 43792 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_411
timestamp 1669390400
transform 1 0 47376 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_419
timestamp 1669390400
transform 1 0 48272 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_423
timestamp 1669390400
transform 1 0 48720 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1669390400
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_428
timestamp 1669390400
transform 1 0 49280 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_492
timestamp 1669390400
transform 1 0 56448 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1669390400
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_499
timestamp 1669390400
transform 1 0 57232 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_563
timestamp 1669390400
transform 1 0 64400 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_567
timestamp 1669390400
transform 1 0 64848 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_570
timestamp 1669390400
transform 1 0 65184 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_634
timestamp 1669390400
transform 1 0 72352 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_638
timestamp 1669390400
transform 1 0 72800 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_641
timestamp 1669390400
transform 1 0 73136 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_649
timestamp 1669390400
transform 1 0 74032 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_651
timestamp 1669390400
transform 1 0 74256 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_654
timestamp 1669390400
transform 1 0 74592 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_670
timestamp 1669390400
transform 1 0 76384 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_686
timestamp 1669390400
transform 1 0 78176 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_17
timestamp 1669390400
transform 1 0 3248 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_21
timestamp 1669390400
transform 1 0 3696 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_29
timestamp 1669390400
transform 1 0 4592 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_33
timestamp 1669390400
transform 1 0 5040 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1669390400
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1669390400
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1669390400
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1669390400
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1669390400
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_353
timestamp 1669390400
transform 1 0 40880 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_363
timestamp 1669390400
transform 1 0 42000 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_371
timestamp 1669390400
transform 1 0 42896 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_373
timestamp 1669390400
transform 1 0 43120 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_380
timestamp 1669390400
transform 1 0 43904 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_384
timestamp 1669390400
transform 1 0 44352 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_388
timestamp 1669390400
transform 1 0 44800 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_456
timestamp 1669390400
transform 1 0 52416 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_460
timestamp 1669390400
transform 1 0 52864 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_463
timestamp 1669390400
transform 1 0 53200 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_527
timestamp 1669390400
transform 1 0 60368 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_531
timestamp 1669390400
transform 1 0 60816 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_534
timestamp 1669390400
transform 1 0 61152 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_598
timestamp 1669390400
transform 1 0 68320 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_602
timestamp 1669390400
transform 1 0 68768 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_605
timestamp 1669390400
transform 1 0 69104 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_637
timestamp 1669390400
transform 1 0 72688 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_645
timestamp 1669390400
transform 1 0 73584 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_649
timestamp 1669390400
transform 1 0 74032 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_651
timestamp 1669390400
transform 1 0 74256 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_654
timestamp 1669390400
transform 1 0 74592 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_670
timestamp 1669390400
transform 1 0 76384 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_676
timestamp 1669390400
transform 1 0 77056 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_684
timestamp 1669390400
transform 1 0 77952 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_17
timestamp 1669390400
transform 1 0 3248 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_21
timestamp 1669390400
transform 1 0 3696 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_53
timestamp 1669390400
transform 1 0 7280 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_69
timestamp 1669390400
transform 1 0 9072 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1669390400
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1669390400
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1669390400
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1669390400
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1669390400
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1669390400
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1669390400
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_365
timestamp 1669390400
transform 1 0 42224 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_369
timestamp 1669390400
transform 1 0 42672 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_377
timestamp 1669390400
transform 1 0 43568 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_387
timestamp 1669390400
transform 1 0 44688 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_391
timestamp 1669390400
transform 1 0 45136 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_423
timestamp 1669390400
transform 1 0 48720 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1669390400
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_428
timestamp 1669390400
transform 1 0 49280 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_492
timestamp 1669390400
transform 1 0 56448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1669390400
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_499
timestamp 1669390400
transform 1 0 57232 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_563
timestamp 1669390400
transform 1 0 64400 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_567
timestamp 1669390400
transform 1 0 64848 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_570
timestamp 1669390400
transform 1 0 65184 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_634
timestamp 1669390400
transform 1 0 72352 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_638
timestamp 1669390400
transform 1 0 72800 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_641
timestamp 1669390400
transform 1 0 73136 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_649
timestamp 1669390400
transform 1 0 74032 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_651
timestamp 1669390400
transform 1 0 74256 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_654
timestamp 1669390400
transform 1 0 74592 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_670
timestamp 1669390400
transform 1 0 76384 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_686
timestamp 1669390400
transform 1 0 78176 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_17
timestamp 1669390400
transform 1 0 3248 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_21
timestamp 1669390400
transform 1 0 3696 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_29
timestamp 1669390400
transform 1 0 4592 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_33
timestamp 1669390400
transform 1 0 5040 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1669390400
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1669390400
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1669390400
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1669390400
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1669390400
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1669390400
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1669390400
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_353
timestamp 1669390400
transform 1 0 40880 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_369
timestamp 1669390400
transform 1 0 42672 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_383
timestamp 1669390400
transform 1 0 44240 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_387
timestamp 1669390400
transform 1 0 44688 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1669390400
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_399
timestamp 1669390400
transform 1 0 46032 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_403
timestamp 1669390400
transform 1 0 46480 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_407
timestamp 1669390400
transform 1 0 46928 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_439
timestamp 1669390400
transform 1 0 50512 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_455
timestamp 1669390400
transform 1 0 52304 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_459
timestamp 1669390400
transform 1 0 52752 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_463
timestamp 1669390400
transform 1 0 53200 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_527
timestamp 1669390400
transform 1 0 60368 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_531
timestamp 1669390400
transform 1 0 60816 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_534
timestamp 1669390400
transform 1 0 61152 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_598
timestamp 1669390400
transform 1 0 68320 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_602
timestamp 1669390400
transform 1 0 68768 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_605
timestamp 1669390400
transform 1 0 69104 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_637
timestamp 1669390400
transform 1 0 72688 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_645
timestamp 1669390400
transform 1 0 73584 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_649
timestamp 1669390400
transform 1 0 74032 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_651
timestamp 1669390400
transform 1 0 74256 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_654
timestamp 1669390400
transform 1 0 74592 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_670
timestamp 1669390400
transform 1 0 76384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_676
timestamp 1669390400
transform 1 0 77056 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_684
timestamp 1669390400
transform 1 0 77952 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_17
timestamp 1669390400
transform 1 0 3248 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_21
timestamp 1669390400
transform 1 0 3696 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_53
timestamp 1669390400
transform 1 0 7280 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_69
timestamp 1669390400
transform 1 0 9072 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1669390400
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1669390400
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1669390400
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1669390400
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1669390400
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1669390400
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1669390400
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_373
timestamp 1669390400
transform 1 0 43120 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_377
timestamp 1669390400
transform 1 0 43568 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_381
timestamp 1669390400
transform 1 0 44016 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_389
timestamp 1669390400
transform 1 0 44912 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_397
timestamp 1669390400
transform 1 0 45808 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_405
timestamp 1669390400
transform 1 0 46704 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_413
timestamp 1669390400
transform 1 0 47600 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_417
timestamp 1669390400
transform 1 0 48048 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_421
timestamp 1669390400
transform 1 0 48496 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1669390400
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_428
timestamp 1669390400
transform 1 0 49280 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_492
timestamp 1669390400
transform 1 0 56448 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_496
timestamp 1669390400
transform 1 0 56896 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_499
timestamp 1669390400
transform 1 0 57232 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_563
timestamp 1669390400
transform 1 0 64400 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_567
timestamp 1669390400
transform 1 0 64848 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_570
timestamp 1669390400
transform 1 0 65184 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_634
timestamp 1669390400
transform 1 0 72352 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_638
timestamp 1669390400
transform 1 0 72800 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_641
timestamp 1669390400
transform 1 0 73136 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_649
timestamp 1669390400
transform 1 0 74032 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_651
timestamp 1669390400
transform 1 0 74256 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_654
timestamp 1669390400
transform 1 0 74592 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_670
timestamp 1669390400
transform 1 0 76384 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_686
timestamp 1669390400
transform 1 0 78176 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_17
timestamp 1669390400
transform 1 0 3248 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_21
timestamp 1669390400
transform 1 0 3696 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_29
timestamp 1669390400
transform 1 0 4592 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_33
timestamp 1669390400
transform 1 0 5040 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1669390400
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1669390400
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_108
timestamp 1669390400
transform 1 0 13440 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_172
timestamp 1669390400
transform 1 0 20608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1669390400
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_179
timestamp 1669390400
transform 1 0 21392 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_243
timestamp 1669390400
transform 1 0 28560 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1669390400
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_250
timestamp 1669390400
transform 1 0 29344 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_314
timestamp 1669390400
transform 1 0 36512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1669390400
transform 1 0 36960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_321
timestamp 1669390400
transform 1 0 37296 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_385
timestamp 1669390400
transform 1 0 44464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_389
timestamp 1669390400
transform 1 0 44912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_392
timestamp 1669390400
transform 1 0 45248 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_394
timestamp 1669390400
transform 1 0 45472 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_401
timestamp 1669390400
transform 1 0 46256 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_411
timestamp 1669390400
transform 1 0 47376 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_415
timestamp 1669390400
transform 1 0 47824 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_419
timestamp 1669390400
transform 1 0 48272 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_451
timestamp 1669390400
transform 1 0 51856 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_459
timestamp 1669390400
transform 1 0 52752 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_463
timestamp 1669390400
transform 1 0 53200 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_527
timestamp 1669390400
transform 1 0 60368 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_531
timestamp 1669390400
transform 1 0 60816 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_534
timestamp 1669390400
transform 1 0 61152 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_598
timestamp 1669390400
transform 1 0 68320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_602
timestamp 1669390400
transform 1 0 68768 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_605
timestamp 1669390400
transform 1 0 69104 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_637
timestamp 1669390400
transform 1 0 72688 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_645
timestamp 1669390400
transform 1 0 73584 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_649
timestamp 1669390400
transform 1 0 74032 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_651
timestamp 1669390400
transform 1 0 74256 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_654
timestamp 1669390400
transform 1 0 74592 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_670
timestamp 1669390400
transform 1 0 76384 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_676
timestamp 1669390400
transform 1 0 77056 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_684
timestamp 1669390400
transform 1 0 77952 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_17
timestamp 1669390400
transform 1 0 3248 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_21
timestamp 1669390400
transform 1 0 3696 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_53
timestamp 1669390400
transform 1 0 7280 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_69
timestamp 1669390400
transform 1 0 9072 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_73
timestamp 1669390400
transform 1 0 9520 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_137
timestamp 1669390400
transform 1 0 16688 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1669390400
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_144
timestamp 1669390400
transform 1 0 17472 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_208
timestamp 1669390400
transform 1 0 24640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1669390400
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_215
timestamp 1669390400
transform 1 0 25424 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_279
timestamp 1669390400
transform 1 0 32592 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1669390400
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_286
timestamp 1669390400
transform 1 0 33376 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_350
timestamp 1669390400
transform 1 0 40544 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1669390400
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_357
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_389
timestamp 1669390400
transform 1 0 44912 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_399
timestamp 1669390400
transform 1 0 46032 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_407
timestamp 1669390400
transform 1 0 46928 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_409
timestamp 1669390400
transform 1 0 47152 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_416
timestamp 1669390400
transform 1 0 47936 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_420
timestamp 1669390400
transform 1 0 48384 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_424
timestamp 1669390400
transform 1 0 48832 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_428
timestamp 1669390400
transform 1 0 49280 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_492
timestamp 1669390400
transform 1 0 56448 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1669390400
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_499
timestamp 1669390400
transform 1 0 57232 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_563
timestamp 1669390400
transform 1 0 64400 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_567
timestamp 1669390400
transform 1 0 64848 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_570
timestamp 1669390400
transform 1 0 65184 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_634
timestamp 1669390400
transform 1 0 72352 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_638
timestamp 1669390400
transform 1 0 72800 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_641
timestamp 1669390400
transform 1 0 73136 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_649
timestamp 1669390400
transform 1 0 74032 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_651
timestamp 1669390400
transform 1 0 74256 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_654
timestamp 1669390400
transform 1 0 74592 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_670
timestamp 1669390400
transform 1 0 76384 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_686
timestamp 1669390400
transform 1 0 78176 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_17
timestamp 1669390400
transform 1 0 3248 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_21
timestamp 1669390400
transform 1 0 3696 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_29
timestamp 1669390400
transform 1 0 4592 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_33
timestamp 1669390400
transform 1 0 5040 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1669390400
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1669390400
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1669390400
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_108
timestamp 1669390400
transform 1 0 13440 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_172
timestamp 1669390400
transform 1 0 20608 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1669390400
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_179
timestamp 1669390400
transform 1 0 21392 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_243
timestamp 1669390400
transform 1 0 28560 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1669390400
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_250
timestamp 1669390400
transform 1 0 29344 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_314
timestamp 1669390400
transform 1 0 36512 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1669390400
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_321
timestamp 1669390400
transform 1 0 37296 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_385
timestamp 1669390400
transform 1 0 44464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1669390400
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_392
timestamp 1669390400
transform 1 0 45248 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_400
timestamp 1669390400
transform 1 0 46144 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_404
timestamp 1669390400
transform 1 0 46592 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_406
timestamp 1669390400
transform 1 0 46816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_413
timestamp 1669390400
transform 1 0 47600 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_415
timestamp 1669390400
transform 1 0 47824 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_422
timestamp 1669390400
transform 1 0 48608 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_426
timestamp 1669390400
transform 1 0 49056 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_428
timestamp 1669390400
transform 1 0 49280 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_433
timestamp 1669390400
transform 1 0 49840 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_437
timestamp 1669390400
transform 1 0 50288 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_453
timestamp 1669390400
transform 1 0 52080 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_463
timestamp 1669390400
transform 1 0 53200 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_527
timestamp 1669390400
transform 1 0 60368 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_531
timestamp 1669390400
transform 1 0 60816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_534
timestamp 1669390400
transform 1 0 61152 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_598
timestamp 1669390400
transform 1 0 68320 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_602
timestamp 1669390400
transform 1 0 68768 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_605
timestamp 1669390400
transform 1 0 69104 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_637
timestamp 1669390400
transform 1 0 72688 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_645
timestamp 1669390400
transform 1 0 73584 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_649
timestamp 1669390400
transform 1 0 74032 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_651
timestamp 1669390400
transform 1 0 74256 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_654
timestamp 1669390400
transform 1 0 74592 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_670
timestamp 1669390400
transform 1 0 76384 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_676
timestamp 1669390400
transform 1 0 77056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_679
timestamp 1669390400
transform 1 0 77392 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_687
timestamp 1669390400
transform 1 0 78288 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_17
timestamp 1669390400
transform 1 0 3248 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_33
timestamp 1669390400
transform 1 0 5040 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_37
timestamp 1669390400
transform 1 0 5488 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_69
timestamp 1669390400
transform 1 0 9072 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_73
timestamp 1669390400
transform 1 0 9520 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_137
timestamp 1669390400
transform 1 0 16688 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1669390400
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_144
timestamp 1669390400
transform 1 0 17472 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_208
timestamp 1669390400
transform 1 0 24640 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1669390400
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_215
timestamp 1669390400
transform 1 0 25424 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_279
timestamp 1669390400
transform 1 0 32592 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1669390400
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_286
timestamp 1669390400
transform 1 0 33376 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_350
timestamp 1669390400
transform 1 0 40544 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1669390400
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_357
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_389
timestamp 1669390400
transform 1 0 44912 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_405
timestamp 1669390400
transform 1 0 46704 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_415
timestamp 1669390400
transform 1 0 47824 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_423
timestamp 1669390400
transform 1 0 48720 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_425
timestamp 1669390400
transform 1 0 48944 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_428
timestamp 1669390400
transform 1 0 49280 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_439
timestamp 1669390400
transform 1 0 50512 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_471
timestamp 1669390400
transform 1 0 54096 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_487
timestamp 1669390400
transform 1 0 55888 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_495
timestamp 1669390400
transform 1 0 56784 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_499
timestamp 1669390400
transform 1 0 57232 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_563
timestamp 1669390400
transform 1 0 64400 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_567
timestamp 1669390400
transform 1 0 64848 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_570
timestamp 1669390400
transform 1 0 65184 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_604
timestamp 1669390400
transform 1 0 68992 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_636
timestamp 1669390400
transform 1 0 72576 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_638
timestamp 1669390400
transform 1 0 72800 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_641
timestamp 1669390400
transform 1 0 73136 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_649
timestamp 1669390400
transform 1 0 74032 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_651
timestamp 1669390400
transform 1 0 74256 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_654
timestamp 1669390400
transform 1 0 74592 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_670
timestamp 1669390400
transform 1 0 76384 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_686
timestamp 1669390400
transform 1 0 78176 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_19
timestamp 1669390400
transform 1 0 3472 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_23
timestamp 1669390400
transform 1 0 3920 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_27
timestamp 1669390400
transform 1 0 4368 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1669390400
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1669390400
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1669390400
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_108
timestamp 1669390400
transform 1 0 13440 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_172
timestamp 1669390400
transform 1 0 20608 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1669390400
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_179
timestamp 1669390400
transform 1 0 21392 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_243
timestamp 1669390400
transform 1 0 28560 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1669390400
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_250
timestamp 1669390400
transform 1 0 29344 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_314
timestamp 1669390400
transform 1 0 36512 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1669390400
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_321
timestamp 1669390400
transform 1 0 37296 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_385
timestamp 1669390400
transform 1 0 44464 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1669390400
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_392
timestamp 1669390400
transform 1 0 45248 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_408
timestamp 1669390400
transform 1 0 47040 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_416
timestamp 1669390400
transform 1 0 47936 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_419
timestamp 1669390400
transform 1 0 48272 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_423
timestamp 1669390400
transform 1 0 48720 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_425
timestamp 1669390400
transform 1 0 48944 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_436
timestamp 1669390400
transform 1 0 50176 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_442
timestamp 1669390400
transform 1 0 50848 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_446
timestamp 1669390400
transform 1 0 51296 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_454
timestamp 1669390400
transform 1 0 52192 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_458
timestamp 1669390400
transform 1 0 52640 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1669390400
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_463
timestamp 1669390400
transform 1 0 53200 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_527
timestamp 1669390400
transform 1 0 60368 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_531
timestamp 1669390400
transform 1 0 60816 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_534
timestamp 1669390400
transform 1 0 61152 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_566
timestamp 1669390400
transform 1 0 64736 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_584
timestamp 1669390400
transform 1 0 66752 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_590
timestamp 1669390400
transform 1 0 67424 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_602
timestamp 1669390400
transform 1 0 68768 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_605
timestamp 1669390400
transform 1 0 69104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_610
timestamp 1669390400
transform 1 0 69664 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_614
timestamp 1669390400
transform 1 0 70112 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_630
timestamp 1669390400
transform 1 0 71904 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_638
timestamp 1669390400
transform 1 0 72800 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_642
timestamp 1669390400
transform 1 0 73248 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_650
timestamp 1669390400
transform 1 0 74144 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_654
timestamp 1669390400
transform 1 0 74592 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_672
timestamp 1669390400
transform 1 0 76608 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_676
timestamp 1669390400
transform 1 0 77056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_679
timestamp 1669390400
transform 1 0 77392 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_687
timestamp 1669390400
transform 1 0 78288 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_19
timestamp 1669390400
transform 1 0 3472 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_23
timestamp 1669390400
transform 1 0 3920 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_55
timestamp 1669390400
transform 1 0 7504 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_73
timestamp 1669390400
transform 1 0 9520 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_137
timestamp 1669390400
transform 1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1669390400
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_144
timestamp 1669390400
transform 1 0 17472 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_208
timestamp 1669390400
transform 1 0 24640 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1669390400
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_215
timestamp 1669390400
transform 1 0 25424 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_279
timestamp 1669390400
transform 1 0 32592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1669390400
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_286
timestamp 1669390400
transform 1 0 33376 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_350
timestamp 1669390400
transform 1 0 40544 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1669390400
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_357
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_389
timestamp 1669390400
transform 1 0 44912 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_397
timestamp 1669390400
transform 1 0 45808 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_401
timestamp 1669390400
transform 1 0 46256 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_407
timestamp 1669390400
transform 1 0 46928 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_411
timestamp 1669390400
transform 1 0 47376 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_415
timestamp 1669390400
transform 1 0 47824 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_421
timestamp 1669390400
transform 1 0 48496 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1669390400
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_428
timestamp 1669390400
transform 1 0 49280 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_432
timestamp 1669390400
transform 1 0 49728 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_444
timestamp 1669390400
transform 1 0 51072 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_450
timestamp 1669390400
transform 1 0 51744 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_454
timestamp 1669390400
transform 1 0 52192 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_486
timestamp 1669390400
transform 1 0 55776 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_494
timestamp 1669390400
transform 1 0 56672 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_496
timestamp 1669390400
transform 1 0 56896 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_499
timestamp 1669390400
transform 1 0 57232 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_563
timestamp 1669390400
transform 1 0 64400 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_567
timestamp 1669390400
transform 1 0 64848 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_570
timestamp 1669390400
transform 1 0 65184 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_634
timestamp 1669390400
transform 1 0 72352 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_638
timestamp 1669390400
transform 1 0 72800 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_641
timestamp 1669390400
transform 1 0 73136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_652
timestamp 1669390400
transform 1 0 74368 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_672
timestamp 1669390400
transform 1 0 76608 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_676
timestamp 1669390400
transform 1 0 77056 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_684
timestamp 1669390400
transform 1 0 77952 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_19
timestamp 1669390400
transform 1 0 3472 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_23
timestamp 1669390400
transform 1 0 3920 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_31
timestamp 1669390400
transform 1 0 4816 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1669390400
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1669390400
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1669390400
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_108
timestamp 1669390400
transform 1 0 13440 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_172
timestamp 1669390400
transform 1 0 20608 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1669390400
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1669390400
transform 1 0 21392 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1669390400
transform 1 0 28560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1669390400
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_250
timestamp 1669390400
transform 1 0 29344 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_314
timestamp 1669390400
transform 1 0 36512 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1669390400
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_321
timestamp 1669390400
transform 1 0 37296 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_385
timestamp 1669390400
transform 1 0 44464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1669390400
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_392
timestamp 1669390400
transform 1 0 45248 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_426
timestamp 1669390400
transform 1 0 49056 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_432
timestamp 1669390400
transform 1 0 49728 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_446
timestamp 1669390400
transform 1 0 51296 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_452
timestamp 1669390400
transform 1 0 51968 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_456
timestamp 1669390400
transform 1 0 52416 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1669390400
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_463
timestamp 1669390400
transform 1 0 53200 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_470
timestamp 1669390400
transform 1 0 53984 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_502
timestamp 1669390400
transform 1 0 57568 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_518
timestamp 1669390400
transform 1 0 59360 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_526
timestamp 1669390400
transform 1 0 60256 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_530
timestamp 1669390400
transform 1 0 60704 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_534
timestamp 1669390400
transform 1 0 61152 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_598
timestamp 1669390400
transform 1 0 68320 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_602
timestamp 1669390400
transform 1 0 68768 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_605
timestamp 1669390400
transform 1 0 69104 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_621
timestamp 1669390400
transform 1 0 70896 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_629
timestamp 1669390400
transform 1 0 71792 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_633
timestamp 1669390400
transform 1 0 72240 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_639
timestamp 1669390400
transform 1 0 72912 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_641
timestamp 1669390400
transform 1 0 73136 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_646
timestamp 1669390400
transform 1 0 73696 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_650
timestamp 1669390400
transform 1 0 74144 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_654
timestamp 1669390400
transform 1 0 74592 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_672
timestamp 1669390400
transform 1 0 76608 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_676
timestamp 1669390400
transform 1 0 77056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_679
timestamp 1669390400
transform 1 0 77392 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_687
timestamp 1669390400
transform 1 0 78288 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_19
timestamp 1669390400
transform 1 0 3472 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_23
timestamp 1669390400
transform 1 0 3920 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_55
timestamp 1669390400
transform 1 0 7504 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_73
timestamp 1669390400
transform 1 0 9520 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_137
timestamp 1669390400
transform 1 0 16688 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1669390400
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_144
timestamp 1669390400
transform 1 0 17472 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_208
timestamp 1669390400
transform 1 0 24640 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1669390400
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1669390400
transform 1 0 25424 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1669390400
transform 1 0 32592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1669390400
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_286
timestamp 1669390400
transform 1 0 33376 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_350
timestamp 1669390400
transform 1 0 40544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1669390400
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_357
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_421
timestamp 1669390400
transform 1 0 48496 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1669390400
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_428
timestamp 1669390400
transform 1 0 49280 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_431
timestamp 1669390400
transform 1 0 49616 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_447
timestamp 1669390400
transform 1 0 51408 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_459
timestamp 1669390400
transform 1 0 52752 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_469
timestamp 1669390400
transform 1 0 53872 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_487
timestamp 1669390400
transform 1 0 55888 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_495
timestamp 1669390400
transform 1 0 56784 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_499
timestamp 1669390400
transform 1 0 57232 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_563
timestamp 1669390400
transform 1 0 64400 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_567
timestamp 1669390400
transform 1 0 64848 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_570
timestamp 1669390400
transform 1 0 65184 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_634
timestamp 1669390400
transform 1 0 72352 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_638
timestamp 1669390400
transform 1 0 72800 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_641
timestamp 1669390400
transform 1 0 73136 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_649
timestamp 1669390400
transform 1 0 74032 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_653
timestamp 1669390400
transform 1 0 74480 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_655
timestamp 1669390400
transform 1 0 74704 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_672
timestamp 1669390400
transform 1 0 76608 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_676
timestamp 1669390400
transform 1 0 77056 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_684
timestamp 1669390400
transform 1 0 77952 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_19
timestamp 1669390400
transform 1 0 3472 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_23
timestamp 1669390400
transform 1 0 3920 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_31
timestamp 1669390400
transform 1 0 4816 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1669390400
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1669390400
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1669390400
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1669390400
transform 1 0 13440 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_172
timestamp 1669390400
transform 1 0 20608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1669390400
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1669390400
transform 1 0 21392 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_243
timestamp 1669390400
transform 1 0 28560 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1669390400
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1669390400
transform 1 0 29344 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1669390400
transform 1 0 36512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1669390400
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_321
timestamp 1669390400
transform 1 0 37296 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_385
timestamp 1669390400
transform 1 0 44464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1669390400
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_392
timestamp 1669390400
transform 1 0 45248 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_408
timestamp 1669390400
transform 1 0 47040 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_416
timestamp 1669390400
transform 1 0 47936 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_422
timestamp 1669390400
transform 1 0 48608 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_426
timestamp 1669390400
transform 1 0 49056 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_428
timestamp 1669390400
transform 1 0 49280 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_433
timestamp 1669390400
transform 1 0 49840 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_437
timestamp 1669390400
transform 1 0 50288 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_444
timestamp 1669390400
transform 1 0 51072 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_448
timestamp 1669390400
transform 1 0 51520 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_460
timestamp 1669390400
transform 1 0 52864 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_463
timestamp 1669390400
transform 1 0 53200 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_474
timestamp 1669390400
transform 1 0 54432 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_482
timestamp 1669390400
transform 1 0 55328 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_485
timestamp 1669390400
transform 1 0 55664 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_493
timestamp 1669390400
transform 1 0 56560 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_501
timestamp 1669390400
transform 1 0 57456 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_509
timestamp 1669390400
transform 1 0 58352 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_513
timestamp 1669390400
transform 1 0 58800 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_515
timestamp 1669390400
transform 1 0 59024 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_520
timestamp 1669390400
transform 1 0 59584 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_524
timestamp 1669390400
transform 1 0 60032 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_526
timestamp 1669390400
transform 1 0 60256 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_531
timestamp 1669390400
transform 1 0 60816 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_534
timestamp 1669390400
transform 1 0 61152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_537
timestamp 1669390400
transform 1 0 61488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_601
timestamp 1669390400
transform 1 0 68656 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_605
timestamp 1669390400
transform 1 0 69104 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_637
timestamp 1669390400
transform 1 0 72688 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_653
timestamp 1669390400
transform 1 0 74480 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_655
timestamp 1669390400
transform 1 0 74704 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_672
timestamp 1669390400
transform 1 0 76608 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_676
timestamp 1669390400
transform 1 0 77056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_679
timestamp 1669390400
transform 1 0 77392 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_687
timestamp 1669390400
transform 1 0 78288 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_19
timestamp 1669390400
transform 1 0 3472 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_23
timestamp 1669390400
transform 1 0 3920 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_55
timestamp 1669390400
transform 1 0 7504 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1669390400
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_137
timestamp 1669390400
transform 1 0 16688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1669390400
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1669390400
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1669390400
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1669390400
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1669390400
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1669390400
transform 1 0 32592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1669390400
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_286
timestamp 1669390400
transform 1 0 33376 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_350
timestamp 1669390400
transform 1 0 40544 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1669390400
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_357
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_389
timestamp 1669390400
transform 1 0 44912 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_405
timestamp 1669390400
transform 1 0 46704 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_413
timestamp 1669390400
transform 1 0 47600 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_416
timestamp 1669390400
transform 1 0 47936 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_422
timestamp 1669390400
transform 1 0 48608 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_428
timestamp 1669390400
transform 1 0 49280 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_436
timestamp 1669390400
transform 1 0 50176 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_441
timestamp 1669390400
transform 1 0 50736 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_445
timestamp 1669390400
transform 1 0 51184 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_447
timestamp 1669390400
transform 1 0 51408 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_454
timestamp 1669390400
transform 1 0 52192 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_468
timestamp 1669390400
transform 1 0 53760 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_472
timestamp 1669390400
transform 1 0 54208 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_488
timestamp 1669390400
transform 1 0 56000 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_492
timestamp 1669390400
transform 1 0 56448 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_495
timestamp 1669390400
transform 1 0 56784 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_499
timestamp 1669390400
transform 1 0 57232 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_504
timestamp 1669390400
transform 1 0 57792 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_508
timestamp 1669390400
transform 1 0 58240 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_540
timestamp 1669390400
transform 1 0 61824 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_556
timestamp 1669390400
transform 1 0 63616 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_564
timestamp 1669390400
transform 1 0 64512 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_570
timestamp 1669390400
transform 1 0 65184 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_634
timestamp 1669390400
transform 1 0 72352 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_638
timestamp 1669390400
transform 1 0 72800 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_641
timestamp 1669390400
transform 1 0 73136 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_649
timestamp 1669390400
transform 1 0 74032 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_653
timestamp 1669390400
transform 1 0 74480 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_655
timestamp 1669390400
transform 1 0 74704 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_672
timestamp 1669390400
transform 1 0 76608 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_676
timestamp 1669390400
transform 1 0 77056 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_684
timestamp 1669390400
transform 1 0 77952 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_19
timestamp 1669390400
transform 1 0 3472 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_23
timestamp 1669390400
transform 1 0 3920 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_31
timestamp 1669390400
transform 1 0 4816 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1669390400
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1669390400
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1669390400
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1669390400
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1669390400
transform 1 0 20608 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1669390400
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1669390400
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1669390400
transform 1 0 28560 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1669390400
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1669390400
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1669390400
transform 1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1669390400
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_321
timestamp 1669390400
transform 1 0 37296 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_385
timestamp 1669390400
transform 1 0 44464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1669390400
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_392
timestamp 1669390400
transform 1 0 45248 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_424
timestamp 1669390400
transform 1 0 48832 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_440
timestamp 1669390400
transform 1 0 50624 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_448
timestamp 1669390400
transform 1 0 51520 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_452
timestamp 1669390400
transform 1 0 51968 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_456
timestamp 1669390400
transform 1 0 52416 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_460
timestamp 1669390400
transform 1 0 52864 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_463
timestamp 1669390400
transform 1 0 53200 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_468
timestamp 1669390400
transform 1 0 53760 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_470
timestamp 1669390400
transform 1 0 53984 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_481
timestamp 1669390400
transform 1 0 55216 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_489
timestamp 1669390400
transform 1 0 56112 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_493
timestamp 1669390400
transform 1 0 56560 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_495
timestamp 1669390400
transform 1 0 56784 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_502
timestamp 1669390400
transform 1 0 57568 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_518
timestamp 1669390400
transform 1 0 59360 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_526
timestamp 1669390400
transform 1 0 60256 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_530
timestamp 1669390400
transform 1 0 60704 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_534
timestamp 1669390400
transform 1 0 61152 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_598
timestamp 1669390400
transform 1 0 68320 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_602
timestamp 1669390400
transform 1 0 68768 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_605
timestamp 1669390400
transform 1 0 69104 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_637
timestamp 1669390400
transform 1 0 72688 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_653
timestamp 1669390400
transform 1 0 74480 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_655
timestamp 1669390400
transform 1 0 74704 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_672
timestamp 1669390400
transform 1 0 76608 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_676
timestamp 1669390400
transform 1 0 77056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_679
timestamp 1669390400
transform 1 0 77392 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_687
timestamp 1669390400
transform 1 0 78288 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_19
timestamp 1669390400
transform 1 0 3472 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_23
timestamp 1669390400
transform 1 0 3920 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_55
timestamp 1669390400
transform 1 0 7504 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1669390400
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1669390400
transform 1 0 16688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1669390400
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1669390400
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1669390400
transform 1 0 24640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1669390400
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1669390400
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1669390400
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1669390400
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1669390400
transform 1 0 33376 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_350
timestamp 1669390400
transform 1 0 40544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1669390400
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_357
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_421
timestamp 1669390400
transform 1 0 48496 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1669390400
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_428
timestamp 1669390400
transform 1 0 49280 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_444
timestamp 1669390400
transform 1 0 51072 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_450
timestamp 1669390400
transform 1 0 51744 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_456
timestamp 1669390400
transform 1 0 52416 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_462
timestamp 1669390400
transform 1 0 53088 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_466
timestamp 1669390400
transform 1 0 53536 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_472
timestamp 1669390400
transform 1 0 54208 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_484
timestamp 1669390400
transform 1 0 55552 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_490
timestamp 1669390400
transform 1 0 56224 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_496
timestamp 1669390400
transform 1 0 56896 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_499
timestamp 1669390400
transform 1 0 57232 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_502
timestamp 1669390400
transform 1 0 57568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_566
timestamp 1669390400
transform 1 0 64736 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_570
timestamp 1669390400
transform 1 0 65184 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_634
timestamp 1669390400
transform 1 0 72352 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_638
timestamp 1669390400
transform 1 0 72800 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_641
timestamp 1669390400
transform 1 0 73136 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_649
timestamp 1669390400
transform 1 0 74032 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_653
timestamp 1669390400
transform 1 0 74480 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_655
timestamp 1669390400
transform 1 0 74704 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_672
timestamp 1669390400
transform 1 0 76608 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_676
timestamp 1669390400
transform 1 0 77056 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_684
timestamp 1669390400
transform 1 0 77952 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_19
timestamp 1669390400
transform 1 0 3472 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_23
timestamp 1669390400
transform 1 0 3920 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_31
timestamp 1669390400
transform 1 0 4816 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1669390400
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1669390400
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1669390400
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_108
timestamp 1669390400
transform 1 0 13440 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_172
timestamp 1669390400
transform 1 0 20608 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1669390400
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1669390400
transform 1 0 21392 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_243
timestamp 1669390400
transform 1 0 28560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1669390400
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1669390400
transform 1 0 29344 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1669390400
transform 1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1669390400
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_321
timestamp 1669390400
transform 1 0 37296 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_385
timestamp 1669390400
transform 1 0 44464 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1669390400
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_392
timestamp 1669390400
transform 1 0 45248 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_424
timestamp 1669390400
transform 1 0 48832 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_432
timestamp 1669390400
transform 1 0 49728 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_436
timestamp 1669390400
transform 1 0 50176 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_438
timestamp 1669390400
transform 1 0 50400 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_443
timestamp 1669390400
transform 1 0 50960 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_447
timestamp 1669390400
transform 1 0 51408 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_455
timestamp 1669390400
transform 1 0 52304 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_459
timestamp 1669390400
transform 1 0 52752 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_463
timestamp 1669390400
transform 1 0 53200 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_465
timestamp 1669390400
transform 1 0 53424 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_468
timestamp 1669390400
transform 1 0 53760 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_476
timestamp 1669390400
transform 1 0 54656 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_478
timestamp 1669390400
transform 1 0 54880 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_489
timestamp 1669390400
transform 1 0 56112 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_493
timestamp 1669390400
transform 1 0 56560 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_501
timestamp 1669390400
transform 1 0 57456 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_505
timestamp 1669390400
transform 1 0 57904 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_521
timestamp 1669390400
transform 1 0 59696 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_529
timestamp 1669390400
transform 1 0 60592 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_531
timestamp 1669390400
transform 1 0 60816 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_534
timestamp 1669390400
transform 1 0 61152 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_598
timestamp 1669390400
transform 1 0 68320 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_602
timestamp 1669390400
transform 1 0 68768 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_605
timestamp 1669390400
transform 1 0 69104 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_637
timestamp 1669390400
transform 1 0 72688 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_653
timestamp 1669390400
transform 1 0 74480 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_655
timestamp 1669390400
transform 1 0 74704 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_672
timestamp 1669390400
transform 1 0 76608 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_676
timestamp 1669390400
transform 1 0 77056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_679
timestamp 1669390400
transform 1 0 77392 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_687
timestamp 1669390400
transform 1 0 78288 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_19
timestamp 1669390400
transform 1 0 3472 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_23
timestamp 1669390400
transform 1 0 3920 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_55
timestamp 1669390400
transform 1 0 7504 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_73
timestamp 1669390400
transform 1 0 9520 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_137
timestamp 1669390400
transform 1 0 16688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_141
timestamp 1669390400
transform 1 0 17136 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_144
timestamp 1669390400
transform 1 0 17472 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_208
timestamp 1669390400
transform 1 0 24640 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1669390400
transform 1 0 25088 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_215
timestamp 1669390400
transform 1 0 25424 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_279
timestamp 1669390400
transform 1 0 32592 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_283
timestamp 1669390400
transform 1 0 33040 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_286
timestamp 1669390400
transform 1 0 33376 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_350
timestamp 1669390400
transform 1 0 40544 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1669390400
transform 1 0 40992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_357
timestamp 1669390400
transform 1 0 41328 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_421
timestamp 1669390400
transform 1 0 48496 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_425
timestamp 1669390400
transform 1 0 48944 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_428
timestamp 1669390400
transform 1 0 49280 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_460
timestamp 1669390400
transform 1 0 52864 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_465
timestamp 1669390400
transform 1 0 53424 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_469
timestamp 1669390400
transform 1 0 53872 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_473
timestamp 1669390400
transform 1 0 54320 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_475
timestamp 1669390400
transform 1 0 54544 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_478
timestamp 1669390400
transform 1 0 54880 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_490
timestamp 1669390400
transform 1 0 56224 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_496
timestamp 1669390400
transform 1 0 56896 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_499
timestamp 1669390400
transform 1 0 57232 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_510
timestamp 1669390400
transform 1 0 58464 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_542
timestamp 1669390400
transform 1 0 62048 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_558
timestamp 1669390400
transform 1 0 63840 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_566
timestamp 1669390400
transform 1 0 64736 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_570
timestamp 1669390400
transform 1 0 65184 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_634
timestamp 1669390400
transform 1 0 72352 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_638
timestamp 1669390400
transform 1 0 72800 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_641
timestamp 1669390400
transform 1 0 73136 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_649
timestamp 1669390400
transform 1 0 74032 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_653
timestamp 1669390400
transform 1 0 74480 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_655
timestamp 1669390400
transform 1 0 74704 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_672
timestamp 1669390400
transform 1 0 76608 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_676
timestamp 1669390400
transform 1 0 77056 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_684
timestamp 1669390400
transform 1 0 77952 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_2
timestamp 1669390400
transform 1 0 1568 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_19
timestamp 1669390400
transform 1 0 3472 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_23
timestamp 1669390400
transform 1 0 3920 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_31
timestamp 1669390400
transform 1 0 4816 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_37
timestamp 1669390400
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_101
timestamp 1669390400
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_105
timestamp 1669390400
transform 1 0 13104 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_108
timestamp 1669390400
transform 1 0 13440 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_172
timestamp 1669390400
transform 1 0 20608 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_176
timestamp 1669390400
transform 1 0 21056 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_179
timestamp 1669390400
transform 1 0 21392 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_243
timestamp 1669390400
transform 1 0 28560 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_247
timestamp 1669390400
transform 1 0 29008 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_250
timestamp 1669390400
transform 1 0 29344 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_314
timestamp 1669390400
transform 1 0 36512 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_318
timestamp 1669390400
transform 1 0 36960 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_321
timestamp 1669390400
transform 1 0 37296 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_385
timestamp 1669390400
transform 1 0 44464 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_389
timestamp 1669390400
transform 1 0 44912 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_392
timestamp 1669390400
transform 1 0 45248 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_456
timestamp 1669390400
transform 1 0 52416 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_460
timestamp 1669390400
transform 1 0 52864 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_463
timestamp 1669390400
transform 1 0 53200 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_479
timestamp 1669390400
transform 1 0 54992 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_487
timestamp 1669390400
transform 1 0 55888 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_490
timestamp 1669390400
transform 1 0 56224 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_496
timestamp 1669390400
transform 1 0 56896 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_508
timestamp 1669390400
transform 1 0 58240 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_516
timestamp 1669390400
transform 1 0 59136 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_520
timestamp 1669390400
transform 1 0 59584 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_528
timestamp 1669390400
transform 1 0 60480 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_534
timestamp 1669390400
transform 1 0 61152 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_598
timestamp 1669390400
transform 1 0 68320 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_602
timestamp 1669390400
transform 1 0 68768 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_605
timestamp 1669390400
transform 1 0 69104 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_637
timestamp 1669390400
transform 1 0 72688 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_653
timestamp 1669390400
transform 1 0 74480 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_655
timestamp 1669390400
transform 1 0 74704 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_672
timestamp 1669390400
transform 1 0 76608 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_676
timestamp 1669390400
transform 1 0 77056 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_679
timestamp 1669390400
transform 1 0 77392 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_687
timestamp 1669390400
transform 1 0 78288 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_2
timestamp 1669390400
transform 1 0 1568 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_19
timestamp 1669390400
transform 1 0 3472 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_23
timestamp 1669390400
transform 1 0 3920 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_55
timestamp 1669390400
transform 1 0 7504 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_73
timestamp 1669390400
transform 1 0 9520 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_137
timestamp 1669390400
transform 1 0 16688 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_141
timestamp 1669390400
transform 1 0 17136 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_144
timestamp 1669390400
transform 1 0 17472 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_208
timestamp 1669390400
transform 1 0 24640 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1669390400
transform 1 0 25088 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_215
timestamp 1669390400
transform 1 0 25424 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_279
timestamp 1669390400
transform 1 0 32592 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_283
timestamp 1669390400
transform 1 0 33040 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_286
timestamp 1669390400
transform 1 0 33376 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_350
timestamp 1669390400
transform 1 0 40544 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_354
timestamp 1669390400
transform 1 0 40992 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_357
timestamp 1669390400
transform 1 0 41328 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_421
timestamp 1669390400
transform 1 0 48496 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_425
timestamp 1669390400
transform 1 0 48944 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_428
timestamp 1669390400
transform 1 0 49280 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_460
timestamp 1669390400
transform 1 0 52864 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_468
timestamp 1669390400
transform 1 0 53760 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_472
timestamp 1669390400
transform 1 0 54208 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_474
timestamp 1669390400
transform 1 0 54432 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_477
timestamp 1669390400
transform 1 0 54768 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_483
timestamp 1669390400
transform 1 0 55440 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_491
timestamp 1669390400
transform 1 0 56336 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_495
timestamp 1669390400
transform 1 0 56784 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_499
timestamp 1669390400
transform 1 0 57232 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_501
timestamp 1669390400
transform 1 0 57456 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_512
timestamp 1669390400
transform 1 0 58688 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_544
timestamp 1669390400
transform 1 0 62272 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_546
timestamp 1669390400
transform 1 0 62496 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_551
timestamp 1669390400
transform 1 0 63056 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_555
timestamp 1669390400
transform 1 0 63504 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_563
timestamp 1669390400
transform 1 0 64400 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_567
timestamp 1669390400
transform 1 0 64848 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_570
timestamp 1669390400
transform 1 0 65184 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_634
timestamp 1669390400
transform 1 0 72352 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_638
timestamp 1669390400
transform 1 0 72800 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_641
timestamp 1669390400
transform 1 0 73136 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_649
timestamp 1669390400
transform 1 0 74032 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_653
timestamp 1669390400
transform 1 0 74480 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_655
timestamp 1669390400
transform 1 0 74704 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_672
timestamp 1669390400
transform 1 0 76608 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_676
timestamp 1669390400
transform 1 0 77056 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_684
timestamp 1669390400
transform 1 0 77952 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_2
timestamp 1669390400
transform 1 0 1568 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_19
timestamp 1669390400
transform 1 0 3472 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_23
timestamp 1669390400
transform 1 0 3920 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_27
timestamp 1669390400
transform 1 0 4368 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_37
timestamp 1669390400
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_101
timestamp 1669390400
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_105
timestamp 1669390400
transform 1 0 13104 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_108
timestamp 1669390400
transform 1 0 13440 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_172
timestamp 1669390400
transform 1 0 20608 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_176
timestamp 1669390400
transform 1 0 21056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_179
timestamp 1669390400
transform 1 0 21392 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_243
timestamp 1669390400
transform 1 0 28560 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_247
timestamp 1669390400
transform 1 0 29008 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_250
timestamp 1669390400
transform 1 0 29344 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_314
timestamp 1669390400
transform 1 0 36512 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_318
timestamp 1669390400
transform 1 0 36960 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_321
timestamp 1669390400
transform 1 0 37296 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_385
timestamp 1669390400
transform 1 0 44464 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_389
timestamp 1669390400
transform 1 0 44912 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_392
timestamp 1669390400
transform 1 0 45248 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_456
timestamp 1669390400
transform 1 0 52416 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_460
timestamp 1669390400
transform 1 0 52864 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_463
timestamp 1669390400
transform 1 0 53200 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_479
timestamp 1669390400
transform 1 0 54992 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_487
timestamp 1669390400
transform 1 0 55888 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_491
timestamp 1669390400
transform 1 0 56336 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_495
timestamp 1669390400
transform 1 0 56784 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_501
timestamp 1669390400
transform 1 0 57456 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_513
timestamp 1669390400
transform 1 0 58800 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_519
timestamp 1669390400
transform 1 0 59472 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_523
timestamp 1669390400
transform 1 0 59920 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_531
timestamp 1669390400
transform 1 0 60816 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_534
timestamp 1669390400
transform 1 0 61152 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_598
timestamp 1669390400
transform 1 0 68320 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_602
timestamp 1669390400
transform 1 0 68768 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_605
timestamp 1669390400
transform 1 0 69104 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_637
timestamp 1669390400
transform 1 0 72688 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_653
timestamp 1669390400
transform 1 0 74480 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_655
timestamp 1669390400
transform 1 0 74704 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_672
timestamp 1669390400
transform 1 0 76608 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_676
timestamp 1669390400
transform 1 0 77056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_679
timestamp 1669390400
transform 1 0 77392 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_687
timestamp 1669390400
transform 1 0 78288 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_2
timestamp 1669390400
transform 1 0 1568 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_19
timestamp 1669390400
transform 1 0 3472 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_37
timestamp 1669390400
transform 1 0 5488 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_69
timestamp 1669390400
transform 1 0 9072 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_73
timestamp 1669390400
transform 1 0 9520 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_137
timestamp 1669390400
transform 1 0 16688 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_141
timestamp 1669390400
transform 1 0 17136 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_144
timestamp 1669390400
transform 1 0 17472 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_208
timestamp 1669390400
transform 1 0 24640 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_212
timestamp 1669390400
transform 1 0 25088 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_215
timestamp 1669390400
transform 1 0 25424 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_279
timestamp 1669390400
transform 1 0 32592 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_283
timestamp 1669390400
transform 1 0 33040 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_286
timestamp 1669390400
transform 1 0 33376 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_350
timestamp 1669390400
transform 1 0 40544 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_354
timestamp 1669390400
transform 1 0 40992 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_357
timestamp 1669390400
transform 1 0 41328 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_421
timestamp 1669390400
transform 1 0 48496 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_425
timestamp 1669390400
transform 1 0 48944 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_428
timestamp 1669390400
transform 1 0 49280 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_492
timestamp 1669390400
transform 1 0 56448 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_496
timestamp 1669390400
transform 1 0 56896 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_499
timestamp 1669390400
transform 1 0 57232 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_505
timestamp 1669390400
transform 1 0 57904 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_507
timestamp 1669390400
transform 1 0 58128 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_512
timestamp 1669390400
transform 1 0 58688 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_516
timestamp 1669390400
transform 1 0 59136 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_528
timestamp 1669390400
transform 1 0 60480 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_538
timestamp 1669390400
transform 1 0 61600 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_542
timestamp 1669390400
transform 1 0 62048 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_558
timestamp 1669390400
transform 1 0 63840 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_566
timestamp 1669390400
transform 1 0 64736 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_570
timestamp 1669390400
transform 1 0 65184 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_634
timestamp 1669390400
transform 1 0 72352 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_638
timestamp 1669390400
transform 1 0 72800 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_641
timestamp 1669390400
transform 1 0 73136 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_649
timestamp 1669390400
transform 1 0 74032 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_651
timestamp 1669390400
transform 1 0 74256 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_654
timestamp 1669390400
transform 1 0 74592 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_672
timestamp 1669390400
transform 1 0 76608 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_676
timestamp 1669390400
transform 1 0 77056 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_684
timestamp 1669390400
transform 1 0 77952 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_2
timestamp 1669390400
transform 1 0 1568 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_19
timestamp 1669390400
transform 1 0 3472 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_23
timestamp 1669390400
transform 1 0 3920 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_27
timestamp 1669390400
transform 1 0 4368 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_37
timestamp 1669390400
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_101
timestamp 1669390400
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_105
timestamp 1669390400
transform 1 0 13104 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_108
timestamp 1669390400
transform 1 0 13440 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_172
timestamp 1669390400
transform 1 0 20608 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_176
timestamp 1669390400
transform 1 0 21056 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_179
timestamp 1669390400
transform 1 0 21392 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_243
timestamp 1669390400
transform 1 0 28560 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_247
timestamp 1669390400
transform 1 0 29008 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_250
timestamp 1669390400
transform 1 0 29344 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_314
timestamp 1669390400
transform 1 0 36512 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_318
timestamp 1669390400
transform 1 0 36960 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_321
timestamp 1669390400
transform 1 0 37296 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_385
timestamp 1669390400
transform 1 0 44464 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_389
timestamp 1669390400
transform 1 0 44912 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_392
timestamp 1669390400
transform 1 0 45248 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_456
timestamp 1669390400
transform 1 0 52416 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_460
timestamp 1669390400
transform 1 0 52864 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_463
timestamp 1669390400
transform 1 0 53200 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_479
timestamp 1669390400
transform 1 0 54992 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_487
timestamp 1669390400
transform 1 0 55888 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_489
timestamp 1669390400
transform 1 0 56112 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_492
timestamp 1669390400
transform 1 0 56448 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_500
timestamp 1669390400
transform 1 0 57344 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_504
timestamp 1669390400
transform 1 0 57792 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_509
timestamp 1669390400
transform 1 0 58352 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_511
timestamp 1669390400
transform 1 0 58576 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_516
timestamp 1669390400
transform 1 0 59136 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_520
timestamp 1669390400
transform 1 0 59584 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_531
timestamp 1669390400
transform 1 0 60816 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_534
timestamp 1669390400
transform 1 0 61152 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_539
timestamp 1669390400
transform 1 0 61712 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_543
timestamp 1669390400
transform 1 0 62160 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_575
timestamp 1669390400
transform 1 0 65744 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_579
timestamp 1669390400
transform 1 0 66192 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_584
timestamp 1669390400
transform 1 0 66752 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_588
timestamp 1669390400
transform 1 0 67200 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_596
timestamp 1669390400
transform 1 0 68096 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_600
timestamp 1669390400
transform 1 0 68544 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_602
timestamp 1669390400
transform 1 0 68768 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_605
timestamp 1669390400
transform 1 0 69104 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_637
timestamp 1669390400
transform 1 0 72688 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_654
timestamp 1669390400
transform 1 0 74592 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_672
timestamp 1669390400
transform 1 0 76608 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_676
timestamp 1669390400
transform 1 0 77056 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_679
timestamp 1669390400
transform 1 0 77392 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_687
timestamp 1669390400
transform 1 0 78288 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_2
timestamp 1669390400
transform 1 0 1568 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_19
timestamp 1669390400
transform 1 0 3472 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_23
timestamp 1669390400
transform 1 0 3920 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_55
timestamp 1669390400
transform 1 0 7504 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_73
timestamp 1669390400
transform 1 0 9520 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_137
timestamp 1669390400
transform 1 0 16688 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_141
timestamp 1669390400
transform 1 0 17136 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_144
timestamp 1669390400
transform 1 0 17472 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_208
timestamp 1669390400
transform 1 0 24640 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_212
timestamp 1669390400
transform 1 0 25088 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_215
timestamp 1669390400
transform 1 0 25424 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_279
timestamp 1669390400
transform 1 0 32592 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_283
timestamp 1669390400
transform 1 0 33040 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_286
timestamp 1669390400
transform 1 0 33376 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_350
timestamp 1669390400
transform 1 0 40544 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_354
timestamp 1669390400
transform 1 0 40992 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_357
timestamp 1669390400
transform 1 0 41328 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_421
timestamp 1669390400
transform 1 0 48496 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_425
timestamp 1669390400
transform 1 0 48944 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_428
timestamp 1669390400
transform 1 0 49280 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_492
timestamp 1669390400
transform 1 0 56448 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_496
timestamp 1669390400
transform 1 0 56896 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_499
timestamp 1669390400
transform 1 0 57232 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_504
timestamp 1669390400
transform 1 0 57792 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_508
timestamp 1669390400
transform 1 0 58240 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_512
timestamp 1669390400
transform 1 0 58688 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_516
timestamp 1669390400
transform 1 0 59136 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_523
timestamp 1669390400
transform 1 0 59920 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_527
timestamp 1669390400
transform 1 0 60368 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_538
timestamp 1669390400
transform 1 0 61600 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_550
timestamp 1669390400
transform 1 0 62944 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_558
timestamp 1669390400
transform 1 0 63840 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_566
timestamp 1669390400
transform 1 0 64736 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_570
timestamp 1669390400
transform 1 0 65184 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_573
timestamp 1669390400
transform 1 0 65520 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_637
timestamp 1669390400
transform 1 0 72688 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_641
timestamp 1669390400
transform 1 0 73136 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_649
timestamp 1669390400
transform 1 0 74032 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_653
timestamp 1669390400
transform 1 0 74480 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_655
timestamp 1669390400
transform 1 0 74704 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_672
timestamp 1669390400
transform 1 0 76608 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_676
timestamp 1669390400
transform 1 0 77056 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_684
timestamp 1669390400
transform 1 0 77952 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_2
timestamp 1669390400
transform 1 0 1568 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_19
timestamp 1669390400
transform 1 0 3472 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_23
timestamp 1669390400
transform 1 0 3920 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_31
timestamp 1669390400
transform 1 0 4816 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_37
timestamp 1669390400
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_101
timestamp 1669390400
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_105
timestamp 1669390400
transform 1 0 13104 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_108
timestamp 1669390400
transform 1 0 13440 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_172
timestamp 1669390400
transform 1 0 20608 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_176
timestamp 1669390400
transform 1 0 21056 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_179
timestamp 1669390400
transform 1 0 21392 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_243
timestamp 1669390400
transform 1 0 28560 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_247
timestamp 1669390400
transform 1 0 29008 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_250
timestamp 1669390400
transform 1 0 29344 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_314
timestamp 1669390400
transform 1 0 36512 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_318
timestamp 1669390400
transform 1 0 36960 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_321
timestamp 1669390400
transform 1 0 37296 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_385
timestamp 1669390400
transform 1 0 44464 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_389
timestamp 1669390400
transform 1 0 44912 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_392
timestamp 1669390400
transform 1 0 45248 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_456
timestamp 1669390400
transform 1 0 52416 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_460
timestamp 1669390400
transform 1 0 52864 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_463
timestamp 1669390400
transform 1 0 53200 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_495
timestamp 1669390400
transform 1 0 56784 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_511
timestamp 1669390400
transform 1 0 58576 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_517
timestamp 1669390400
transform 1 0 59248 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_523
timestamp 1669390400
transform 1 0 59920 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_529
timestamp 1669390400
transform 1 0 60592 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_531
timestamp 1669390400
transform 1 0 60816 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_534
timestamp 1669390400
transform 1 0 61152 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_540
timestamp 1669390400
transform 1 0 61824 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_544
timestamp 1669390400
transform 1 0 62272 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_550
timestamp 1669390400
transform 1 0 62944 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_558
timestamp 1669390400
transform 1 0 63840 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_590
timestamp 1669390400
transform 1 0 67424 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_598
timestamp 1669390400
transform 1 0 68320 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_602
timestamp 1669390400
transform 1 0 68768 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_605
timestamp 1669390400
transform 1 0 69104 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_637
timestamp 1669390400
transform 1 0 72688 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_653
timestamp 1669390400
transform 1 0 74480 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_655
timestamp 1669390400
transform 1 0 74704 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_672
timestamp 1669390400
transform 1 0 76608 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_676
timestamp 1669390400
transform 1 0 77056 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_679
timestamp 1669390400
transform 1 0 77392 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_687
timestamp 1669390400
transform 1 0 78288 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_2
timestamp 1669390400
transform 1 0 1568 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_19
timestamp 1669390400
transform 1 0 3472 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_23
timestamp 1669390400
transform 1 0 3920 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_55
timestamp 1669390400
transform 1 0 7504 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_73
timestamp 1669390400
transform 1 0 9520 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_137
timestamp 1669390400
transform 1 0 16688 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_141
timestamp 1669390400
transform 1 0 17136 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_144
timestamp 1669390400
transform 1 0 17472 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_208
timestamp 1669390400
transform 1 0 24640 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_212
timestamp 1669390400
transform 1 0 25088 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_215
timestamp 1669390400
transform 1 0 25424 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_279
timestamp 1669390400
transform 1 0 32592 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_283
timestamp 1669390400
transform 1 0 33040 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_286
timestamp 1669390400
transform 1 0 33376 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_350
timestamp 1669390400
transform 1 0 40544 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_354
timestamp 1669390400
transform 1 0 40992 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_357
timestamp 1669390400
transform 1 0 41328 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_421
timestamp 1669390400
transform 1 0 48496 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_425
timestamp 1669390400
transform 1 0 48944 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_428
timestamp 1669390400
transform 1 0 49280 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_492
timestamp 1669390400
transform 1 0 56448 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_496
timestamp 1669390400
transform 1 0 56896 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_499
timestamp 1669390400
transform 1 0 57232 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_515
timestamp 1669390400
transform 1 0 59024 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_523
timestamp 1669390400
transform 1 0 59920 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_527
timestamp 1669390400
transform 1 0 60368 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_531
timestamp 1669390400
transform 1 0 60816 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_535
timestamp 1669390400
transform 1 0 61264 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_541
timestamp 1669390400
transform 1 0 61936 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_553
timestamp 1669390400
transform 1 0 63280 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_565
timestamp 1669390400
transform 1 0 64624 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_567
timestamp 1669390400
transform 1 0 64848 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_570
timestamp 1669390400
transform 1 0 65184 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_586
timestamp 1669390400
transform 1 0 66976 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_594
timestamp 1669390400
transform 1 0 67872 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_599
timestamp 1669390400
transform 1 0 68432 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_603
timestamp 1669390400
transform 1 0 68880 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_635
timestamp 1669390400
transform 1 0 72464 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_641
timestamp 1669390400
transform 1 0 73136 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_649
timestamp 1669390400
transform 1 0 74032 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_653
timestamp 1669390400
transform 1 0 74480 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_655
timestamp 1669390400
transform 1 0 74704 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_672
timestamp 1669390400
transform 1 0 76608 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_676
timestamp 1669390400
transform 1 0 77056 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_684
timestamp 1669390400
transform 1 0 77952 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_2
timestamp 1669390400
transform 1 0 1568 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_19
timestamp 1669390400
transform 1 0 3472 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_23
timestamp 1669390400
transform 1 0 3920 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_27
timestamp 1669390400
transform 1 0 4368 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_37
timestamp 1669390400
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_101
timestamp 1669390400
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_105
timestamp 1669390400
transform 1 0 13104 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_108
timestamp 1669390400
transform 1 0 13440 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_172
timestamp 1669390400
transform 1 0 20608 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_176
timestamp 1669390400
transform 1 0 21056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_179
timestamp 1669390400
transform 1 0 21392 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_243
timestamp 1669390400
transform 1 0 28560 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_247
timestamp 1669390400
transform 1 0 29008 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_250
timestamp 1669390400
transform 1 0 29344 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_314
timestamp 1669390400
transform 1 0 36512 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_318
timestamp 1669390400
transform 1 0 36960 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_321
timestamp 1669390400
transform 1 0 37296 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_385
timestamp 1669390400
transform 1 0 44464 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_389
timestamp 1669390400
transform 1 0 44912 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_392
timestamp 1669390400
transform 1 0 45248 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_456
timestamp 1669390400
transform 1 0 52416 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_460
timestamp 1669390400
transform 1 0 52864 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_463
timestamp 1669390400
transform 1 0 53200 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_495
timestamp 1669390400
transform 1 0 56784 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_511
timestamp 1669390400
transform 1 0 58576 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_515
timestamp 1669390400
transform 1 0 59024 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_520
timestamp 1669390400
transform 1 0 59584 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_524
timestamp 1669390400
transform 1 0 60032 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_534
timestamp 1669390400
transform 1 0 61152 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_539
timestamp 1669390400
transform 1 0 61712 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_543
timestamp 1669390400
transform 1 0 62160 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_547
timestamp 1669390400
transform 1 0 62608 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_549
timestamp 1669390400
transform 1 0 62832 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_560
timestamp 1669390400
transform 1 0 64064 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_564
timestamp 1669390400
transform 1 0 64512 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_566
timestamp 1669390400
transform 1 0 64736 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_569
timestamp 1669390400
transform 1 0 65072 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_573
timestamp 1669390400
transform 1 0 65520 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_579
timestamp 1669390400
transform 1 0 66192 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_583
timestamp 1669390400
transform 1 0 66640 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_585
timestamp 1669390400
transform 1 0 66864 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_588
timestamp 1669390400
transform 1 0 67200 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_596
timestamp 1669390400
transform 1 0 68096 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_600
timestamp 1669390400
transform 1 0 68544 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_602
timestamp 1669390400
transform 1 0 68768 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_605
timestamp 1669390400
transform 1 0 69104 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_637
timestamp 1669390400
transform 1 0 72688 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_653
timestamp 1669390400
transform 1 0 74480 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_655
timestamp 1669390400
transform 1 0 74704 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_672
timestamp 1669390400
transform 1 0 76608 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_676
timestamp 1669390400
transform 1 0 77056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_679
timestamp 1669390400
transform 1 0 77392 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_687
timestamp 1669390400
transform 1 0 78288 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_2
timestamp 1669390400
transform 1 0 1568 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_19
timestamp 1669390400
transform 1 0 3472 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_37
timestamp 1669390400
transform 1 0 5488 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_69
timestamp 1669390400
transform 1 0 9072 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_73
timestamp 1669390400
transform 1 0 9520 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_137
timestamp 1669390400
transform 1 0 16688 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_141
timestamp 1669390400
transform 1 0 17136 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_144
timestamp 1669390400
transform 1 0 17472 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_208
timestamp 1669390400
transform 1 0 24640 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_212
timestamp 1669390400
transform 1 0 25088 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_215
timestamp 1669390400
transform 1 0 25424 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_279
timestamp 1669390400
transform 1 0 32592 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_283
timestamp 1669390400
transform 1 0 33040 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_286
timestamp 1669390400
transform 1 0 33376 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_350
timestamp 1669390400
transform 1 0 40544 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_354
timestamp 1669390400
transform 1 0 40992 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_357
timestamp 1669390400
transform 1 0 41328 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_421
timestamp 1669390400
transform 1 0 48496 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_425
timestamp 1669390400
transform 1 0 48944 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_428
timestamp 1669390400
transform 1 0 49280 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_492
timestamp 1669390400
transform 1 0 56448 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_496
timestamp 1669390400
transform 1 0 56896 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_499
timestamp 1669390400
transform 1 0 57232 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_531
timestamp 1669390400
transform 1 0 60816 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_536
timestamp 1669390400
transform 1 0 61376 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_540
timestamp 1669390400
transform 1 0 61824 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_548
timestamp 1669390400
transform 1 0 62720 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_550
timestamp 1669390400
transform 1 0 62944 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_561
timestamp 1669390400
transform 1 0 64176 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_567
timestamp 1669390400
transform 1 0 64848 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_570
timestamp 1669390400
transform 1 0 65184 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_577
timestamp 1669390400
transform 1 0 65968 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_585
timestamp 1669390400
transform 1 0 66864 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_587
timestamp 1669390400
transform 1 0 67088 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_594
timestamp 1669390400
transform 1 0 67872 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_626
timestamp 1669390400
transform 1 0 71456 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_634
timestamp 1669390400
transform 1 0 72352 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_638
timestamp 1669390400
transform 1 0 72800 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_641
timestamp 1669390400
transform 1 0 73136 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_649
timestamp 1669390400
transform 1 0 74032 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_651
timestamp 1669390400
transform 1 0 74256 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_654
timestamp 1669390400
transform 1 0 74592 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_672
timestamp 1669390400
transform 1 0 76608 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_676
timestamp 1669390400
transform 1 0 77056 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_684
timestamp 1669390400
transform 1 0 77952 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_2
timestamp 1669390400
transform 1 0 1568 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_19
timestamp 1669390400
transform 1 0 3472 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_23
timestamp 1669390400
transform 1 0 3920 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_27
timestamp 1669390400
transform 1 0 4368 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_37
timestamp 1669390400
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_101
timestamp 1669390400
transform 1 0 12656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_105
timestamp 1669390400
transform 1 0 13104 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_108
timestamp 1669390400
transform 1 0 13440 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_172
timestamp 1669390400
transform 1 0 20608 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_176
timestamp 1669390400
transform 1 0 21056 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_179
timestamp 1669390400
transform 1 0 21392 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_243
timestamp 1669390400
transform 1 0 28560 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_247
timestamp 1669390400
transform 1 0 29008 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_250
timestamp 1669390400
transform 1 0 29344 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_314
timestamp 1669390400
transform 1 0 36512 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_318
timestamp 1669390400
transform 1 0 36960 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_321
timestamp 1669390400
transform 1 0 37296 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_385
timestamp 1669390400
transform 1 0 44464 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_389
timestamp 1669390400
transform 1 0 44912 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_392
timestamp 1669390400
transform 1 0 45248 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_456
timestamp 1669390400
transform 1 0 52416 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_460
timestamp 1669390400
transform 1 0 52864 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_463
timestamp 1669390400
transform 1 0 53200 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_527
timestamp 1669390400
transform 1 0 60368 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_531
timestamp 1669390400
transform 1 0 60816 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_534
timestamp 1669390400
transform 1 0 61152 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_542
timestamp 1669390400
transform 1 0 62048 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_546
timestamp 1669390400
transform 1 0 62496 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_554
timestamp 1669390400
transform 1 0 63392 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_558
timestamp 1669390400
transform 1 0 63840 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_564
timestamp 1669390400
transform 1 0 64512 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_566
timestamp 1669390400
transform 1 0 64736 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_577
timestamp 1669390400
transform 1 0 65968 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_583
timestamp 1669390400
transform 1 0 66640 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_591
timestamp 1669390400
transform 1 0 67536 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_595
timestamp 1669390400
transform 1 0 67984 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_602
timestamp 1669390400
transform 1 0 68768 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_605
timestamp 1669390400
transform 1 0 69104 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_612
timestamp 1669390400
transform 1 0 69888 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_628
timestamp 1669390400
transform 1 0 71680 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_636
timestamp 1669390400
transform 1 0 72576 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_654
timestamp 1669390400
transform 1 0 74592 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_672
timestamp 1669390400
transform 1 0 76608 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_676
timestamp 1669390400
transform 1 0 77056 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_679
timestamp 1669390400
transform 1 0 77392 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_687
timestamp 1669390400
transform 1 0 78288 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_2
timestamp 1669390400
transform 1 0 1568 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_19
timestamp 1669390400
transform 1 0 3472 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_23
timestamp 1669390400
transform 1 0 3920 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_55
timestamp 1669390400
transform 1 0 7504 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_73
timestamp 1669390400
transform 1 0 9520 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_137
timestamp 1669390400
transform 1 0 16688 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_141
timestamp 1669390400
transform 1 0 17136 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_144
timestamp 1669390400
transform 1 0 17472 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_208
timestamp 1669390400
transform 1 0 24640 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_212
timestamp 1669390400
transform 1 0 25088 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_215
timestamp 1669390400
transform 1 0 25424 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_279
timestamp 1669390400
transform 1 0 32592 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_283
timestamp 1669390400
transform 1 0 33040 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_286
timestamp 1669390400
transform 1 0 33376 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_350
timestamp 1669390400
transform 1 0 40544 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_354
timestamp 1669390400
transform 1 0 40992 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_357
timestamp 1669390400
transform 1 0 41328 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_421
timestamp 1669390400
transform 1 0 48496 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_425
timestamp 1669390400
transform 1 0 48944 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_428
timestamp 1669390400
transform 1 0 49280 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_492
timestamp 1669390400
transform 1 0 56448 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_496
timestamp 1669390400
transform 1 0 56896 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_499
timestamp 1669390400
transform 1 0 57232 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_531
timestamp 1669390400
transform 1 0 60816 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_539
timestamp 1669390400
transform 1 0 61712 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_544
timestamp 1669390400
transform 1 0 62272 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_548
timestamp 1669390400
transform 1 0 62720 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_556
timestamp 1669390400
transform 1 0 63616 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_560
timestamp 1669390400
transform 1 0 64064 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_562
timestamp 1669390400
transform 1 0 64288 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_567
timestamp 1669390400
transform 1 0 64848 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_570
timestamp 1669390400
transform 1 0 65184 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_581
timestamp 1669390400
transform 1 0 66416 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_585
timestamp 1669390400
transform 1 0 66864 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_589
timestamp 1669390400
transform 1 0 67312 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_603
timestamp 1669390400
transform 1 0 68880 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_635
timestamp 1669390400
transform 1 0 72464 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_641
timestamp 1669390400
transform 1 0 73136 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_649
timestamp 1669390400
transform 1 0 74032 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_653
timestamp 1669390400
transform 1 0 74480 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_655
timestamp 1669390400
transform 1 0 74704 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_672
timestamp 1669390400
transform 1 0 76608 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_676
timestamp 1669390400
transform 1 0 77056 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_684
timestamp 1669390400
transform 1 0 77952 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_2
timestamp 1669390400
transform 1 0 1568 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_19
timestamp 1669390400
transform 1 0 3472 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_23
timestamp 1669390400
transform 1 0 3920 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_31
timestamp 1669390400
transform 1 0 4816 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_37
timestamp 1669390400
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_101
timestamp 1669390400
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_105
timestamp 1669390400
transform 1 0 13104 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_108
timestamp 1669390400
transform 1 0 13440 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_172
timestamp 1669390400
transform 1 0 20608 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_176
timestamp 1669390400
transform 1 0 21056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_179
timestamp 1669390400
transform 1 0 21392 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_243
timestamp 1669390400
transform 1 0 28560 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_247
timestamp 1669390400
transform 1 0 29008 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_250
timestamp 1669390400
transform 1 0 29344 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_314
timestamp 1669390400
transform 1 0 36512 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_318
timestamp 1669390400
transform 1 0 36960 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_321
timestamp 1669390400
transform 1 0 37296 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_385
timestamp 1669390400
transform 1 0 44464 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_389
timestamp 1669390400
transform 1 0 44912 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_392
timestamp 1669390400
transform 1 0 45248 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_456
timestamp 1669390400
transform 1 0 52416 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_460
timestamp 1669390400
transform 1 0 52864 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_463
timestamp 1669390400
transform 1 0 53200 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_527
timestamp 1669390400
transform 1 0 60368 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_531
timestamp 1669390400
transform 1 0 60816 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_80_534
timestamp 1669390400
transform 1 0 61152 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_550
timestamp 1669390400
transform 1 0 62944 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_556
timestamp 1669390400
transform 1 0 63616 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_560
timestamp 1669390400
transform 1 0 64064 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_564
timestamp 1669390400
transform 1 0 64512 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_566
timestamp 1669390400
transform 1 0 64736 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_569
timestamp 1669390400
transform 1 0 65072 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_581
timestamp 1669390400
transform 1 0 66416 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_587
timestamp 1669390400
transform 1 0 67088 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_589
timestamp 1669390400
transform 1 0 67312 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_600
timestamp 1669390400
transform 1 0 68544 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_602
timestamp 1669390400
transform 1 0 68768 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_605
timestamp 1669390400
transform 1 0 69104 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_80_637
timestamp 1669390400
transform 1 0 72688 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_653
timestamp 1669390400
transform 1 0 74480 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_655
timestamp 1669390400
transform 1 0 74704 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_672
timestamp 1669390400
transform 1 0 76608 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_676
timestamp 1669390400
transform 1 0 77056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_679
timestamp 1669390400
transform 1 0 77392 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_687
timestamp 1669390400
transform 1 0 78288 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_2
timestamp 1669390400
transform 1 0 1568 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_19
timestamp 1669390400
transform 1 0 3472 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_23
timestamp 1669390400
transform 1 0 3920 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_55
timestamp 1669390400
transform 1 0 7504 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_73
timestamp 1669390400
transform 1 0 9520 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_137
timestamp 1669390400
transform 1 0 16688 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_141
timestamp 1669390400
transform 1 0 17136 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_144
timestamp 1669390400
transform 1 0 17472 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_208
timestamp 1669390400
transform 1 0 24640 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_212
timestamp 1669390400
transform 1 0 25088 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_215
timestamp 1669390400
transform 1 0 25424 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_279
timestamp 1669390400
transform 1 0 32592 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_283
timestamp 1669390400
transform 1 0 33040 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_286
timestamp 1669390400
transform 1 0 33376 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_350
timestamp 1669390400
transform 1 0 40544 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_354
timestamp 1669390400
transform 1 0 40992 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_357
timestamp 1669390400
transform 1 0 41328 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_421
timestamp 1669390400
transform 1 0 48496 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_425
timestamp 1669390400
transform 1 0 48944 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_428
timestamp 1669390400
transform 1 0 49280 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_492
timestamp 1669390400
transform 1 0 56448 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_496
timestamp 1669390400
transform 1 0 56896 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_499
timestamp 1669390400
transform 1 0 57232 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_531
timestamp 1669390400
transform 1 0 60816 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_547
timestamp 1669390400
transform 1 0 62608 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_551
timestamp 1669390400
transform 1 0 63056 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_557
timestamp 1669390400
transform 1 0 63728 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_561
timestamp 1669390400
transform 1 0 64176 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_565
timestamp 1669390400
transform 1 0 64624 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_567
timestamp 1669390400
transform 1 0 64848 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_570
timestamp 1669390400
transform 1 0 65184 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_582
timestamp 1669390400
transform 1 0 66528 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_588
timestamp 1669390400
transform 1 0 67200 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_592
timestamp 1669390400
transform 1 0 67648 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_604
timestamp 1669390400
transform 1 0 68992 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_610
timestamp 1669390400
transform 1 0 69664 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_626
timestamp 1669390400
transform 1 0 71456 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_634
timestamp 1669390400
transform 1 0 72352 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_638
timestamp 1669390400
transform 1 0 72800 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_641
timestamp 1669390400
transform 1 0 73136 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_649
timestamp 1669390400
transform 1 0 74032 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_653
timestamp 1669390400
transform 1 0 74480 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_655
timestamp 1669390400
transform 1 0 74704 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_672
timestamp 1669390400
transform 1 0 76608 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_676
timestamp 1669390400
transform 1 0 77056 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_684
timestamp 1669390400
transform 1 0 77952 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_2
timestamp 1669390400
transform 1 0 1568 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_19
timestamp 1669390400
transform 1 0 3472 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_23
timestamp 1669390400
transform 1 0 3920 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_27
timestamp 1669390400
transform 1 0 4368 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_37
timestamp 1669390400
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_101
timestamp 1669390400
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_105
timestamp 1669390400
transform 1 0 13104 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_108
timestamp 1669390400
transform 1 0 13440 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_172
timestamp 1669390400
transform 1 0 20608 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_176
timestamp 1669390400
transform 1 0 21056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_179
timestamp 1669390400
transform 1 0 21392 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_243
timestamp 1669390400
transform 1 0 28560 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_247
timestamp 1669390400
transform 1 0 29008 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_250
timestamp 1669390400
transform 1 0 29344 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_314
timestamp 1669390400
transform 1 0 36512 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_318
timestamp 1669390400
transform 1 0 36960 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_321
timestamp 1669390400
transform 1 0 37296 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_385
timestamp 1669390400
transform 1 0 44464 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_389
timestamp 1669390400
transform 1 0 44912 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_392
timestamp 1669390400
transform 1 0 45248 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_456
timestamp 1669390400
transform 1 0 52416 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_460
timestamp 1669390400
transform 1 0 52864 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_463
timestamp 1669390400
transform 1 0 53200 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_527
timestamp 1669390400
transform 1 0 60368 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_531
timestamp 1669390400
transform 1 0 60816 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_534
timestamp 1669390400
transform 1 0 61152 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_566
timestamp 1669390400
transform 1 0 64736 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_574
timestamp 1669390400
transform 1 0 65632 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_578
timestamp 1669390400
transform 1 0 66080 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_581
timestamp 1669390400
transform 1 0 66416 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_585
timestamp 1669390400
transform 1 0 66864 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_591
timestamp 1669390400
transform 1 0 67536 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_597
timestamp 1669390400
transform 1 0 68208 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_601
timestamp 1669390400
transform 1 0 68656 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_605
timestamp 1669390400
transform 1 0 69104 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_610
timestamp 1669390400
transform 1 0 69664 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_642
timestamp 1669390400
transform 1 0 73248 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_650
timestamp 1669390400
transform 1 0 74144 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_654
timestamp 1669390400
transform 1 0 74592 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_672
timestamp 1669390400
transform 1 0 76608 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_676
timestamp 1669390400
transform 1 0 77056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_679
timestamp 1669390400
transform 1 0 77392 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_687
timestamp 1669390400
transform 1 0 78288 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_2
timestamp 1669390400
transform 1 0 1568 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_19
timestamp 1669390400
transform 1 0 3472 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_37
timestamp 1669390400
transform 1 0 5488 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_69
timestamp 1669390400
transform 1 0 9072 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_73
timestamp 1669390400
transform 1 0 9520 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_137
timestamp 1669390400
transform 1 0 16688 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_141
timestamp 1669390400
transform 1 0 17136 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_144
timestamp 1669390400
transform 1 0 17472 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_208
timestamp 1669390400
transform 1 0 24640 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_212
timestamp 1669390400
transform 1 0 25088 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_215
timestamp 1669390400
transform 1 0 25424 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_279
timestamp 1669390400
transform 1 0 32592 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_283
timestamp 1669390400
transform 1 0 33040 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_286
timestamp 1669390400
transform 1 0 33376 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_350
timestamp 1669390400
transform 1 0 40544 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_354
timestamp 1669390400
transform 1 0 40992 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_357
timestamp 1669390400
transform 1 0 41328 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_421
timestamp 1669390400
transform 1 0 48496 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_425
timestamp 1669390400
transform 1 0 48944 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_428
timestamp 1669390400
transform 1 0 49280 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_492
timestamp 1669390400
transform 1 0 56448 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_496
timestamp 1669390400
transform 1 0 56896 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_499
timestamp 1669390400
transform 1 0 57232 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_563
timestamp 1669390400
transform 1 0 64400 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_567
timestamp 1669390400
transform 1 0 64848 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_570
timestamp 1669390400
transform 1 0 65184 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_586
timestamp 1669390400
transform 1 0 66976 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_589
timestamp 1669390400
transform 1 0 67312 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_595
timestamp 1669390400
transform 1 0 67984 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_603
timestamp 1669390400
transform 1 0 68880 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_611
timestamp 1669390400
transform 1 0 69776 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_614
timestamp 1669390400
transform 1 0 70112 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_630
timestamp 1669390400
transform 1 0 71904 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_638
timestamp 1669390400
transform 1 0 72800 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_641
timestamp 1669390400
transform 1 0 73136 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_649
timestamp 1669390400
transform 1 0 74032 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_651
timestamp 1669390400
transform 1 0 74256 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_654
timestamp 1669390400
transform 1 0 74592 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_672
timestamp 1669390400
transform 1 0 76608 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_676
timestamp 1669390400
transform 1 0 77056 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_684
timestamp 1669390400
transform 1 0 77952 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_2
timestamp 1669390400
transform 1 0 1568 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_19
timestamp 1669390400
transform 1 0 3472 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_23
timestamp 1669390400
transform 1 0 3920 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_27
timestamp 1669390400
transform 1 0 4368 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_37
timestamp 1669390400
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_101
timestamp 1669390400
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_105
timestamp 1669390400
transform 1 0 13104 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_108
timestamp 1669390400
transform 1 0 13440 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_172
timestamp 1669390400
transform 1 0 20608 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_176
timestamp 1669390400
transform 1 0 21056 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_179
timestamp 1669390400
transform 1 0 21392 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_243
timestamp 1669390400
transform 1 0 28560 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_247
timestamp 1669390400
transform 1 0 29008 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_250
timestamp 1669390400
transform 1 0 29344 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_314
timestamp 1669390400
transform 1 0 36512 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_318
timestamp 1669390400
transform 1 0 36960 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_321
timestamp 1669390400
transform 1 0 37296 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_385
timestamp 1669390400
transform 1 0 44464 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_389
timestamp 1669390400
transform 1 0 44912 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_392
timestamp 1669390400
transform 1 0 45248 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_456
timestamp 1669390400
transform 1 0 52416 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_460
timestamp 1669390400
transform 1 0 52864 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_463
timestamp 1669390400
transform 1 0 53200 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_527
timestamp 1669390400
transform 1 0 60368 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_531
timestamp 1669390400
transform 1 0 60816 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_534
timestamp 1669390400
transform 1 0 61152 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_598
timestamp 1669390400
transform 1 0 68320 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_602
timestamp 1669390400
transform 1 0 68768 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_605
timestamp 1669390400
transform 1 0 69104 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_612
timestamp 1669390400
transform 1 0 69888 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_620
timestamp 1669390400
transform 1 0 70784 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_624
timestamp 1669390400
transform 1 0 71232 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_632
timestamp 1669390400
transform 1 0 72128 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_636
timestamp 1669390400
transform 1 0 72576 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_654
timestamp 1669390400
transform 1 0 74592 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_672
timestamp 1669390400
transform 1 0 76608 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_676
timestamp 1669390400
transform 1 0 77056 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_679
timestamp 1669390400
transform 1 0 77392 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_687
timestamp 1669390400
transform 1 0 78288 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_2
timestamp 1669390400
transform 1 0 1568 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_19
timestamp 1669390400
transform 1 0 3472 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_23
timestamp 1669390400
transform 1 0 3920 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_85_55
timestamp 1669390400
transform 1 0 7504 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_73
timestamp 1669390400
transform 1 0 9520 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_137
timestamp 1669390400
transform 1 0 16688 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_141
timestamp 1669390400
transform 1 0 17136 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_144
timestamp 1669390400
transform 1 0 17472 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_208
timestamp 1669390400
transform 1 0 24640 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_212
timestamp 1669390400
transform 1 0 25088 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_215
timestamp 1669390400
transform 1 0 25424 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_279
timestamp 1669390400
transform 1 0 32592 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_283
timestamp 1669390400
transform 1 0 33040 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_286
timestamp 1669390400
transform 1 0 33376 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_350
timestamp 1669390400
transform 1 0 40544 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_354
timestamp 1669390400
transform 1 0 40992 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_357
timestamp 1669390400
transform 1 0 41328 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_421
timestamp 1669390400
transform 1 0 48496 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_425
timestamp 1669390400
transform 1 0 48944 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_428
timestamp 1669390400
transform 1 0 49280 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_492
timestamp 1669390400
transform 1 0 56448 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_496
timestamp 1669390400
transform 1 0 56896 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_499
timestamp 1669390400
transform 1 0 57232 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_563
timestamp 1669390400
transform 1 0 64400 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_567
timestamp 1669390400
transform 1 0 64848 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_570
timestamp 1669390400
transform 1 0 65184 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_602
timestamp 1669390400
transform 1 0 68768 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_606
timestamp 1669390400
transform 1 0 69216 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_609
timestamp 1669390400
transform 1 0 69552 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_617
timestamp 1669390400
transform 1 0 70448 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_619
timestamp 1669390400
transform 1 0 70672 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_626
timestamp 1669390400
transform 1 0 71456 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_630
timestamp 1669390400
transform 1 0 71904 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_638
timestamp 1669390400
transform 1 0 72800 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_641
timestamp 1669390400
transform 1 0 73136 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_649
timestamp 1669390400
transform 1 0 74032 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_653
timestamp 1669390400
transform 1 0 74480 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_655
timestamp 1669390400
transform 1 0 74704 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_672
timestamp 1669390400
transform 1 0 76608 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_676
timestamp 1669390400
transform 1 0 77056 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_684
timestamp 1669390400
transform 1 0 77952 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_2
timestamp 1669390400
transform 1 0 1568 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_19
timestamp 1669390400
transform 1 0 3472 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_23
timestamp 1669390400
transform 1 0 3920 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_31
timestamp 1669390400
transform 1 0 4816 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_37
timestamp 1669390400
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_101
timestamp 1669390400
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_105
timestamp 1669390400
transform 1 0 13104 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_108
timestamp 1669390400
transform 1 0 13440 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_172
timestamp 1669390400
transform 1 0 20608 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_176
timestamp 1669390400
transform 1 0 21056 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_179
timestamp 1669390400
transform 1 0 21392 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_243
timestamp 1669390400
transform 1 0 28560 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_247
timestamp 1669390400
transform 1 0 29008 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_250
timestamp 1669390400
transform 1 0 29344 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_314
timestamp 1669390400
transform 1 0 36512 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_318
timestamp 1669390400
transform 1 0 36960 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_321
timestamp 1669390400
transform 1 0 37296 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_385
timestamp 1669390400
transform 1 0 44464 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_389
timestamp 1669390400
transform 1 0 44912 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_392
timestamp 1669390400
transform 1 0 45248 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_456
timestamp 1669390400
transform 1 0 52416 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_460
timestamp 1669390400
transform 1 0 52864 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_463
timestamp 1669390400
transform 1 0 53200 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_527
timestamp 1669390400
transform 1 0 60368 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_531
timestamp 1669390400
transform 1 0 60816 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_534
timestamp 1669390400
transform 1 0 61152 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_598
timestamp 1669390400
transform 1 0 68320 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_602
timestamp 1669390400
transform 1 0 68768 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_605
timestamp 1669390400
transform 1 0 69104 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_615
timestamp 1669390400
transform 1 0 70224 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_623
timestamp 1669390400
transform 1 0 71120 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_625
timestamp 1669390400
transform 1 0 71344 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_632
timestamp 1669390400
transform 1 0 72128 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_636
timestamp 1669390400
transform 1 0 72576 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_640
timestamp 1669390400
transform 1 0 73024 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_644
timestamp 1669390400
transform 1 0 73472 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_648
timestamp 1669390400
transform 1 0 73920 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_654
timestamp 1669390400
transform 1 0 74592 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_672
timestamp 1669390400
transform 1 0 76608 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_676
timestamp 1669390400
transform 1 0 77056 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_679
timestamp 1669390400
transform 1 0 77392 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_687
timestamp 1669390400
transform 1 0 78288 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_2
timestamp 1669390400
transform 1 0 1568 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_17
timestamp 1669390400
transform 1 0 3248 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_33
timestamp 1669390400
transform 1 0 5040 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_37
timestamp 1669390400
transform 1 0 5488 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_69
timestamp 1669390400
transform 1 0 9072 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_73
timestamp 1669390400
transform 1 0 9520 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_137
timestamp 1669390400
transform 1 0 16688 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_141
timestamp 1669390400
transform 1 0 17136 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_144
timestamp 1669390400
transform 1 0 17472 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_208
timestamp 1669390400
transform 1 0 24640 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_212
timestamp 1669390400
transform 1 0 25088 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_215
timestamp 1669390400
transform 1 0 25424 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_279
timestamp 1669390400
transform 1 0 32592 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_283
timestamp 1669390400
transform 1 0 33040 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_286
timestamp 1669390400
transform 1 0 33376 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_350
timestamp 1669390400
transform 1 0 40544 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_354
timestamp 1669390400
transform 1 0 40992 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_357
timestamp 1669390400
transform 1 0 41328 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_421
timestamp 1669390400
transform 1 0 48496 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_425
timestamp 1669390400
transform 1 0 48944 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_428
timestamp 1669390400
transform 1 0 49280 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_492
timestamp 1669390400
transform 1 0 56448 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_496
timestamp 1669390400
transform 1 0 56896 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_499
timestamp 1669390400
transform 1 0 57232 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_563
timestamp 1669390400
transform 1 0 64400 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_567
timestamp 1669390400
transform 1 0 64848 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_570
timestamp 1669390400
transform 1 0 65184 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_87_602
timestamp 1669390400
transform 1 0 68768 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_618
timestamp 1669390400
transform 1 0 70560 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_621
timestamp 1669390400
transform 1 0 70896 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_629
timestamp 1669390400
transform 1 0 71792 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_637
timestamp 1669390400
transform 1 0 72688 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_641
timestamp 1669390400
transform 1 0 73136 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_646
timestamp 1669390400
transform 1 0 73696 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_652
timestamp 1669390400
transform 1 0 74368 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_670
timestamp 1669390400
transform 1 0 76384 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_686
timestamp 1669390400
transform 1 0 78176 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_2
timestamp 1669390400
transform 1 0 1568 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_17
timestamp 1669390400
transform 1 0 3248 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_21
timestamp 1669390400
transform 1 0 3696 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_25
timestamp 1669390400
transform 1 0 4144 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_33
timestamp 1669390400
transform 1 0 5040 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_37
timestamp 1669390400
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_101
timestamp 1669390400
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_105
timestamp 1669390400
transform 1 0 13104 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_108
timestamp 1669390400
transform 1 0 13440 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_172
timestamp 1669390400
transform 1 0 20608 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_176
timestamp 1669390400
transform 1 0 21056 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_179
timestamp 1669390400
transform 1 0 21392 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_243
timestamp 1669390400
transform 1 0 28560 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_247
timestamp 1669390400
transform 1 0 29008 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_250
timestamp 1669390400
transform 1 0 29344 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_314
timestamp 1669390400
transform 1 0 36512 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_318
timestamp 1669390400
transform 1 0 36960 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_321
timestamp 1669390400
transform 1 0 37296 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_385
timestamp 1669390400
transform 1 0 44464 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_389
timestamp 1669390400
transform 1 0 44912 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_392
timestamp 1669390400
transform 1 0 45248 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_456
timestamp 1669390400
transform 1 0 52416 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_460
timestamp 1669390400
transform 1 0 52864 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_463
timestamp 1669390400
transform 1 0 53200 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_527
timestamp 1669390400
transform 1 0 60368 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_531
timestamp 1669390400
transform 1 0 60816 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_534
timestamp 1669390400
transform 1 0 61152 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_598
timestamp 1669390400
transform 1 0 68320 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_602
timestamp 1669390400
transform 1 0 68768 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_605
timestamp 1669390400
transform 1 0 69104 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_612
timestamp 1669390400
transform 1 0 69888 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_616
timestamp 1669390400
transform 1 0 70336 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_624
timestamp 1669390400
transform 1 0 71232 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_634
timestamp 1669390400
transform 1 0 72352 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_644
timestamp 1669390400
transform 1 0 73472 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_652
timestamp 1669390400
transform 1 0 74368 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_670
timestamp 1669390400
transform 1 0 76384 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_676
timestamp 1669390400
transform 1 0 77056 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_684
timestamp 1669390400
transform 1 0 77952 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_2
timestamp 1669390400
transform 1 0 1568 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_17
timestamp 1669390400
transform 1 0 3248 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_33
timestamp 1669390400
transform 1 0 5040 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_89_37
timestamp 1669390400
transform 1 0 5488 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_69
timestamp 1669390400
transform 1 0 9072 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_73
timestamp 1669390400
transform 1 0 9520 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_137
timestamp 1669390400
transform 1 0 16688 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_141
timestamp 1669390400
transform 1 0 17136 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_144
timestamp 1669390400
transform 1 0 17472 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_208
timestamp 1669390400
transform 1 0 24640 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_212
timestamp 1669390400
transform 1 0 25088 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_215
timestamp 1669390400
transform 1 0 25424 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_279
timestamp 1669390400
transform 1 0 32592 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_283
timestamp 1669390400
transform 1 0 33040 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_286
timestamp 1669390400
transform 1 0 33376 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_350
timestamp 1669390400
transform 1 0 40544 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_354
timestamp 1669390400
transform 1 0 40992 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_357
timestamp 1669390400
transform 1 0 41328 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_421
timestamp 1669390400
transform 1 0 48496 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_425
timestamp 1669390400
transform 1 0 48944 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_428
timestamp 1669390400
transform 1 0 49280 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_492
timestamp 1669390400
transform 1 0 56448 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_496
timestamp 1669390400
transform 1 0 56896 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_499
timestamp 1669390400
transform 1 0 57232 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_563
timestamp 1669390400
transform 1 0 64400 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_567
timestamp 1669390400
transform 1 0 64848 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_570
timestamp 1669390400
transform 1 0 65184 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_89_586
timestamp 1669390400
transform 1 0 66976 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_594
timestamp 1669390400
transform 1 0 67872 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_598
timestamp 1669390400
transform 1 0 68320 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_600
timestamp 1669390400
transform 1 0 68544 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_607
timestamp 1669390400
transform 1 0 69328 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_611
timestamp 1669390400
transform 1 0 69776 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_627
timestamp 1669390400
transform 1 0 71568 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_631
timestamp 1669390400
transform 1 0 72016 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_633
timestamp 1669390400
transform 1 0 72240 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_636
timestamp 1669390400
transform 1 0 72576 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_638
timestamp 1669390400
transform 1 0 72800 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_641
timestamp 1669390400
transform 1 0 73136 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_643
timestamp 1669390400
transform 1 0 73360 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_650
timestamp 1669390400
transform 1 0 74144 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_654
timestamp 1669390400
transform 1 0 74592 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_670
timestamp 1669390400
transform 1 0 76384 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_686
timestamp 1669390400
transform 1 0 78176 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_2
timestamp 1669390400
transform 1 0 1568 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_19
timestamp 1669390400
transform 1 0 3472 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_23
timestamp 1669390400
transform 1 0 3920 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_27
timestamp 1669390400
transform 1 0 4368 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_37
timestamp 1669390400
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_101
timestamp 1669390400
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_105
timestamp 1669390400
transform 1 0 13104 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_108
timestamp 1669390400
transform 1 0 13440 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_172
timestamp 1669390400
transform 1 0 20608 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_176
timestamp 1669390400
transform 1 0 21056 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_179
timestamp 1669390400
transform 1 0 21392 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_243
timestamp 1669390400
transform 1 0 28560 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_247
timestamp 1669390400
transform 1 0 29008 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_250
timestamp 1669390400
transform 1 0 29344 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_314
timestamp 1669390400
transform 1 0 36512 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_318
timestamp 1669390400
transform 1 0 36960 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_321
timestamp 1669390400
transform 1 0 37296 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_385
timestamp 1669390400
transform 1 0 44464 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_389
timestamp 1669390400
transform 1 0 44912 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_392
timestamp 1669390400
transform 1 0 45248 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_456
timestamp 1669390400
transform 1 0 52416 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_460
timestamp 1669390400
transform 1 0 52864 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_463
timestamp 1669390400
transform 1 0 53200 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_527
timestamp 1669390400
transform 1 0 60368 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_531
timestamp 1669390400
transform 1 0 60816 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_534
timestamp 1669390400
transform 1 0 61152 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_598
timestamp 1669390400
transform 1 0 68320 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_602
timestamp 1669390400
transform 1 0 68768 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_605
timestamp 1669390400
transform 1 0 69104 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_637
timestamp 1669390400
transform 1 0 72688 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_641
timestamp 1669390400
transform 1 0 73136 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_643
timestamp 1669390400
transform 1 0 73360 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_646
timestamp 1669390400
transform 1 0 73696 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_650
timestamp 1669390400
transform 1 0 74144 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_654
timestamp 1669390400
transform 1 0 74592 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_672
timestamp 1669390400
transform 1 0 76608 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_676
timestamp 1669390400
transform 1 0 77056 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_679
timestamp 1669390400
transform 1 0 77392 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_687
timestamp 1669390400
transform 1 0 78288 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_2
timestamp 1669390400
transform 1 0 1568 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_17
timestamp 1669390400
transform 1 0 3248 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_91_21
timestamp 1669390400
transform 1 0 3696 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_53
timestamp 1669390400
transform 1 0 7280 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_69
timestamp 1669390400
transform 1 0 9072 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_73
timestamp 1669390400
transform 1 0 9520 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_137
timestamp 1669390400
transform 1 0 16688 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_141
timestamp 1669390400
transform 1 0 17136 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_144
timestamp 1669390400
transform 1 0 17472 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_208
timestamp 1669390400
transform 1 0 24640 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_212
timestamp 1669390400
transform 1 0 25088 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_215
timestamp 1669390400
transform 1 0 25424 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_279
timestamp 1669390400
transform 1 0 32592 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_283
timestamp 1669390400
transform 1 0 33040 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_286
timestamp 1669390400
transform 1 0 33376 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_350
timestamp 1669390400
transform 1 0 40544 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_354
timestamp 1669390400
transform 1 0 40992 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_357
timestamp 1669390400
transform 1 0 41328 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_421
timestamp 1669390400
transform 1 0 48496 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_425
timestamp 1669390400
transform 1 0 48944 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_428
timestamp 1669390400
transform 1 0 49280 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_492
timestamp 1669390400
transform 1 0 56448 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_496
timestamp 1669390400
transform 1 0 56896 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_499
timestamp 1669390400
transform 1 0 57232 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_563
timestamp 1669390400
transform 1 0 64400 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_567
timestamp 1669390400
transform 1 0 64848 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_570
timestamp 1669390400
transform 1 0 65184 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_634
timestamp 1669390400
transform 1 0 72352 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_638
timestamp 1669390400
transform 1 0 72800 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_91_641
timestamp 1669390400
transform 1 0 73136 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_649
timestamp 1669390400
transform 1 0 74032 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_653
timestamp 1669390400
transform 1 0 74480 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_655
timestamp 1669390400
transform 1 0 74704 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_670
timestamp 1669390400
transform 1 0 76384 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_686
timestamp 1669390400
transform 1 0 78176 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_2
timestamp 1669390400
transform 1 0 1568 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_17
timestamp 1669390400
transform 1 0 3248 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_21
timestamp 1669390400
transform 1 0 3696 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_29
timestamp 1669390400
transform 1 0 4592 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_33
timestamp 1669390400
transform 1 0 5040 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_37
timestamp 1669390400
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_101
timestamp 1669390400
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_105
timestamp 1669390400
transform 1 0 13104 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_108
timestamp 1669390400
transform 1 0 13440 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_172
timestamp 1669390400
transform 1 0 20608 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_176
timestamp 1669390400
transform 1 0 21056 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_179
timestamp 1669390400
transform 1 0 21392 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_243
timestamp 1669390400
transform 1 0 28560 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_247
timestamp 1669390400
transform 1 0 29008 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_250
timestamp 1669390400
transform 1 0 29344 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_314
timestamp 1669390400
transform 1 0 36512 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_318
timestamp 1669390400
transform 1 0 36960 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_321
timestamp 1669390400
transform 1 0 37296 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_385
timestamp 1669390400
transform 1 0 44464 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_389
timestamp 1669390400
transform 1 0 44912 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_392
timestamp 1669390400
transform 1 0 45248 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_456
timestamp 1669390400
transform 1 0 52416 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_460
timestamp 1669390400
transform 1 0 52864 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_463
timestamp 1669390400
transform 1 0 53200 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_527
timestamp 1669390400
transform 1 0 60368 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_531
timestamp 1669390400
transform 1 0 60816 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_534
timestamp 1669390400
transform 1 0 61152 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_598
timestamp 1669390400
transform 1 0 68320 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_602
timestamp 1669390400
transform 1 0 68768 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_92_605
timestamp 1669390400
transform 1 0 69104 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_92_637
timestamp 1669390400
transform 1 0 72688 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_653
timestamp 1669390400
transform 1 0 74480 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_655
timestamp 1669390400
transform 1 0 74704 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_670
timestamp 1669390400
transform 1 0 76384 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_676
timestamp 1669390400
transform 1 0 77056 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_684
timestamp 1669390400
transform 1 0 77952 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_2
timestamp 1669390400
transform 1 0 1568 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_34
timestamp 1669390400
transform 1 0 5152 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_37
timestamp 1669390400
transform 1 0 5488 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_69
timestamp 1669390400
transform 1 0 9072 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_72
timestamp 1669390400
transform 1 0 9408 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_104
timestamp 1669390400
transform 1 0 12992 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_107
timestamp 1669390400
transform 1 0 13328 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_139
timestamp 1669390400
transform 1 0 16912 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_142
timestamp 1669390400
transform 1 0 17248 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_174
timestamp 1669390400
transform 1 0 20832 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_177
timestamp 1669390400
transform 1 0 21168 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_209
timestamp 1669390400
transform 1 0 24752 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_212
timestamp 1669390400
transform 1 0 25088 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_244
timestamp 1669390400
transform 1 0 28672 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_247
timestamp 1669390400
transform 1 0 29008 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_279
timestamp 1669390400
transform 1 0 32592 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_282
timestamp 1669390400
transform 1 0 32928 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_314
timestamp 1669390400
transform 1 0 36512 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_317
timestamp 1669390400
transform 1 0 36848 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_349
timestamp 1669390400
transform 1 0 40432 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_352
timestamp 1669390400
transform 1 0 40768 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_384
timestamp 1669390400
transform 1 0 44352 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_387
timestamp 1669390400
transform 1 0 44688 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_419
timestamp 1669390400
transform 1 0 48272 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_422
timestamp 1669390400
transform 1 0 48608 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_454
timestamp 1669390400
transform 1 0 52192 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_457
timestamp 1669390400
transform 1 0 52528 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_489
timestamp 1669390400
transform 1 0 56112 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_492
timestamp 1669390400
transform 1 0 56448 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_524
timestamp 1669390400
transform 1 0 60032 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_527
timestamp 1669390400
transform 1 0 60368 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_559
timestamp 1669390400
transform 1 0 63952 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_562
timestamp 1669390400
transform 1 0 64288 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_594
timestamp 1669390400
transform 1 0 67872 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_597
timestamp 1669390400
transform 1 0 68208 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_629
timestamp 1669390400
transform 1 0 71792 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_632
timestamp 1669390400
transform 1 0 72128 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_664
timestamp 1669390400
transform 1 0 75712 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_93_667
timestamp 1669390400
transform 1 0 76048 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_683
timestamp 1669390400
transform 1 0 77840 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_687
timestamp 1669390400
transform 1 0 78288 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 78624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 78624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 78624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 78624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 78624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 78624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 78624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 78624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 78624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 78624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 78624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 78624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 78624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 78624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 78624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 78624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 78624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 78624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 78624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 78624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 78624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 78624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 78624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 78624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 78624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_136
timestamp 1669390400
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_137
timestamp 1669390400
transform -1 0 78624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_138
timestamp 1669390400
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_139
timestamp 1669390400
transform -1 0 78624 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_140
timestamp 1669390400
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_141
timestamp 1669390400
transform -1 0 78624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_142
timestamp 1669390400
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_143
timestamp 1669390400
transform -1 0 78624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_144
timestamp 1669390400
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_145
timestamp 1669390400
transform -1 0 78624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_146
timestamp 1669390400
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_147
timestamp 1669390400
transform -1 0 78624 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_148
timestamp 1669390400
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_149
timestamp 1669390400
transform -1 0 78624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_150
timestamp 1669390400
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_151
timestamp 1669390400
transform -1 0 78624 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_152
timestamp 1669390400
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_153
timestamp 1669390400
transform -1 0 78624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_154
timestamp 1669390400
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_155
timestamp 1669390400
transform -1 0 78624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_156
timestamp 1669390400
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_157
timestamp 1669390400
transform -1 0 78624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_158
timestamp 1669390400
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_159
timestamp 1669390400
transform -1 0 78624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_160
timestamp 1669390400
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_161
timestamp 1669390400
transform -1 0 78624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_162
timestamp 1669390400
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_163
timestamp 1669390400
transform -1 0 78624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_164
timestamp 1669390400
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_165
timestamp 1669390400
transform -1 0 78624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_166
timestamp 1669390400
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_167
timestamp 1669390400
transform -1 0 78624 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_168
timestamp 1669390400
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_169
timestamp 1669390400
transform -1 0 78624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_170
timestamp 1669390400
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_171
timestamp 1669390400
transform -1 0 78624 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_172
timestamp 1669390400
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_173
timestamp 1669390400
transform -1 0 78624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_174
timestamp 1669390400
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_175
timestamp 1669390400
transform -1 0 78624 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_176
timestamp 1669390400
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_177
timestamp 1669390400
transform -1 0 78624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_178
timestamp 1669390400
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_179
timestamp 1669390400
transform -1 0 78624 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_180
timestamp 1669390400
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_181
timestamp 1669390400
transform -1 0 78624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_182
timestamp 1669390400
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_183
timestamp 1669390400
transform -1 0 78624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_184
timestamp 1669390400
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_185
timestamp 1669390400
transform -1 0 78624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_186
timestamp 1669390400
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_187
timestamp 1669390400
transform -1 0 78624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 60928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 68880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 76832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 64960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 72912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 60928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 68880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 76832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1669390400
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1669390400
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1669390400
transform 1 0 64960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1669390400
transform 1 0 72912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1669390400
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1669390400
transform 1 0 60928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1669390400
transform 1 0 68880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1669390400
transform 1 0 76832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1669390400
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1669390400
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1669390400
transform 1 0 64960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1669390400
transform 1 0 72912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1669390400
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1669390400
transform 1 0 60928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1669390400
transform 1 0 68880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1669390400
transform 1 0 76832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1669390400
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1669390400
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1669390400
transform 1 0 64960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1669390400
transform 1 0 72912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1669390400
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1669390400
transform 1 0 60928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1669390400
transform 1 0 68880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1669390400
transform 1 0 76832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1669390400
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1669390400
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1669390400
transform 1 0 64960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1669390400
transform 1 0 72912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1669390400
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1669390400
transform 1 0 60928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1669390400
transform 1 0 68880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1669390400
transform 1 0 76832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1669390400
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1669390400
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1669390400
transform 1 0 64960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1669390400
transform 1 0 72912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1669390400
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1669390400
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1669390400
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1669390400
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1669390400
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1669390400
transform 1 0 60928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1669390400
transform 1 0 68880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1669390400
transform 1 0 76832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1669390400
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1669390400
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1669390400
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1669390400
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1669390400
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1669390400
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1669390400
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1669390400
transform 1 0 64960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1669390400
transform 1 0 72912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1669390400
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1669390400
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1669390400
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1669390400
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1669390400
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1669390400
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1669390400
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1669390400
transform 1 0 60928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1669390400
transform 1 0 68880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1669390400
transform 1 0 76832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1669390400
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1669390400
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1669390400
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1669390400
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1669390400
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1669390400
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1669390400
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1669390400
transform 1 0 64960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1669390400
transform 1 0 72912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1669390400
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1669390400
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1669390400
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1669390400
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1669390400
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1669390400
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1669390400
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1669390400
transform 1 0 60928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1669390400
transform 1 0 68880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1669390400
transform 1 0 76832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1669390400
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1669390400
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1669390400
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1669390400
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1669390400
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1669390400
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1669390400
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1669390400
transform 1 0 64960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1669390400
transform 1 0 72912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1669390400
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1669390400
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1669390400
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1669390400
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1669390400
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1669390400
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1669390400
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1669390400
transform 1 0 60928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1669390400
transform 1 0 68880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1669390400
transform 1 0 76832 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1669390400
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1669390400
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1669390400
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1669390400
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1669390400
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1669390400
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1669390400
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1669390400
transform 1 0 64960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1669390400
transform 1 0 72912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1669390400
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1669390400
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1669390400
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1669390400
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1669390400
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1669390400
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1669390400
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1669390400
transform 1 0 60928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1669390400
transform 1 0 68880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1669390400
transform 1 0 76832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1669390400
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1669390400
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1669390400
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1669390400
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1669390400
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1669390400
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1669390400
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1669390400
transform 1 0 64960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1669390400
transform 1 0 72912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1669390400
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1669390400
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1669390400
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1669390400
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1669390400
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1669390400
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1669390400
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1669390400
transform 1 0 60928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1669390400
transform 1 0 68880 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1669390400
transform 1 0 76832 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1669390400
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1669390400
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1669390400
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1669390400
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1669390400
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1669390400
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1669390400
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1669390400
transform 1 0 64960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1669390400
transform 1 0 72912 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1669390400
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1669390400
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1669390400
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1669390400
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1669390400
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1669390400
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1669390400
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1669390400
transform 1 0 60928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1669390400
transform 1 0 68880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1669390400
transform 1 0 76832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1669390400
transform 1 0 9296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1669390400
transform 1 0 17248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1669390400
transform 1 0 25200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1669390400
transform 1 0 33152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1669390400
transform 1 0 41104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1669390400
transform 1 0 49056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1669390400
transform 1 0 57008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1669390400
transform 1 0 64960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1669390400
transform 1 0 72912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1669390400
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1669390400
transform 1 0 13216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1669390400
transform 1 0 21168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1669390400
transform 1 0 29120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1669390400
transform 1 0 37072 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1669390400
transform 1 0 45024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1669390400
transform 1 0 52976 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1669390400
transform 1 0 60928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1669390400
transform 1 0 68880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1669390400
transform 1 0 76832 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1669390400
transform 1 0 9296 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1669390400
transform 1 0 17248 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1669390400
transform 1 0 25200 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1669390400
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1669390400
transform 1 0 41104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1669390400
transform 1 0 49056 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1669390400
transform 1 0 57008 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1669390400
transform 1 0 64960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1669390400
transform 1 0 72912 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1669390400
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1669390400
transform 1 0 13216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1669390400
transform 1 0 21168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1669390400
transform 1 0 29120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1669390400
transform 1 0 37072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1669390400
transform 1 0 45024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1669390400
transform 1 0 52976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1669390400
transform 1 0 60928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1669390400
transform 1 0 68880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1669390400
transform 1 0 76832 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1669390400
transform 1 0 9296 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1669390400
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1669390400
transform 1 0 25200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1669390400
transform 1 0 33152 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1669390400
transform 1 0 41104 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1669390400
transform 1 0 49056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1669390400
transform 1 0 57008 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1669390400
transform 1 0 64960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1669390400
transform 1 0 72912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1669390400
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1669390400
transform 1 0 13216 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1669390400
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1669390400
transform 1 0 29120 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1669390400
transform 1 0 37072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1669390400
transform 1 0 45024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1669390400
transform 1 0 52976 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1669390400
transform 1 0 60928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1669390400
transform 1 0 68880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1669390400
transform 1 0 76832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1669390400
transform 1 0 9296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1669390400
transform 1 0 17248 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1669390400
transform 1 0 25200 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1669390400
transform 1 0 33152 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1669390400
transform 1 0 41104 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1669390400
transform 1 0 49056 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1669390400
transform 1 0 57008 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_898
timestamp 1669390400
transform 1 0 64960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_899
timestamp 1669390400
transform 1 0 72912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_900
timestamp 1669390400
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_901
timestamp 1669390400
transform 1 0 13216 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_902
timestamp 1669390400
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_903
timestamp 1669390400
transform 1 0 29120 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_904
timestamp 1669390400
transform 1 0 37072 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_905
timestamp 1669390400
transform 1 0 45024 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_906
timestamp 1669390400
transform 1 0 52976 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_907
timestamp 1669390400
transform 1 0 60928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_908
timestamp 1669390400
transform 1 0 68880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_909
timestamp 1669390400
transform 1 0 76832 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_910
timestamp 1669390400
transform 1 0 9296 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_911
timestamp 1669390400
transform 1 0 17248 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_912
timestamp 1669390400
transform 1 0 25200 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_913
timestamp 1669390400
transform 1 0 33152 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_914
timestamp 1669390400
transform 1 0 41104 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_915
timestamp 1669390400
transform 1 0 49056 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_916
timestamp 1669390400
transform 1 0 57008 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_917
timestamp 1669390400
transform 1 0 64960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_918
timestamp 1669390400
transform 1 0 72912 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_919
timestamp 1669390400
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_920
timestamp 1669390400
transform 1 0 13216 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_921
timestamp 1669390400
transform 1 0 21168 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_922
timestamp 1669390400
transform 1 0 29120 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_923
timestamp 1669390400
transform 1 0 37072 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_924
timestamp 1669390400
transform 1 0 45024 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_925
timestamp 1669390400
transform 1 0 52976 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_926
timestamp 1669390400
transform 1 0 60928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_927
timestamp 1669390400
transform 1 0 68880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_928
timestamp 1669390400
transform 1 0 76832 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_929
timestamp 1669390400
transform 1 0 9296 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_930
timestamp 1669390400
transform 1 0 17248 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_931
timestamp 1669390400
transform 1 0 25200 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_932
timestamp 1669390400
transform 1 0 33152 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_933
timestamp 1669390400
transform 1 0 41104 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_934
timestamp 1669390400
transform 1 0 49056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_935
timestamp 1669390400
transform 1 0 57008 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_936
timestamp 1669390400
transform 1 0 64960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_937
timestamp 1669390400
transform 1 0 72912 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_938
timestamp 1669390400
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_939
timestamp 1669390400
transform 1 0 13216 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_940
timestamp 1669390400
transform 1 0 21168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_941
timestamp 1669390400
transform 1 0 29120 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_942
timestamp 1669390400
transform 1 0 37072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_943
timestamp 1669390400
transform 1 0 45024 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_944
timestamp 1669390400
transform 1 0 52976 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_945
timestamp 1669390400
transform 1 0 60928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_946
timestamp 1669390400
transform 1 0 68880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_947
timestamp 1669390400
transform 1 0 76832 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_948
timestamp 1669390400
transform 1 0 9296 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_949
timestamp 1669390400
transform 1 0 17248 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_950
timestamp 1669390400
transform 1 0 25200 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_951
timestamp 1669390400
transform 1 0 33152 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_952
timestamp 1669390400
transform 1 0 41104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_953
timestamp 1669390400
transform 1 0 49056 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_954
timestamp 1669390400
transform 1 0 57008 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_955
timestamp 1669390400
transform 1 0 64960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_956
timestamp 1669390400
transform 1 0 72912 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_957
timestamp 1669390400
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_958
timestamp 1669390400
transform 1 0 13216 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_959
timestamp 1669390400
transform 1 0 21168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_960
timestamp 1669390400
transform 1 0 29120 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_961
timestamp 1669390400
transform 1 0 37072 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_962
timestamp 1669390400
transform 1 0 45024 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_963
timestamp 1669390400
transform 1 0 52976 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_964
timestamp 1669390400
transform 1 0 60928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_965
timestamp 1669390400
transform 1 0 68880 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_966
timestamp 1669390400
transform 1 0 76832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_967
timestamp 1669390400
transform 1 0 9296 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_968
timestamp 1669390400
transform 1 0 17248 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_969
timestamp 1669390400
transform 1 0 25200 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_970
timestamp 1669390400
transform 1 0 33152 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_971
timestamp 1669390400
transform 1 0 41104 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_972
timestamp 1669390400
transform 1 0 49056 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_973
timestamp 1669390400
transform 1 0 57008 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_974
timestamp 1669390400
transform 1 0 64960 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_975
timestamp 1669390400
transform 1 0 72912 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_976
timestamp 1669390400
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_977
timestamp 1669390400
transform 1 0 13216 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_978
timestamp 1669390400
transform 1 0 21168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_979
timestamp 1669390400
transform 1 0 29120 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_980
timestamp 1669390400
transform 1 0 37072 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_981
timestamp 1669390400
transform 1 0 45024 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_982
timestamp 1669390400
transform 1 0 52976 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_983
timestamp 1669390400
transform 1 0 60928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_984
timestamp 1669390400
transform 1 0 68880 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_985
timestamp 1669390400
transform 1 0 76832 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_986
timestamp 1669390400
transform 1 0 9296 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_987
timestamp 1669390400
transform 1 0 17248 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_988
timestamp 1669390400
transform 1 0 25200 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_989
timestamp 1669390400
transform 1 0 33152 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_990
timestamp 1669390400
transform 1 0 41104 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_991
timestamp 1669390400
transform 1 0 49056 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_992
timestamp 1669390400
transform 1 0 57008 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_993
timestamp 1669390400
transform 1 0 64960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_994
timestamp 1669390400
transform 1 0 72912 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_995
timestamp 1669390400
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_996
timestamp 1669390400
transform 1 0 13216 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_997
timestamp 1669390400
transform 1 0 21168 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_998
timestamp 1669390400
transform 1 0 29120 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_999
timestamp 1669390400
transform 1 0 37072 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1000
timestamp 1669390400
transform 1 0 45024 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1001
timestamp 1669390400
transform 1 0 52976 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1002
timestamp 1669390400
transform 1 0 60928 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1003
timestamp 1669390400
transform 1 0 68880 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1004
timestamp 1669390400
transform 1 0 76832 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1005
timestamp 1669390400
transform 1 0 9296 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1006
timestamp 1669390400
transform 1 0 17248 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1007
timestamp 1669390400
transform 1 0 25200 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1008
timestamp 1669390400
transform 1 0 33152 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1009
timestamp 1669390400
transform 1 0 41104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1010
timestamp 1669390400
transform 1 0 49056 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1011
timestamp 1669390400
transform 1 0 57008 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1012
timestamp 1669390400
transform 1 0 64960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1013
timestamp 1669390400
transform 1 0 72912 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1014
timestamp 1669390400
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1015
timestamp 1669390400
transform 1 0 13216 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1016
timestamp 1669390400
transform 1 0 21168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1017
timestamp 1669390400
transform 1 0 29120 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1018
timestamp 1669390400
transform 1 0 37072 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1019
timestamp 1669390400
transform 1 0 45024 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1020
timestamp 1669390400
transform 1 0 52976 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1021
timestamp 1669390400
transform 1 0 60928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1022
timestamp 1669390400
transform 1 0 68880 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1023
timestamp 1669390400
transform 1 0 76832 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1024
timestamp 1669390400
transform 1 0 9296 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1025
timestamp 1669390400
transform 1 0 17248 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1026
timestamp 1669390400
transform 1 0 25200 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1027
timestamp 1669390400
transform 1 0 33152 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1028
timestamp 1669390400
transform 1 0 41104 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1029
timestamp 1669390400
transform 1 0 49056 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1030
timestamp 1669390400
transform 1 0 57008 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1031
timestamp 1669390400
transform 1 0 64960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1032
timestamp 1669390400
transform 1 0 72912 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1033
timestamp 1669390400
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1034
timestamp 1669390400
transform 1 0 13216 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1035
timestamp 1669390400
transform 1 0 21168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1036
timestamp 1669390400
transform 1 0 29120 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1037
timestamp 1669390400
transform 1 0 37072 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1038
timestamp 1669390400
transform 1 0 45024 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1039
timestamp 1669390400
transform 1 0 52976 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1040
timestamp 1669390400
transform 1 0 60928 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1041
timestamp 1669390400
transform 1 0 68880 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1042
timestamp 1669390400
transform 1 0 76832 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1043
timestamp 1669390400
transform 1 0 9296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1044
timestamp 1669390400
transform 1 0 17248 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1045
timestamp 1669390400
transform 1 0 25200 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1046
timestamp 1669390400
transform 1 0 33152 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1047
timestamp 1669390400
transform 1 0 41104 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1048
timestamp 1669390400
transform 1 0 49056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1049
timestamp 1669390400
transform 1 0 57008 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1050
timestamp 1669390400
transform 1 0 64960 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1051
timestamp 1669390400
transform 1 0 72912 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1052
timestamp 1669390400
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1053
timestamp 1669390400
transform 1 0 13216 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1054
timestamp 1669390400
transform 1 0 21168 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1055
timestamp 1669390400
transform 1 0 29120 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1056
timestamp 1669390400
transform 1 0 37072 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1057
timestamp 1669390400
transform 1 0 45024 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1058
timestamp 1669390400
transform 1 0 52976 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1059
timestamp 1669390400
transform 1 0 60928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1060
timestamp 1669390400
transform 1 0 68880 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1061
timestamp 1669390400
transform 1 0 76832 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1062
timestamp 1669390400
transform 1 0 9296 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1063
timestamp 1669390400
transform 1 0 17248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1064
timestamp 1669390400
transform 1 0 25200 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1065
timestamp 1669390400
transform 1 0 33152 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1066
timestamp 1669390400
transform 1 0 41104 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1067
timestamp 1669390400
transform 1 0 49056 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1068
timestamp 1669390400
transform 1 0 57008 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1069
timestamp 1669390400
transform 1 0 64960 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1070
timestamp 1669390400
transform 1 0 72912 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1071
timestamp 1669390400
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1072
timestamp 1669390400
transform 1 0 13216 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1073
timestamp 1669390400
transform 1 0 21168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1074
timestamp 1669390400
transform 1 0 29120 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1075
timestamp 1669390400
transform 1 0 37072 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1076
timestamp 1669390400
transform 1 0 45024 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1077
timestamp 1669390400
transform 1 0 52976 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1078
timestamp 1669390400
transform 1 0 60928 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1079
timestamp 1669390400
transform 1 0 68880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1080
timestamp 1669390400
transform 1 0 76832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1081
timestamp 1669390400
transform 1 0 5264 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1082
timestamp 1669390400
transform 1 0 9184 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1083
timestamp 1669390400
transform 1 0 13104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1084
timestamp 1669390400
transform 1 0 17024 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1085
timestamp 1669390400
transform 1 0 20944 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1086
timestamp 1669390400
transform 1 0 24864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1087
timestamp 1669390400
transform 1 0 28784 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1088
timestamp 1669390400
transform 1 0 32704 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1089
timestamp 1669390400
transform 1 0 36624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1090
timestamp 1669390400
transform 1 0 40544 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1091
timestamp 1669390400
transform 1 0 44464 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1092
timestamp 1669390400
transform 1 0 48384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1093
timestamp 1669390400
transform 1 0 52304 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1094
timestamp 1669390400
transform 1 0 56224 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1095
timestamp 1669390400
transform 1 0 60144 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1096
timestamp 1669390400
transform 1 0 64064 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1097
timestamp 1669390400
transform 1 0 67984 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1098
timestamp 1669390400
transform 1 0 71904 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1099
timestamp 1669390400
transform 1 0 75824 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _100_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 72464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _101_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 19936 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _102_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 25760 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _103_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 25536 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _104_
timestamp 1669390400
transform 1 0 17920 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _105_
timestamp 1669390400
transform -1 0 23856 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _106_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22512 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _107_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 54768 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _108_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 54768 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _109_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 56784 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _110_
timestamp 1669390400
transform 1 0 67200 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _111_
timestamp 1669390400
transform 1 0 69216 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _112_
timestamp 1669390400
transform 1 0 56000 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _113_
timestamp 1669390400
transform 1 0 55440 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _114_
timestamp 1669390400
transform 1 0 56672 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _115_
timestamp 1669390400
transform 1 0 66864 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _116_
timestamp 1669390400
transform 1 0 68096 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _117_
timestamp 1669390400
transform -1 0 73696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _118_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 73248 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _119_
timestamp 1669390400
transform 1 0 66976 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _120_
timestamp 1669390400
transform -1 0 69664 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _121_
timestamp 1669390400
transform -1 0 68768 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _122_
timestamp 1669390400
transform 1 0 48272 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _123_
timestamp 1669390400
transform 1 0 56112 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _124_
timestamp 1669390400
transform -1 0 53984 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _125_
timestamp 1669390400
transform 1 0 55888 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_
timestamp 1669390400
transform -1 0 51072 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _127_
timestamp 1669390400
transform -1 0 49840 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _128_
timestamp 1669390400
transform 1 0 49056 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _129_
timestamp 1669390400
transform 1 0 48048 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _130_
timestamp 1669390400
transform -1 0 50848 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _131_
timestamp 1669390400
transform -1 0 50512 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _132_
timestamp 1669390400
transform 1 0 46480 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _133_
timestamp 1669390400
transform -1 0 51744 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _134_
timestamp 1669390400
transform -1 0 51072 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _135_
timestamp 1669390400
transform 1 0 49280 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _136_
timestamp 1669390400
transform -1 0 51968 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _137_
timestamp 1669390400
transform -1 0 51296 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _138_
timestamp 1669390400
transform 1 0 49392 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _139_
timestamp 1669390400
transform -1 0 53872 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _140_
timestamp 1669390400
transform 1 0 51520 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _141_
timestamp 1669390400
transform -1 0 59584 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _142_
timestamp 1669390400
transform -1 0 52752 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _143_
timestamp 1669390400
transform 1 0 48160 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _144_
timestamp 1669390400
transform -1 0 60816 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _145_
timestamp 1669390400
transform -1 0 52864 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _146_
timestamp 1669390400
transform 1 0 48160 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _147_
timestamp 1669390400
transform -1 0 57792 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _148_
timestamp 1669390400
transform -1 0 54432 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _149_
timestamp 1669390400
transform 1 0 50288 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _150_
timestamp 1669390400
transform -1 0 53760 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _151_
timestamp 1669390400
transform -1 0 53760 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _152_
timestamp 1669390400
transform 1 0 52640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _153_
timestamp 1669390400
transform -1 0 56112 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _154_
timestamp 1669390400
transform 1 0 53984 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _155_
timestamp 1669390400
transform 1 0 53760 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _156_
timestamp 1669390400
transform 1 0 54096 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _157_
timestamp 1669390400
transform 1 0 51968 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _158_
timestamp 1669390400
transform -1 0 56224 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _159_
timestamp 1669390400
transform -1 0 55552 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _160_
timestamp 1669390400
transform 1 0 50512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _161_
timestamp 1669390400
transform -1 0 56896 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _162_
timestamp 1669390400
transform -1 0 56112 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _163_
timestamp 1669390400
transform 1 0 52976 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _164_
timestamp 1669390400
transform -1 0 56896 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _165_
timestamp 1669390400
transform -1 0 56224 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _166_
timestamp 1669390400
transform 1 0 56448 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _167_
timestamp 1669390400
transform 1 0 56896 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _168_
timestamp 1669390400
transform 1 0 56784 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _169_
timestamp 1669390400
transform -1 0 59136 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _170_
timestamp 1669390400
transform -1 0 58464 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _171_
timestamp 1669390400
transform 1 0 54992 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _172_
timestamp 1669390400
transform -1 0 63056 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _173_
timestamp 1669390400
transform -1 0 58240 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _174_
timestamp 1669390400
transform 1 0 55888 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _175_
timestamp 1669390400
transform -1 0 59472 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _176_
timestamp 1669390400
transform -1 0 58688 0 -1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _177_
timestamp 1669390400
transform 1 0 57008 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _178_
timestamp 1669390400
transform 1 0 58240 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _179_
timestamp 1669390400
transform -1 0 58800 0 1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _180_
timestamp 1669390400
transform 1 0 58688 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _181_
timestamp 1669390400
transform -1 0 61600 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _182_
timestamp 1669390400
transform 1 0 59248 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _183_
timestamp 1669390400
transform -1 0 61712 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _184_
timestamp 1669390400
transform -1 0 60480 0 -1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _185_
timestamp 1669390400
transform 1 0 57904 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _186_
timestamp 1669390400
transform -1 0 66752 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _187_
timestamp 1669390400
transform -1 0 60816 0 1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _188_
timestamp 1669390400
transform 1 0 57344 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _189_
timestamp 1669390400
transform -1 0 64736 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _190_
timestamp 1669390400
transform -1 0 61600 0 -1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _191_
timestamp 1669390400
transform 1 0 60144 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _192_
timestamp 1669390400
transform 1 0 61376 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _193_
timestamp 1669390400
transform 1 0 61824 0 -1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _194_
timestamp 1669390400
transform 1 0 61264 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _195_
timestamp 1669390400
transform -1 0 63840 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _196_
timestamp 1669390400
transform 1 0 62048 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _197_
timestamp 1669390400
transform 1 0 61488 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _198_
timestamp 1669390400
transform 1 0 62160 0 -1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _199_
timestamp 1669390400
transform 1 0 59472 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _200_
timestamp 1669390400
transform -1 0 68432 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _201_
timestamp 1669390400
transform -1 0 64624 0 -1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _202_
timestamp 1669390400
transform 1 0 59136 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _203_
timestamp 1669390400
transform -1 0 64512 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _204_
timestamp 1669390400
transform -1 0 64064 0 1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _205_
timestamp 1669390400
transform 1 0 60928 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _206_
timestamp 1669390400
transform -1 0 64848 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _207_
timestamp 1669390400
transform -1 0 64176 0 -1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _208_
timestamp 1669390400
transform 1 0 61600 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _209_
timestamp 1669390400
transform -1 0 66864 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _210_
timestamp 1669390400
transform 1 0 65296 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _211_
timestamp 1669390400
transform -1 0 66640 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _212_
timestamp 1669390400
transform -1 0 65968 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _213_
timestamp 1669390400
transform 1 0 61824 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _214_
timestamp 1669390400
transform 1 0 64400 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _215_
timestamp 1669390400
transform 1 0 65296 0 -1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _216_
timestamp 1669390400
transform 1 0 63168 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _217_
timestamp 1669390400
transform -1 0 67088 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _218_
timestamp 1669390400
transform -1 0 66416 0 1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _219_
timestamp 1669390400
transform 1 0 63280 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _220_
timestamp 1669390400
transform -1 0 67200 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _221_
timestamp 1669390400
transform -1 0 66528 0 -1 67424
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _222_
timestamp 1669390400
transform 1 0 67088 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _223_
timestamp 1669390400
transform -1 0 69664 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _224_
timestamp 1669390400
transform -1 0 68544 0 1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _225_
timestamp 1669390400
transform 1 0 67760 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _226_
timestamp 1669390400
transform -1 0 69664 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _227_
timestamp 1669390400
transform -1 0 68880 0 -1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _228_
timestamp 1669390400
transform 1 0 67536 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _229_
timestamp 1669390400
transform 1 0 68432 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _230_
timestamp 1669390400
transform -1 0 68992 0 -1 67424
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _231_
timestamp 1669390400
transform -1 0 73696 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _232_
timestamp 1669390400
transform -1 0 74368 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _233_
timestamp 1669390400
transform -1 0 74368 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _234_
timestamp 1669390400
transform 1 0 73472 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _235_
timestamp 1669390400
transform 1 0 69216 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _236_
timestamp 1669390400
transform 1 0 68656 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _237_
timestamp 1669390400
transform 1 0 4480 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _238_
timestamp 1669390400
transform 1 0 6272 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _239_
timestamp 1669390400
transform 1 0 6832 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _240_
timestamp 1669390400
transform 1 0 7728 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _241_
timestamp 1669390400
transform 1 0 8288 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _242_
timestamp 1669390400
transform 1 0 8960 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _243_
timestamp 1669390400
transform 1 0 9744 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _244_
timestamp 1669390400
transform 1 0 10416 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _245_
timestamp 1669390400
transform 1 0 10976 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _246_
timestamp 1669390400
transform 1 0 11424 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _247_
timestamp 1669390400
transform 1 0 12320 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _248_
timestamp 1669390400
transform 1 0 12992 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _249_
timestamp 1669390400
transform 1 0 57344 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _250_
timestamp 1669390400
transform 1 0 55216 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _251_
timestamp 1669390400
transform 1 0 55888 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _252_
timestamp 1669390400
transform 1 0 55888 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _253_
timestamp 1669390400
transform 1 0 19264 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _254_
timestamp 1669390400
transform 1 0 19040 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _255_
timestamp 1669390400
transform 1 0 18032 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _256_
timestamp 1669390400
transform 1 0 18368 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _257_
timestamp 1669390400
transform 1 0 20608 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _258_
timestamp 1669390400
transform 1 0 21504 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _259_
timestamp 1669390400
transform 1 0 20384 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _260_
timestamp 1669390400
transform 1 0 20720 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _261_
timestamp 1669390400
transform 1 0 23072 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _262_
timestamp 1669390400
transform 1 0 23520 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _263_
timestamp 1669390400
transform 1 0 22848 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _264_
timestamp 1669390400
transform 1 0 23408 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _265_
timestamp 1669390400
transform 1 0 25200 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _266_
timestamp 1669390400
transform 1 0 24416 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _267_
timestamp 1669390400
transform 1 0 25648 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _268_
timestamp 1669390400
transform 1 0 26208 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _269_
timestamp 1669390400
transform -1 0 5152 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _270_
timestamp 1669390400
transform -1 0 5152 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _271_
timestamp 1669390400
transform -1 0 6608 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _272_
timestamp 1669390400
transform -1 0 7056 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _273_
timestamp 1669390400
transform -1 0 7952 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _274_
timestamp 1669390400
transform -1 0 8624 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _275_
timestamp 1669390400
transform -1 0 9184 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _276_
timestamp 1669390400
transform -1 0 9968 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _277_
timestamp 1669390400
transform -1 0 10640 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _278_
timestamp 1669390400
transform -1 0 11200 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _279_
timestamp 1669390400
transform -1 0 11872 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _280_
timestamp 1669390400
transform -1 0 12768 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _281_
timestamp 1669390400
transform -1 0 12992 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _282_
timestamp 1669390400
transform -1 0 13888 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _283_
timestamp 1669390400
transform -1 0 14560 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _284_
timestamp 1669390400
transform -1 0 15232 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _285_
timestamp 1669390400
transform -1 0 16352 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _286_
timestamp 1669390400
transform -1 0 16240 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _287_
timestamp 1669390400
transform -1 0 17136 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _288_
timestamp 1669390400
transform -1 0 18144 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _289_
timestamp 1669390400
transform -1 0 19152 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _290_
timestamp 1669390400
transform -1 0 19264 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _291_
timestamp 1669390400
transform -1 0 20160 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _292_
timestamp 1669390400
transform -1 0 20496 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _293_
timestamp 1669390400
transform -1 0 22176 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _294_
timestamp 1669390400
transform -1 0 22288 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _295_
timestamp 1669390400
transform -1 0 22624 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _296_
timestamp 1669390400
transform -1 0 22960 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _297_
timestamp 1669390400
transform -1 0 24192 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _298_
timestamp 1669390400
transform -1 0 24192 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _299_
timestamp 1669390400
transform -1 0 24864 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _300_
timestamp 1669390400
transform -1 0 25760 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _301_
timestamp 1669390400
transform 1 0 27216 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _302_
timestamp 1669390400
transform 1 0 27776 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _303_
timestamp 1669390400
transform 1 0 28448 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _304_
timestamp 1669390400
transform 1 0 29456 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _305_
timestamp 1669390400
transform 1 0 29904 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _306_
timestamp 1669390400
transform 1 0 30352 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _307_
timestamp 1669390400
transform 1 0 31248 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _308_
timestamp 1669390400
transform 1 0 31808 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _309_
timestamp 1669390400
transform 1 0 32592 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _310_
timestamp 1669390400
transform 1 0 33488 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _311_
timestamp 1669390400
transform 1 0 33936 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _312_
timestamp 1669390400
transform 1 0 34608 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _313_
timestamp 1669390400
transform 1 0 35056 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _314_
timestamp 1669390400
transform 1 0 35952 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _315_
timestamp 1669390400
transform 1 0 36512 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _316_
timestamp 1669390400
transform 1 0 37408 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _317_
timestamp 1669390400
transform 1 0 37968 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _318_
timestamp 1669390400
transform 1 0 38640 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _319_
timestamp 1669390400
transform 1 0 39200 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _320_
timestamp 1669390400
transform 1 0 39648 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _321_
timestamp 1669390400
transform 1 0 40544 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _322_
timestamp 1669390400
transform 1 0 41440 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _323_
timestamp 1669390400
transform 1 0 42000 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _324_
timestamp 1669390400
transform 1 0 42672 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _325_
timestamp 1669390400
transform 1 0 43232 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _326_
timestamp 1669390400
transform 1 0 44016 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _327_
timestamp 1669390400
transform 1 0 45360 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _328_
timestamp 1669390400
transform 1 0 45136 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _329_
timestamp 1669390400
transform 1 0 46928 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _330_
timestamp 1669390400
transform 1 0 46704 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _331_
timestamp 1669390400
transform 1 0 47264 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _332_
timestamp 1669390400
transform 1 0 47936 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _333_
timestamp 1669390400
transform -1 0 26768 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _334_
timestamp 1669390400
transform -1 0 27440 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _335_
timestamp 1669390400
transform -1 0 28112 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _336_
timestamp 1669390400
transform -1 0 28784 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _337_
timestamp 1669390400
transform -1 0 29456 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _338_
timestamp 1669390400
transform -1 0 30128 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _339_
timestamp 1669390400
transform -1 0 30576 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _340_
timestamp 1669390400
transform -1 0 31472 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _341_
timestamp 1669390400
transform -1 0 32144 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _342_
timestamp 1669390400
transform -1 0 32816 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _343_
timestamp 1669390400
transform -1 0 33488 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _344_
timestamp 1669390400
transform -1 0 34272 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _345_
timestamp 1669390400
transform -1 0 34832 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _346_
timestamp 1669390400
transform -1 0 35280 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _347_
timestamp 1669390400
transform -1 0 36176 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _348_
timestamp 1669390400
transform -1 0 36848 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _349_
timestamp 1669390400
transform -1 0 37520 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _350_
timestamp 1669390400
transform -1 0 38192 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _351_
timestamp 1669390400
transform -1 0 38864 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _352_
timestamp 1669390400
transform -1 0 39424 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _353_
timestamp 1669390400
transform -1 0 39984 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _354_
timestamp 1669390400
transform -1 0 40880 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _355_
timestamp 1669390400
transform -1 0 41552 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _356_
timestamp 1669390400
transform -1 0 42336 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _357_
timestamp 1669390400
transform -1 0 42896 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _358_
timestamp 1669390400
transform -1 0 43568 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _359_
timestamp 1669390400
transform -1 0 44240 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _360_
timestamp 1669390400
transform -1 0 44912 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _361_
timestamp 1669390400
transform -1 0 46704 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _362_
timestamp 1669390400
transform -1 0 46256 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _363_
timestamp 1669390400
transform -1 0 46928 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _364_
timestamp 1669390400
transform -1 0 47600 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _365_
timestamp 1669390400
transform 1 0 70784 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _366_
timestamp 1669390400
transform 1 0 71456 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _367_
timestamp 1669390400
transform 1 0 72016 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _368_
timestamp 1669390400
transform 1 0 72800 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _369_
timestamp 1669390400
transform -1 0 70448 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _370_
timestamp 1669390400
transform -1 0 71120 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _371_
timestamp 1669390400
transform -1 0 71792 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _372_
timestamp 1669390400
transform -1 0 72352 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _373_
timestamp 1669390400
transform 1 0 70112 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _374_
timestamp 1669390400
transform -1 0 69888 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 76608 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform 1 0 1680 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform -1 0 7168 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input4
timestamp 1669390400
transform 1 0 11200 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input5
timestamp 1669390400
transform 1 0 12096 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1669390400
transform 1 0 13552 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input7 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 14112 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input8
timestamp 1669390400
transform 1 0 14112 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input9
timestamp 1669390400
transform 1 0 17360 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input10
timestamp 1669390400
transform 1 0 15344 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input11
timestamp 1669390400
transform -1 0 17920 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input12
timestamp 1669390400
transform 1 0 15232 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input13
timestamp 1669390400
transform 1 0 18144 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input14
timestamp 1669390400
transform 1 0 3360 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input15
timestamp 1669390400
transform 1 0 17248 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input16
timestamp 1669390400
transform -1 0 20608 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input17
timestamp 1669390400
transform 1 0 19264 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input18
timestamp 1669390400
transform -1 0 22624 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input19
timestamp 1669390400
transform 1 0 19264 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input20
timestamp 1669390400
transform 1 0 22176 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input21
timestamp 1669390400
transform 1 0 22848 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input22
timestamp 1669390400
transform 1 0 21280 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input23
timestamp 1669390400
transform 1 0 23184 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input24
timestamp 1669390400
transform -1 0 25088 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input25
timestamp 1669390400
transform -1 0 7168 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input26
timestamp 1669390400
transform 1 0 22960 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input27
timestamp 1669390400
transform -1 0 26992 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input28
timestamp 1669390400
transform -1 0 9184 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input29
timestamp 1669390400
transform -1 0 9072 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input30
timestamp 1669390400
transform 1 0 7392 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input31
timestamp 1669390400
transform 1 0 7280 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input32
timestamp 1669390400
transform -1 0 11088 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input33
timestamp 1669390400
transform -1 0 11872 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input34
timestamp 1669390400
transform -1 0 13104 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input35
timestamp 1669390400
transform -1 0 77056 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input36
timestamp 1669390400
transform -1 0 76608 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input37
timestamp 1669390400
transform -1 0 76608 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input38
timestamp 1669390400
transform -1 0 76608 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input39
timestamp 1669390400
transform -1 0 76608 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input40
timestamp 1669390400
transform -1 0 76608 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input41
timestamp 1669390400
transform -1 0 76608 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input42
timestamp 1669390400
transform -1 0 76608 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input43
timestamp 1669390400
transform -1 0 76608 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input44
timestamp 1669390400
transform -1 0 74592 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input45
timestamp 1669390400
transform -1 0 76608 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input46
timestamp 1669390400
transform -1 0 76608 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input47
timestamp 1669390400
transform -1 0 76608 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input48
timestamp 1669390400
transform -1 0 76608 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input49
timestamp 1669390400
transform -1 0 76608 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input50
timestamp 1669390400
transform -1 0 76608 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input51
timestamp 1669390400
transform -1 0 76608 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input52
timestamp 1669390400
transform -1 0 74592 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input53
timestamp 1669390400
transform -1 0 76608 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input54
timestamp 1669390400
transform -1 0 76608 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input55
timestamp 1669390400
transform -1 0 76608 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input56
timestamp 1669390400
transform -1 0 76608 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input57
timestamp 1669390400
transform -1 0 76608 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input58
timestamp 1669390400
transform -1 0 76608 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input59
timestamp 1669390400
transform -1 0 76608 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input60
timestamp 1669390400
transform -1 0 74592 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input61
timestamp 1669390400
transform -1 0 76608 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input62
timestamp 1669390400
transform -1 0 76608 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input63
timestamp 1669390400
transform -1 0 76608 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input64
timestamp 1669390400
transform -1 0 76608 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input65
timestamp 1669390400
transform -1 0 76608 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input66
timestamp 1669390400
transform -1 0 76608 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input67
timestamp 1669390400
transform -1 0 76608 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input68
timestamp 1669390400
transform 1 0 1680 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input69
timestamp 1669390400
transform 1 0 1680 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input70
timestamp 1669390400
transform 1 0 1680 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input71
timestamp 1669390400
transform 1 0 1680 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input72
timestamp 1669390400
transform 1 0 1680 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input73
timestamp 1669390400
transform 1 0 1680 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input74
timestamp 1669390400
transform 1 0 1680 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input75
timestamp 1669390400
transform 1 0 3696 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input76
timestamp 1669390400
transform 1 0 1680 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input77
timestamp 1669390400
transform 1 0 1680 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input78
timestamp 1669390400
transform 1 0 1680 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input79
timestamp 1669390400
transform 1 0 1680 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input80
timestamp 1669390400
transform 1 0 1680 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input81
timestamp 1669390400
transform 1 0 1680 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input82
timestamp 1669390400
transform 1 0 1680 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input83
timestamp 1669390400
transform 1 0 3696 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input84
timestamp 1669390400
transform 1 0 1680 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input85
timestamp 1669390400
transform 1 0 1680 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input86
timestamp 1669390400
transform 1 0 1680 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input87
timestamp 1669390400
transform 1 0 1680 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input88
timestamp 1669390400
transform 1 0 1680 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input89
timestamp 1669390400
transform 1 0 1680 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input90
timestamp 1669390400
transform 1 0 1680 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input91
timestamp 1669390400
transform 1 0 3696 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input92
timestamp 1669390400
transform 1 0 1680 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input93
timestamp 1669390400
transform 1 0 1680 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input94
timestamp 1669390400
transform 1 0 1680 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input95
timestamp 1669390400
transform 1 0 1680 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input96
timestamp 1669390400
transform 1 0 1680 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input97
timestamp 1669390400
transform 1 0 1680 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input98
timestamp 1669390400
transform 1 0 1680 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input99
timestamp 1669390400
transform 1 0 1680 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input100
timestamp 1669390400
transform -1 0 28672 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input101
timestamp 1669390400
transform 1 0 30800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input102
timestamp 1669390400
transform 1 0 33152 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input103
timestamp 1669390400
transform 1 0 34944 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input104
timestamp 1669390400
transform -1 0 36960 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input105
timestamp 1669390400
transform 1 0 34944 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input106
timestamp 1669390400
transform 1 0 34720 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input107
timestamp 1669390400
transform -1 0 38752 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input108
timestamp 1669390400
transform 1 0 38304 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input109
timestamp 1669390400
transform -1 0 40768 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input110
timestamp 1669390400
transform -1 0 40432 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input111
timestamp 1669390400
transform -1 0 29008 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input112
timestamp 1669390400
transform -1 0 42112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input113
timestamp 1669390400
transform 1 0 41440 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input114
timestamp 1669390400
transform -1 0 43456 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input115
timestamp 1669390400
transform 1 0 42336 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input116
timestamp 1669390400
transform -1 0 45248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input117
timestamp 1669390400
transform -1 0 46592 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input118
timestamp 1669390400
transform 1 0 45472 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input119
timestamp 1669390400
transform 1 0 45360 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input120
timestamp 1669390400
transform -1 0 50512 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input121
timestamp 1669390400
transform 1 0 47376 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input122
timestamp 1669390400
transform -1 0 29008 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input123
timestamp 1669390400
transform 1 0 47040 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input124
timestamp 1669390400
transform -1 0 51184 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input125
timestamp 1669390400
transform -1 0 29008 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input126
timestamp 1669390400
transform -1 0 31024 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input127
timestamp 1669390400
transform 1 0 26880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input128
timestamp 1669390400
transform 1 0 29232 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input129
timestamp 1669390400
transform -1 0 33040 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input130
timestamp 1669390400
transform -1 0 32928 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input131
timestamp 1669390400
transform -1 0 33040 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input132
timestamp 1669390400
transform 1 0 70560 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input133
timestamp 1669390400
transform -1 0 74032 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input134
timestamp 1669390400
transform 1 0 71904 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input135
timestamp 1669390400
transform -1 0 75040 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input136
timestamp 1669390400
transform -1 0 75712 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input137
timestamp 1669390400
transform 1 0 69888 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output138 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 76160 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output139
timestamp 1669390400
transform 1 0 76608 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output140
timestamp 1669390400
transform 1 0 74816 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output141
timestamp 1669390400
transform 1 0 74816 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output142
timestamp 1669390400
transform 1 0 74816 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output143
timestamp 1669390400
transform 1 0 74816 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output144
timestamp 1669390400
transform 1 0 74816 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output145
timestamp 1669390400
transform 1 0 74816 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output146
timestamp 1669390400
transform 1 0 76608 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output147
timestamp 1669390400
transform 1 0 74816 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output148
timestamp 1669390400
transform 1 0 74816 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output149
timestamp 1669390400
transform 1 0 74816 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output150
timestamp 1669390400
transform 1 0 74816 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output151
timestamp 1669390400
transform 1 0 74816 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output152
timestamp 1669390400
transform 1 0 74816 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output153
timestamp 1669390400
transform 1 0 74816 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output154
timestamp 1669390400
transform 1 0 76608 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output155
timestamp 1669390400
transform 1 0 74816 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output156
timestamp 1669390400
transform 1 0 74816 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output157
timestamp 1669390400
transform 1 0 74816 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output158
timestamp 1669390400
transform 1 0 74816 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output159
timestamp 1669390400
transform 1 0 74816 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output160
timestamp 1669390400
transform 1 0 74816 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output161
timestamp 1669390400
transform 1 0 76608 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output162
timestamp 1669390400
transform 1 0 76608 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output163
timestamp 1669390400
transform 1 0 74816 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output164
timestamp 1669390400
transform 1 0 74816 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output165
timestamp 1669390400
transform 1 0 74816 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output166
timestamp 1669390400
transform 1 0 74816 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output167
timestamp 1669390400
transform 1 0 74816 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output168
timestamp 1669390400
transform 1 0 74816 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output169
timestamp 1669390400
transform 1 0 74816 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output170
timestamp 1669390400
transform 1 0 76608 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output171
timestamp 1669390400
transform -1 0 3248 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output172
timestamp 1669390400
transform -1 0 3248 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output173
timestamp 1669390400
transform -1 0 3248 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output174
timestamp 1669390400
transform -1 0 3248 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output175
timestamp 1669390400
transform -1 0 3248 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output176
timestamp 1669390400
transform -1 0 3248 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output177
timestamp 1669390400
transform -1 0 3248 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output178
timestamp 1669390400
transform -1 0 5040 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output179
timestamp 1669390400
transform -1 0 3248 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output180
timestamp 1669390400
transform -1 0 3248 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output181
timestamp 1669390400
transform -1 0 3248 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output182
timestamp 1669390400
transform -1 0 3248 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output183
timestamp 1669390400
transform -1 0 3248 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output184
timestamp 1669390400
transform -1 0 3248 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output185
timestamp 1669390400
transform -1 0 3248 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output186
timestamp 1669390400
transform -1 0 5040 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output187
timestamp 1669390400
transform -1 0 3248 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output188
timestamp 1669390400
transform -1 0 3248 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output189
timestamp 1669390400
transform -1 0 3248 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output190
timestamp 1669390400
transform -1 0 3248 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output191
timestamp 1669390400
transform -1 0 3248 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output192
timestamp 1669390400
transform -1 0 3248 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output193
timestamp 1669390400
transform -1 0 5040 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output194
timestamp 1669390400
transform -1 0 5040 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output195
timestamp 1669390400
transform -1 0 3248 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output196
timestamp 1669390400
transform -1 0 3248 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output197
timestamp 1669390400
transform -1 0 3248 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output198
timestamp 1669390400
transform -1 0 3248 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output199
timestamp 1669390400
transform -1 0 3248 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output200
timestamp 1669390400
transform -1 0 3248 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output201
timestamp 1669390400
transform -1 0 3248 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output202
timestamp 1669390400
transform -1 0 5040 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output203
timestamp 1669390400
transform 1 0 74816 0 1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output204
timestamp 1669390400
transform -1 0 3248 0 1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output205
timestamp 1669390400
transform -1 0 50960 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output206
timestamp 1669390400
transform 1 0 55104 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output207
timestamp 1669390400
transform 1 0 57344 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output208
timestamp 1669390400
transform 1 0 58352 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output209
timestamp 1669390400
transform -1 0 58688 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output210
timestamp 1669390400
transform 1 0 59136 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output211
timestamp 1669390400
transform 1 0 60480 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output212
timestamp 1669390400
transform 1 0 59136 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output213
timestamp 1669390400
transform 1 0 60928 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output214
timestamp 1669390400
transform 1 0 62272 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output215
timestamp 1669390400
transform 1 0 61264 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output216
timestamp 1669390400
transform -1 0 50960 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output217
timestamp 1669390400
transform -1 0 64288 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output218
timestamp 1669390400
transform 1 0 64400 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output219
timestamp 1669390400
transform -1 0 64736 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output220
timestamp 1669390400
transform 1 0 65296 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output221
timestamp 1669390400
transform -1 0 67760 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output222
timestamp 1669390400
transform -1 0 66752 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output223
timestamp 1669390400
transform -1 0 68656 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output224
timestamp 1669390400
transform 1 0 66976 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output225
timestamp 1669390400
transform 1 0 67200 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output226
timestamp 1669390400
transform 1 0 69216 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output227
timestamp 1669390400
transform 1 0 51408 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output228
timestamp 1669390400
transform -1 0 70560 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output229
timestamp 1669390400
transform 1 0 69216 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output230
timestamp 1669390400
transform 1 0 52640 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output231
timestamp 1669390400
transform 1 0 51184 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output232
timestamp 1669390400
transform 1 0 53200 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output233
timestamp 1669390400
transform 1 0 54432 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output234
timestamp 1669390400
transform -1 0 54880 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output235
timestamp 1669390400
transform -1 0 56560 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output236
timestamp 1669390400
transform 1 0 56560 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output237
timestamp 1669390400
transform 1 0 74816 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output238
timestamp 1669390400
transform 1 0 74816 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output239
timestamp 1669390400
transform 1 0 74816 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output240
timestamp 1669390400
transform 1 0 76608 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output241
timestamp 1669390400
transform 1 0 74816 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output242
timestamp 1669390400
transform 1 0 74816 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output243
timestamp 1669390400
transform 1 0 74816 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output244
timestamp 1669390400
transform 1 0 74816 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output245
timestamp 1669390400
transform 1 0 74816 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output246
timestamp 1669390400
transform 1 0 74816 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output247
timestamp 1669390400
transform 1 0 74816 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output248
timestamp 1669390400
transform 1 0 74816 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output249
timestamp 1669390400
transform 1 0 74816 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output250
timestamp 1669390400
transform 1 0 74816 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output251
timestamp 1669390400
transform 1 0 74816 0 -1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output252
timestamp 1669390400
transform 1 0 74816 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output253
timestamp 1669390400
transform 1 0 74816 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output254
timestamp 1669390400
transform 1 0 74816 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output255
timestamp 1669390400
transform 1 0 74816 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output256
timestamp 1669390400
transform 1 0 74816 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output257
timestamp 1669390400
transform 1 0 74816 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output258
timestamp 1669390400
transform 1 0 74816 0 1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output259
timestamp 1669390400
transform 1 0 74816 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output260
timestamp 1669390400
transform 1 0 74816 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output261
timestamp 1669390400
transform 1 0 76608 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output262
timestamp 1669390400
transform 1 0 74816 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output263
timestamp 1669390400
transform 1 0 74816 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output264
timestamp 1669390400
transform 1 0 76608 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output265
timestamp 1669390400
transform 1 0 74816 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output266
timestamp 1669390400
transform 1 0 74816 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output267
timestamp 1669390400
transform 1 0 74816 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output268
timestamp 1669390400
transform 1 0 74816 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output269
timestamp 1669390400
transform -1 0 3248 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output270
timestamp 1669390400
transform -1 0 3248 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output271
timestamp 1669390400
transform -1 0 3248 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output272
timestamp 1669390400
transform -1 0 5040 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output273
timestamp 1669390400
transform -1 0 3248 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output274
timestamp 1669390400
transform -1 0 3248 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output275
timestamp 1669390400
transform -1 0 3248 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output276
timestamp 1669390400
transform -1 0 3248 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output277
timestamp 1669390400
transform -1 0 3248 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output278
timestamp 1669390400
transform -1 0 3248 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output279
timestamp 1669390400
transform -1 0 3248 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output280
timestamp 1669390400
transform -1 0 3248 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output281
timestamp 1669390400
transform -1 0 3248 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output282
timestamp 1669390400
transform -1 0 3248 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output283
timestamp 1669390400
transform -1 0 3248 0 -1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output284
timestamp 1669390400
transform -1 0 3248 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output285
timestamp 1669390400
transform -1 0 3248 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output286
timestamp 1669390400
transform -1 0 3248 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output287
timestamp 1669390400
transform -1 0 3248 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output288
timestamp 1669390400
transform -1 0 3248 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output289
timestamp 1669390400
transform -1 0 3248 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output290
timestamp 1669390400
transform -1 0 3248 0 1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output291
timestamp 1669390400
transform -1 0 3248 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output292
timestamp 1669390400
transform -1 0 3248 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output293
timestamp 1669390400
transform -1 0 5040 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output294
timestamp 1669390400
transform -1 0 3248 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output295
timestamp 1669390400
transform -1 0 3248 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output296
timestamp 1669390400
transform -1 0 5040 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output297
timestamp 1669390400
transform -1 0 3248 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output298
timestamp 1669390400
transform -1 0 3248 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output299
timestamp 1669390400
transform -1 0 3248 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output300
timestamp 1669390400
transform -1 0 3248 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output301
timestamp 1669390400
transform 1 0 74816 0 1 72128
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output302
timestamp 1669390400
transform 1 0 76608 0 -1 72128
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output303
timestamp 1669390400
transform 1 0 74816 0 -1 73696
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output304
timestamp 1669390400
transform 1 0 76608 0 -1 73696
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output305
timestamp 1669390400
transform -1 0 3248 0 1 72128
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output306
timestamp 1669390400
transform -1 0 5040 0 -1 72128
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output307
timestamp 1669390400
transform -1 0 3248 0 -1 73696
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output308
timestamp 1669390400
transform -1 0 5040 0 -1 73696
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output309
timestamp 1669390400
transform 1 0 74816 0 -1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output310
timestamp 1669390400
transform -1 0 3248 0 -1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output311
timestamp 1669390400
transform 1 0 74816 0 -1 72128
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output312
timestamp 1669390400
transform -1 0 3248 0 -1 72128
box -86 -86 1654 870
<< labels >>
flabel metal2 s 73808 0 73920 800 0 FreeSans 448 90 0 0 io_wbs_ack
port 0 nsew signal tristate
flabel metal3 s 79200 73808 80000 73920 0 FreeSans 448 0 0 0 io_wbs_ack_0
port 1 nsew signal input
flabel metal3 s 0 73808 800 73920 0 FreeSans 448 0 0 0 io_wbs_ack_1
port 2 nsew signal input
flabel metal2 s 5264 0 5376 800 0 FreeSans 448 90 0 0 io_wbs_adr[0]
port 3 nsew signal input
flabel metal2 s 11984 0 12096 800 0 FreeSans 448 90 0 0 io_wbs_adr[10]
port 4 nsew signal input
flabel metal2 s 12656 0 12768 800 0 FreeSans 448 90 0 0 io_wbs_adr[11]
port 5 nsew signal input
flabel metal2 s 13328 0 13440 800 0 FreeSans 448 90 0 0 io_wbs_adr[12]
port 6 nsew signal input
flabel metal2 s 14000 0 14112 800 0 FreeSans 448 90 0 0 io_wbs_adr[13]
port 7 nsew signal input
flabel metal2 s 14672 0 14784 800 0 FreeSans 448 90 0 0 io_wbs_adr[14]
port 8 nsew signal input
flabel metal2 s 15344 0 15456 800 0 FreeSans 448 90 0 0 io_wbs_adr[15]
port 9 nsew signal input
flabel metal2 s 16016 0 16128 800 0 FreeSans 448 90 0 0 io_wbs_adr[16]
port 10 nsew signal input
flabel metal2 s 16688 0 16800 800 0 FreeSans 448 90 0 0 io_wbs_adr[17]
port 11 nsew signal input
flabel metal2 s 17360 0 17472 800 0 FreeSans 448 90 0 0 io_wbs_adr[18]
port 12 nsew signal input
flabel metal2 s 18032 0 18144 800 0 FreeSans 448 90 0 0 io_wbs_adr[19]
port 13 nsew signal input
flabel metal2 s 5936 0 6048 800 0 FreeSans 448 90 0 0 io_wbs_adr[1]
port 14 nsew signal input
flabel metal2 s 18704 0 18816 800 0 FreeSans 448 90 0 0 io_wbs_adr[20]
port 15 nsew signal input
flabel metal2 s 19376 0 19488 800 0 FreeSans 448 90 0 0 io_wbs_adr[21]
port 16 nsew signal input
flabel metal2 s 20048 0 20160 800 0 FreeSans 448 90 0 0 io_wbs_adr[22]
port 17 nsew signal input
flabel metal2 s 20720 0 20832 800 0 FreeSans 448 90 0 0 io_wbs_adr[23]
port 18 nsew signal input
flabel metal2 s 21392 0 21504 800 0 FreeSans 448 90 0 0 io_wbs_adr[24]
port 19 nsew signal input
flabel metal2 s 22064 0 22176 800 0 FreeSans 448 90 0 0 io_wbs_adr[25]
port 20 nsew signal input
flabel metal2 s 22736 0 22848 800 0 FreeSans 448 90 0 0 io_wbs_adr[26]
port 21 nsew signal input
flabel metal2 s 23408 0 23520 800 0 FreeSans 448 90 0 0 io_wbs_adr[27]
port 22 nsew signal input
flabel metal2 s 24080 0 24192 800 0 FreeSans 448 90 0 0 io_wbs_adr[28]
port 23 nsew signal input
flabel metal2 s 24752 0 24864 800 0 FreeSans 448 90 0 0 io_wbs_adr[29]
port 24 nsew signal input
flabel metal2 s 6608 0 6720 800 0 FreeSans 448 90 0 0 io_wbs_adr[2]
port 25 nsew signal input
flabel metal2 s 25424 0 25536 800 0 FreeSans 448 90 0 0 io_wbs_adr[30]
port 26 nsew signal input
flabel metal2 s 26096 0 26208 800 0 FreeSans 448 90 0 0 io_wbs_adr[31]
port 27 nsew signal input
flabel metal2 s 7280 0 7392 800 0 FreeSans 448 90 0 0 io_wbs_adr[3]
port 28 nsew signal input
flabel metal2 s 7952 0 8064 800 0 FreeSans 448 90 0 0 io_wbs_adr[4]
port 29 nsew signal input
flabel metal2 s 8624 0 8736 800 0 FreeSans 448 90 0 0 io_wbs_adr[5]
port 30 nsew signal input
flabel metal2 s 9296 0 9408 800 0 FreeSans 448 90 0 0 io_wbs_adr[6]
port 31 nsew signal input
flabel metal2 s 9968 0 10080 800 0 FreeSans 448 90 0 0 io_wbs_adr[7]
port 32 nsew signal input
flabel metal2 s 10640 0 10752 800 0 FreeSans 448 90 0 0 io_wbs_adr[8]
port 33 nsew signal input
flabel metal2 s 11312 0 11424 800 0 FreeSans 448 90 0 0 io_wbs_adr[9]
port 34 nsew signal input
flabel metal3 s 79200 5264 80000 5376 0 FreeSans 448 0 0 0 io_wbs_adr_0[0]
port 35 nsew signal tristate
flabel metal3 s 79200 11984 80000 12096 0 FreeSans 448 0 0 0 io_wbs_adr_0[10]
port 36 nsew signal tristate
flabel metal3 s 79200 12656 80000 12768 0 FreeSans 448 0 0 0 io_wbs_adr_0[11]
port 37 nsew signal tristate
flabel metal3 s 79200 13328 80000 13440 0 FreeSans 448 0 0 0 io_wbs_adr_0[12]
port 38 nsew signal tristate
flabel metal3 s 79200 14000 80000 14112 0 FreeSans 448 0 0 0 io_wbs_adr_0[13]
port 39 nsew signal tristate
flabel metal3 s 79200 14672 80000 14784 0 FreeSans 448 0 0 0 io_wbs_adr_0[14]
port 40 nsew signal tristate
flabel metal3 s 79200 15344 80000 15456 0 FreeSans 448 0 0 0 io_wbs_adr_0[15]
port 41 nsew signal tristate
flabel metal3 s 79200 16016 80000 16128 0 FreeSans 448 0 0 0 io_wbs_adr_0[16]
port 42 nsew signal tristate
flabel metal3 s 79200 16688 80000 16800 0 FreeSans 448 0 0 0 io_wbs_adr_0[17]
port 43 nsew signal tristate
flabel metal3 s 79200 17360 80000 17472 0 FreeSans 448 0 0 0 io_wbs_adr_0[18]
port 44 nsew signal tristate
flabel metal3 s 79200 18032 80000 18144 0 FreeSans 448 0 0 0 io_wbs_adr_0[19]
port 45 nsew signal tristate
flabel metal3 s 79200 5936 80000 6048 0 FreeSans 448 0 0 0 io_wbs_adr_0[1]
port 46 nsew signal tristate
flabel metal3 s 79200 18704 80000 18816 0 FreeSans 448 0 0 0 io_wbs_adr_0[20]
port 47 nsew signal tristate
flabel metal3 s 79200 19376 80000 19488 0 FreeSans 448 0 0 0 io_wbs_adr_0[21]
port 48 nsew signal tristate
flabel metal3 s 79200 20048 80000 20160 0 FreeSans 448 0 0 0 io_wbs_adr_0[22]
port 49 nsew signal tristate
flabel metal3 s 79200 20720 80000 20832 0 FreeSans 448 0 0 0 io_wbs_adr_0[23]
port 50 nsew signal tristate
flabel metal3 s 79200 21392 80000 21504 0 FreeSans 448 0 0 0 io_wbs_adr_0[24]
port 51 nsew signal tristate
flabel metal3 s 79200 22064 80000 22176 0 FreeSans 448 0 0 0 io_wbs_adr_0[25]
port 52 nsew signal tristate
flabel metal3 s 79200 22736 80000 22848 0 FreeSans 448 0 0 0 io_wbs_adr_0[26]
port 53 nsew signal tristate
flabel metal3 s 79200 23408 80000 23520 0 FreeSans 448 0 0 0 io_wbs_adr_0[27]
port 54 nsew signal tristate
flabel metal3 s 79200 24080 80000 24192 0 FreeSans 448 0 0 0 io_wbs_adr_0[28]
port 55 nsew signal tristate
flabel metal3 s 79200 24752 80000 24864 0 FreeSans 448 0 0 0 io_wbs_adr_0[29]
port 56 nsew signal tristate
flabel metal3 s 79200 6608 80000 6720 0 FreeSans 448 0 0 0 io_wbs_adr_0[2]
port 57 nsew signal tristate
flabel metal3 s 79200 25424 80000 25536 0 FreeSans 448 0 0 0 io_wbs_adr_0[30]
port 58 nsew signal tristate
flabel metal3 s 79200 26096 80000 26208 0 FreeSans 448 0 0 0 io_wbs_adr_0[31]
port 59 nsew signal tristate
flabel metal3 s 79200 7280 80000 7392 0 FreeSans 448 0 0 0 io_wbs_adr_0[3]
port 60 nsew signal tristate
flabel metal3 s 79200 7952 80000 8064 0 FreeSans 448 0 0 0 io_wbs_adr_0[4]
port 61 nsew signal tristate
flabel metal3 s 79200 8624 80000 8736 0 FreeSans 448 0 0 0 io_wbs_adr_0[5]
port 62 nsew signal tristate
flabel metal3 s 79200 9296 80000 9408 0 FreeSans 448 0 0 0 io_wbs_adr_0[6]
port 63 nsew signal tristate
flabel metal3 s 79200 9968 80000 10080 0 FreeSans 448 0 0 0 io_wbs_adr_0[7]
port 64 nsew signal tristate
flabel metal3 s 79200 10640 80000 10752 0 FreeSans 448 0 0 0 io_wbs_adr_0[8]
port 65 nsew signal tristate
flabel metal3 s 79200 11312 80000 11424 0 FreeSans 448 0 0 0 io_wbs_adr_0[9]
port 66 nsew signal tristate
flabel metal3 s 0 5264 800 5376 0 FreeSans 448 0 0 0 io_wbs_adr_1[0]
port 67 nsew signal tristate
flabel metal3 s 0 11984 800 12096 0 FreeSans 448 0 0 0 io_wbs_adr_1[10]
port 68 nsew signal tristate
flabel metal3 s 0 12656 800 12768 0 FreeSans 448 0 0 0 io_wbs_adr_1[11]
port 69 nsew signal tristate
flabel metal3 s 0 13328 800 13440 0 FreeSans 448 0 0 0 io_wbs_adr_1[12]
port 70 nsew signal tristate
flabel metal3 s 0 14000 800 14112 0 FreeSans 448 0 0 0 io_wbs_adr_1[13]
port 71 nsew signal tristate
flabel metal3 s 0 14672 800 14784 0 FreeSans 448 0 0 0 io_wbs_adr_1[14]
port 72 nsew signal tristate
flabel metal3 s 0 15344 800 15456 0 FreeSans 448 0 0 0 io_wbs_adr_1[15]
port 73 nsew signal tristate
flabel metal3 s 0 16016 800 16128 0 FreeSans 448 0 0 0 io_wbs_adr_1[16]
port 74 nsew signal tristate
flabel metal3 s 0 16688 800 16800 0 FreeSans 448 0 0 0 io_wbs_adr_1[17]
port 75 nsew signal tristate
flabel metal3 s 0 17360 800 17472 0 FreeSans 448 0 0 0 io_wbs_adr_1[18]
port 76 nsew signal tristate
flabel metal3 s 0 18032 800 18144 0 FreeSans 448 0 0 0 io_wbs_adr_1[19]
port 77 nsew signal tristate
flabel metal3 s 0 5936 800 6048 0 FreeSans 448 0 0 0 io_wbs_adr_1[1]
port 78 nsew signal tristate
flabel metal3 s 0 18704 800 18816 0 FreeSans 448 0 0 0 io_wbs_adr_1[20]
port 79 nsew signal tristate
flabel metal3 s 0 19376 800 19488 0 FreeSans 448 0 0 0 io_wbs_adr_1[21]
port 80 nsew signal tristate
flabel metal3 s 0 20048 800 20160 0 FreeSans 448 0 0 0 io_wbs_adr_1[22]
port 81 nsew signal tristate
flabel metal3 s 0 20720 800 20832 0 FreeSans 448 0 0 0 io_wbs_adr_1[23]
port 82 nsew signal tristate
flabel metal3 s 0 21392 800 21504 0 FreeSans 448 0 0 0 io_wbs_adr_1[24]
port 83 nsew signal tristate
flabel metal3 s 0 22064 800 22176 0 FreeSans 448 0 0 0 io_wbs_adr_1[25]
port 84 nsew signal tristate
flabel metal3 s 0 22736 800 22848 0 FreeSans 448 0 0 0 io_wbs_adr_1[26]
port 85 nsew signal tristate
flabel metal3 s 0 23408 800 23520 0 FreeSans 448 0 0 0 io_wbs_adr_1[27]
port 86 nsew signal tristate
flabel metal3 s 0 24080 800 24192 0 FreeSans 448 0 0 0 io_wbs_adr_1[28]
port 87 nsew signal tristate
flabel metal3 s 0 24752 800 24864 0 FreeSans 448 0 0 0 io_wbs_adr_1[29]
port 88 nsew signal tristate
flabel metal3 s 0 6608 800 6720 0 FreeSans 448 0 0 0 io_wbs_adr_1[2]
port 89 nsew signal tristate
flabel metal3 s 0 25424 800 25536 0 FreeSans 448 0 0 0 io_wbs_adr_1[30]
port 90 nsew signal tristate
flabel metal3 s 0 26096 800 26208 0 FreeSans 448 0 0 0 io_wbs_adr_1[31]
port 91 nsew signal tristate
flabel metal3 s 0 7280 800 7392 0 FreeSans 448 0 0 0 io_wbs_adr_1[3]
port 92 nsew signal tristate
flabel metal3 s 0 7952 800 8064 0 FreeSans 448 0 0 0 io_wbs_adr_1[4]
port 93 nsew signal tristate
flabel metal3 s 0 8624 800 8736 0 FreeSans 448 0 0 0 io_wbs_adr_1[5]
port 94 nsew signal tristate
flabel metal3 s 0 9296 800 9408 0 FreeSans 448 0 0 0 io_wbs_adr_1[6]
port 95 nsew signal tristate
flabel metal3 s 0 9968 800 10080 0 FreeSans 448 0 0 0 io_wbs_adr_1[7]
port 96 nsew signal tristate
flabel metal3 s 0 10640 800 10752 0 FreeSans 448 0 0 0 io_wbs_adr_1[8]
port 97 nsew signal tristate
flabel metal3 s 0 11312 800 11424 0 FreeSans 448 0 0 0 io_wbs_adr_1[9]
port 98 nsew signal tristate
flabel metal2 s 74480 0 74592 800 0 FreeSans 448 90 0 0 io_wbs_cyc
port 99 nsew signal input
flabel metal3 s 79200 74480 80000 74592 0 FreeSans 448 0 0 0 io_wbs_cyc_0
port 100 nsew signal tristate
flabel metal3 s 0 74480 800 74592 0 FreeSans 448 0 0 0 io_wbs_cyc_1
port 101 nsew signal tristate
flabel metal2 s 48272 0 48384 800 0 FreeSans 448 90 0 0 io_wbs_datrd[0]
port 102 nsew signal tristate
flabel metal2 s 54992 0 55104 800 0 FreeSans 448 90 0 0 io_wbs_datrd[10]
port 103 nsew signal tristate
flabel metal2 s 55664 0 55776 800 0 FreeSans 448 90 0 0 io_wbs_datrd[11]
port 104 nsew signal tristate
flabel metal2 s 56336 0 56448 800 0 FreeSans 448 90 0 0 io_wbs_datrd[12]
port 105 nsew signal tristate
flabel metal2 s 57008 0 57120 800 0 FreeSans 448 90 0 0 io_wbs_datrd[13]
port 106 nsew signal tristate
flabel metal2 s 57680 0 57792 800 0 FreeSans 448 90 0 0 io_wbs_datrd[14]
port 107 nsew signal tristate
flabel metal2 s 58352 0 58464 800 0 FreeSans 448 90 0 0 io_wbs_datrd[15]
port 108 nsew signal tristate
flabel metal2 s 59024 0 59136 800 0 FreeSans 448 90 0 0 io_wbs_datrd[16]
port 109 nsew signal tristate
flabel metal2 s 59696 0 59808 800 0 FreeSans 448 90 0 0 io_wbs_datrd[17]
port 110 nsew signal tristate
flabel metal2 s 60368 0 60480 800 0 FreeSans 448 90 0 0 io_wbs_datrd[18]
port 111 nsew signal tristate
flabel metal2 s 61040 0 61152 800 0 FreeSans 448 90 0 0 io_wbs_datrd[19]
port 112 nsew signal tristate
flabel metal2 s 48944 0 49056 800 0 FreeSans 448 90 0 0 io_wbs_datrd[1]
port 113 nsew signal tristate
flabel metal2 s 61712 0 61824 800 0 FreeSans 448 90 0 0 io_wbs_datrd[20]
port 114 nsew signal tristate
flabel metal2 s 62384 0 62496 800 0 FreeSans 448 90 0 0 io_wbs_datrd[21]
port 115 nsew signal tristate
flabel metal2 s 63056 0 63168 800 0 FreeSans 448 90 0 0 io_wbs_datrd[22]
port 116 nsew signal tristate
flabel metal2 s 63728 0 63840 800 0 FreeSans 448 90 0 0 io_wbs_datrd[23]
port 117 nsew signal tristate
flabel metal2 s 64400 0 64512 800 0 FreeSans 448 90 0 0 io_wbs_datrd[24]
port 118 nsew signal tristate
flabel metal2 s 65072 0 65184 800 0 FreeSans 448 90 0 0 io_wbs_datrd[25]
port 119 nsew signal tristate
flabel metal2 s 65744 0 65856 800 0 FreeSans 448 90 0 0 io_wbs_datrd[26]
port 120 nsew signal tristate
flabel metal2 s 66416 0 66528 800 0 FreeSans 448 90 0 0 io_wbs_datrd[27]
port 121 nsew signal tristate
flabel metal2 s 67088 0 67200 800 0 FreeSans 448 90 0 0 io_wbs_datrd[28]
port 122 nsew signal tristate
flabel metal2 s 67760 0 67872 800 0 FreeSans 448 90 0 0 io_wbs_datrd[29]
port 123 nsew signal tristate
flabel metal2 s 49616 0 49728 800 0 FreeSans 448 90 0 0 io_wbs_datrd[2]
port 124 nsew signal tristate
flabel metal2 s 68432 0 68544 800 0 FreeSans 448 90 0 0 io_wbs_datrd[30]
port 125 nsew signal tristate
flabel metal2 s 69104 0 69216 800 0 FreeSans 448 90 0 0 io_wbs_datrd[31]
port 126 nsew signal tristate
flabel metal2 s 50288 0 50400 800 0 FreeSans 448 90 0 0 io_wbs_datrd[3]
port 127 nsew signal tristate
flabel metal2 s 50960 0 51072 800 0 FreeSans 448 90 0 0 io_wbs_datrd[4]
port 128 nsew signal tristate
flabel metal2 s 51632 0 51744 800 0 FreeSans 448 90 0 0 io_wbs_datrd[5]
port 129 nsew signal tristate
flabel metal2 s 52304 0 52416 800 0 FreeSans 448 90 0 0 io_wbs_datrd[6]
port 130 nsew signal tristate
flabel metal2 s 52976 0 53088 800 0 FreeSans 448 90 0 0 io_wbs_datrd[7]
port 131 nsew signal tristate
flabel metal2 s 53648 0 53760 800 0 FreeSans 448 90 0 0 io_wbs_datrd[8]
port 132 nsew signal tristate
flabel metal2 s 54320 0 54432 800 0 FreeSans 448 90 0 0 io_wbs_datrd[9]
port 133 nsew signal tristate
flabel metal3 s 79200 48272 80000 48384 0 FreeSans 448 0 0 0 io_wbs_datrd_0[0]
port 134 nsew signal input
flabel metal3 s 79200 54992 80000 55104 0 FreeSans 448 0 0 0 io_wbs_datrd_0[10]
port 135 nsew signal input
flabel metal3 s 79200 55664 80000 55776 0 FreeSans 448 0 0 0 io_wbs_datrd_0[11]
port 136 nsew signal input
flabel metal3 s 79200 56336 80000 56448 0 FreeSans 448 0 0 0 io_wbs_datrd_0[12]
port 137 nsew signal input
flabel metal3 s 79200 57008 80000 57120 0 FreeSans 448 0 0 0 io_wbs_datrd_0[13]
port 138 nsew signal input
flabel metal3 s 79200 57680 80000 57792 0 FreeSans 448 0 0 0 io_wbs_datrd_0[14]
port 139 nsew signal input
flabel metal3 s 79200 58352 80000 58464 0 FreeSans 448 0 0 0 io_wbs_datrd_0[15]
port 140 nsew signal input
flabel metal3 s 79200 59024 80000 59136 0 FreeSans 448 0 0 0 io_wbs_datrd_0[16]
port 141 nsew signal input
flabel metal3 s 79200 59696 80000 59808 0 FreeSans 448 0 0 0 io_wbs_datrd_0[17]
port 142 nsew signal input
flabel metal3 s 79200 60368 80000 60480 0 FreeSans 448 0 0 0 io_wbs_datrd_0[18]
port 143 nsew signal input
flabel metal3 s 79200 61040 80000 61152 0 FreeSans 448 0 0 0 io_wbs_datrd_0[19]
port 144 nsew signal input
flabel metal3 s 79200 48944 80000 49056 0 FreeSans 448 0 0 0 io_wbs_datrd_0[1]
port 145 nsew signal input
flabel metal3 s 79200 61712 80000 61824 0 FreeSans 448 0 0 0 io_wbs_datrd_0[20]
port 146 nsew signal input
flabel metal3 s 79200 62384 80000 62496 0 FreeSans 448 0 0 0 io_wbs_datrd_0[21]
port 147 nsew signal input
flabel metal3 s 79200 63056 80000 63168 0 FreeSans 448 0 0 0 io_wbs_datrd_0[22]
port 148 nsew signal input
flabel metal3 s 79200 63728 80000 63840 0 FreeSans 448 0 0 0 io_wbs_datrd_0[23]
port 149 nsew signal input
flabel metal3 s 79200 64400 80000 64512 0 FreeSans 448 0 0 0 io_wbs_datrd_0[24]
port 150 nsew signal input
flabel metal3 s 79200 65072 80000 65184 0 FreeSans 448 0 0 0 io_wbs_datrd_0[25]
port 151 nsew signal input
flabel metal3 s 79200 65744 80000 65856 0 FreeSans 448 0 0 0 io_wbs_datrd_0[26]
port 152 nsew signal input
flabel metal3 s 79200 66416 80000 66528 0 FreeSans 448 0 0 0 io_wbs_datrd_0[27]
port 153 nsew signal input
flabel metal3 s 79200 67088 80000 67200 0 FreeSans 448 0 0 0 io_wbs_datrd_0[28]
port 154 nsew signal input
flabel metal3 s 79200 67760 80000 67872 0 FreeSans 448 0 0 0 io_wbs_datrd_0[29]
port 155 nsew signal input
flabel metal3 s 79200 49616 80000 49728 0 FreeSans 448 0 0 0 io_wbs_datrd_0[2]
port 156 nsew signal input
flabel metal3 s 79200 68432 80000 68544 0 FreeSans 448 0 0 0 io_wbs_datrd_0[30]
port 157 nsew signal input
flabel metal3 s 79200 69104 80000 69216 0 FreeSans 448 0 0 0 io_wbs_datrd_0[31]
port 158 nsew signal input
flabel metal3 s 79200 50288 80000 50400 0 FreeSans 448 0 0 0 io_wbs_datrd_0[3]
port 159 nsew signal input
flabel metal3 s 79200 50960 80000 51072 0 FreeSans 448 0 0 0 io_wbs_datrd_0[4]
port 160 nsew signal input
flabel metal3 s 79200 51632 80000 51744 0 FreeSans 448 0 0 0 io_wbs_datrd_0[5]
port 161 nsew signal input
flabel metal3 s 79200 52304 80000 52416 0 FreeSans 448 0 0 0 io_wbs_datrd_0[6]
port 162 nsew signal input
flabel metal3 s 79200 52976 80000 53088 0 FreeSans 448 0 0 0 io_wbs_datrd_0[7]
port 163 nsew signal input
flabel metal3 s 79200 53648 80000 53760 0 FreeSans 448 0 0 0 io_wbs_datrd_0[8]
port 164 nsew signal input
flabel metal3 s 79200 54320 80000 54432 0 FreeSans 448 0 0 0 io_wbs_datrd_0[9]
port 165 nsew signal input
flabel metal3 s 0 48272 800 48384 0 FreeSans 448 0 0 0 io_wbs_datrd_1[0]
port 166 nsew signal input
flabel metal3 s 0 54992 800 55104 0 FreeSans 448 0 0 0 io_wbs_datrd_1[10]
port 167 nsew signal input
flabel metal3 s 0 55664 800 55776 0 FreeSans 448 0 0 0 io_wbs_datrd_1[11]
port 168 nsew signal input
flabel metal3 s 0 56336 800 56448 0 FreeSans 448 0 0 0 io_wbs_datrd_1[12]
port 169 nsew signal input
flabel metal3 s 0 57008 800 57120 0 FreeSans 448 0 0 0 io_wbs_datrd_1[13]
port 170 nsew signal input
flabel metal3 s 0 57680 800 57792 0 FreeSans 448 0 0 0 io_wbs_datrd_1[14]
port 171 nsew signal input
flabel metal3 s 0 58352 800 58464 0 FreeSans 448 0 0 0 io_wbs_datrd_1[15]
port 172 nsew signal input
flabel metal3 s 0 59024 800 59136 0 FreeSans 448 0 0 0 io_wbs_datrd_1[16]
port 173 nsew signal input
flabel metal3 s 0 59696 800 59808 0 FreeSans 448 0 0 0 io_wbs_datrd_1[17]
port 174 nsew signal input
flabel metal3 s 0 60368 800 60480 0 FreeSans 448 0 0 0 io_wbs_datrd_1[18]
port 175 nsew signal input
flabel metal3 s 0 61040 800 61152 0 FreeSans 448 0 0 0 io_wbs_datrd_1[19]
port 176 nsew signal input
flabel metal3 s 0 48944 800 49056 0 FreeSans 448 0 0 0 io_wbs_datrd_1[1]
port 177 nsew signal input
flabel metal3 s 0 61712 800 61824 0 FreeSans 448 0 0 0 io_wbs_datrd_1[20]
port 178 nsew signal input
flabel metal3 s 0 62384 800 62496 0 FreeSans 448 0 0 0 io_wbs_datrd_1[21]
port 179 nsew signal input
flabel metal3 s 0 63056 800 63168 0 FreeSans 448 0 0 0 io_wbs_datrd_1[22]
port 180 nsew signal input
flabel metal3 s 0 63728 800 63840 0 FreeSans 448 0 0 0 io_wbs_datrd_1[23]
port 181 nsew signal input
flabel metal3 s 0 64400 800 64512 0 FreeSans 448 0 0 0 io_wbs_datrd_1[24]
port 182 nsew signal input
flabel metal3 s 0 65072 800 65184 0 FreeSans 448 0 0 0 io_wbs_datrd_1[25]
port 183 nsew signal input
flabel metal3 s 0 65744 800 65856 0 FreeSans 448 0 0 0 io_wbs_datrd_1[26]
port 184 nsew signal input
flabel metal3 s 0 66416 800 66528 0 FreeSans 448 0 0 0 io_wbs_datrd_1[27]
port 185 nsew signal input
flabel metal3 s 0 67088 800 67200 0 FreeSans 448 0 0 0 io_wbs_datrd_1[28]
port 186 nsew signal input
flabel metal3 s 0 67760 800 67872 0 FreeSans 448 0 0 0 io_wbs_datrd_1[29]
port 187 nsew signal input
flabel metal3 s 0 49616 800 49728 0 FreeSans 448 0 0 0 io_wbs_datrd_1[2]
port 188 nsew signal input
flabel metal3 s 0 68432 800 68544 0 FreeSans 448 0 0 0 io_wbs_datrd_1[30]
port 189 nsew signal input
flabel metal3 s 0 69104 800 69216 0 FreeSans 448 0 0 0 io_wbs_datrd_1[31]
port 190 nsew signal input
flabel metal3 s 0 50288 800 50400 0 FreeSans 448 0 0 0 io_wbs_datrd_1[3]
port 191 nsew signal input
flabel metal3 s 0 50960 800 51072 0 FreeSans 448 0 0 0 io_wbs_datrd_1[4]
port 192 nsew signal input
flabel metal3 s 0 51632 800 51744 0 FreeSans 448 0 0 0 io_wbs_datrd_1[5]
port 193 nsew signal input
flabel metal3 s 0 52304 800 52416 0 FreeSans 448 0 0 0 io_wbs_datrd_1[6]
port 194 nsew signal input
flabel metal3 s 0 52976 800 53088 0 FreeSans 448 0 0 0 io_wbs_datrd_1[7]
port 195 nsew signal input
flabel metal3 s 0 53648 800 53760 0 FreeSans 448 0 0 0 io_wbs_datrd_1[8]
port 196 nsew signal input
flabel metal3 s 0 54320 800 54432 0 FreeSans 448 0 0 0 io_wbs_datrd_1[9]
port 197 nsew signal input
flabel metal2 s 26768 0 26880 800 0 FreeSans 448 90 0 0 io_wbs_datwr[0]
port 198 nsew signal input
flabel metal2 s 33488 0 33600 800 0 FreeSans 448 90 0 0 io_wbs_datwr[10]
port 199 nsew signal input
flabel metal2 s 34160 0 34272 800 0 FreeSans 448 90 0 0 io_wbs_datwr[11]
port 200 nsew signal input
flabel metal2 s 34832 0 34944 800 0 FreeSans 448 90 0 0 io_wbs_datwr[12]
port 201 nsew signal input
flabel metal2 s 35504 0 35616 800 0 FreeSans 448 90 0 0 io_wbs_datwr[13]
port 202 nsew signal input
flabel metal2 s 36176 0 36288 800 0 FreeSans 448 90 0 0 io_wbs_datwr[14]
port 203 nsew signal input
flabel metal2 s 36848 0 36960 800 0 FreeSans 448 90 0 0 io_wbs_datwr[15]
port 204 nsew signal input
flabel metal2 s 37520 0 37632 800 0 FreeSans 448 90 0 0 io_wbs_datwr[16]
port 205 nsew signal input
flabel metal2 s 38192 0 38304 800 0 FreeSans 448 90 0 0 io_wbs_datwr[17]
port 206 nsew signal input
flabel metal2 s 38864 0 38976 800 0 FreeSans 448 90 0 0 io_wbs_datwr[18]
port 207 nsew signal input
flabel metal2 s 39536 0 39648 800 0 FreeSans 448 90 0 0 io_wbs_datwr[19]
port 208 nsew signal input
flabel metal2 s 27440 0 27552 800 0 FreeSans 448 90 0 0 io_wbs_datwr[1]
port 209 nsew signal input
flabel metal2 s 40208 0 40320 800 0 FreeSans 448 90 0 0 io_wbs_datwr[20]
port 210 nsew signal input
flabel metal2 s 40880 0 40992 800 0 FreeSans 448 90 0 0 io_wbs_datwr[21]
port 211 nsew signal input
flabel metal2 s 41552 0 41664 800 0 FreeSans 448 90 0 0 io_wbs_datwr[22]
port 212 nsew signal input
flabel metal2 s 42224 0 42336 800 0 FreeSans 448 90 0 0 io_wbs_datwr[23]
port 213 nsew signal input
flabel metal2 s 42896 0 43008 800 0 FreeSans 448 90 0 0 io_wbs_datwr[24]
port 214 nsew signal input
flabel metal2 s 43568 0 43680 800 0 FreeSans 448 90 0 0 io_wbs_datwr[25]
port 215 nsew signal input
flabel metal2 s 44240 0 44352 800 0 FreeSans 448 90 0 0 io_wbs_datwr[26]
port 216 nsew signal input
flabel metal2 s 44912 0 45024 800 0 FreeSans 448 90 0 0 io_wbs_datwr[27]
port 217 nsew signal input
flabel metal2 s 45584 0 45696 800 0 FreeSans 448 90 0 0 io_wbs_datwr[28]
port 218 nsew signal input
flabel metal2 s 46256 0 46368 800 0 FreeSans 448 90 0 0 io_wbs_datwr[29]
port 219 nsew signal input
flabel metal2 s 28112 0 28224 800 0 FreeSans 448 90 0 0 io_wbs_datwr[2]
port 220 nsew signal input
flabel metal2 s 46928 0 47040 800 0 FreeSans 448 90 0 0 io_wbs_datwr[30]
port 221 nsew signal input
flabel metal2 s 47600 0 47712 800 0 FreeSans 448 90 0 0 io_wbs_datwr[31]
port 222 nsew signal input
flabel metal2 s 28784 0 28896 800 0 FreeSans 448 90 0 0 io_wbs_datwr[3]
port 223 nsew signal input
flabel metal2 s 29456 0 29568 800 0 FreeSans 448 90 0 0 io_wbs_datwr[4]
port 224 nsew signal input
flabel metal2 s 30128 0 30240 800 0 FreeSans 448 90 0 0 io_wbs_datwr[5]
port 225 nsew signal input
flabel metal2 s 30800 0 30912 800 0 FreeSans 448 90 0 0 io_wbs_datwr[6]
port 226 nsew signal input
flabel metal2 s 31472 0 31584 800 0 FreeSans 448 90 0 0 io_wbs_datwr[7]
port 227 nsew signal input
flabel metal2 s 32144 0 32256 800 0 FreeSans 448 90 0 0 io_wbs_datwr[8]
port 228 nsew signal input
flabel metal2 s 32816 0 32928 800 0 FreeSans 448 90 0 0 io_wbs_datwr[9]
port 229 nsew signal input
flabel metal3 s 79200 26768 80000 26880 0 FreeSans 448 0 0 0 io_wbs_datwr_0[0]
port 230 nsew signal tristate
flabel metal3 s 79200 33488 80000 33600 0 FreeSans 448 0 0 0 io_wbs_datwr_0[10]
port 231 nsew signal tristate
flabel metal3 s 79200 34160 80000 34272 0 FreeSans 448 0 0 0 io_wbs_datwr_0[11]
port 232 nsew signal tristate
flabel metal3 s 79200 34832 80000 34944 0 FreeSans 448 0 0 0 io_wbs_datwr_0[12]
port 233 nsew signal tristate
flabel metal3 s 79200 35504 80000 35616 0 FreeSans 448 0 0 0 io_wbs_datwr_0[13]
port 234 nsew signal tristate
flabel metal3 s 79200 36176 80000 36288 0 FreeSans 448 0 0 0 io_wbs_datwr_0[14]
port 235 nsew signal tristate
flabel metal3 s 79200 36848 80000 36960 0 FreeSans 448 0 0 0 io_wbs_datwr_0[15]
port 236 nsew signal tristate
flabel metal3 s 79200 37520 80000 37632 0 FreeSans 448 0 0 0 io_wbs_datwr_0[16]
port 237 nsew signal tristate
flabel metal3 s 79200 38192 80000 38304 0 FreeSans 448 0 0 0 io_wbs_datwr_0[17]
port 238 nsew signal tristate
flabel metal3 s 79200 38864 80000 38976 0 FreeSans 448 0 0 0 io_wbs_datwr_0[18]
port 239 nsew signal tristate
flabel metal3 s 79200 39536 80000 39648 0 FreeSans 448 0 0 0 io_wbs_datwr_0[19]
port 240 nsew signal tristate
flabel metal3 s 79200 27440 80000 27552 0 FreeSans 448 0 0 0 io_wbs_datwr_0[1]
port 241 nsew signal tristate
flabel metal3 s 79200 40208 80000 40320 0 FreeSans 448 0 0 0 io_wbs_datwr_0[20]
port 242 nsew signal tristate
flabel metal3 s 79200 40880 80000 40992 0 FreeSans 448 0 0 0 io_wbs_datwr_0[21]
port 243 nsew signal tristate
flabel metal3 s 79200 41552 80000 41664 0 FreeSans 448 0 0 0 io_wbs_datwr_0[22]
port 244 nsew signal tristate
flabel metal3 s 79200 42224 80000 42336 0 FreeSans 448 0 0 0 io_wbs_datwr_0[23]
port 245 nsew signal tristate
flabel metal3 s 79200 42896 80000 43008 0 FreeSans 448 0 0 0 io_wbs_datwr_0[24]
port 246 nsew signal tristate
flabel metal3 s 79200 43568 80000 43680 0 FreeSans 448 0 0 0 io_wbs_datwr_0[25]
port 247 nsew signal tristate
flabel metal3 s 79200 44240 80000 44352 0 FreeSans 448 0 0 0 io_wbs_datwr_0[26]
port 248 nsew signal tristate
flabel metal3 s 79200 44912 80000 45024 0 FreeSans 448 0 0 0 io_wbs_datwr_0[27]
port 249 nsew signal tristate
flabel metal3 s 79200 45584 80000 45696 0 FreeSans 448 0 0 0 io_wbs_datwr_0[28]
port 250 nsew signal tristate
flabel metal3 s 79200 46256 80000 46368 0 FreeSans 448 0 0 0 io_wbs_datwr_0[29]
port 251 nsew signal tristate
flabel metal3 s 79200 28112 80000 28224 0 FreeSans 448 0 0 0 io_wbs_datwr_0[2]
port 252 nsew signal tristate
flabel metal3 s 79200 46928 80000 47040 0 FreeSans 448 0 0 0 io_wbs_datwr_0[30]
port 253 nsew signal tristate
flabel metal3 s 79200 47600 80000 47712 0 FreeSans 448 0 0 0 io_wbs_datwr_0[31]
port 254 nsew signal tristate
flabel metal3 s 79200 28784 80000 28896 0 FreeSans 448 0 0 0 io_wbs_datwr_0[3]
port 255 nsew signal tristate
flabel metal3 s 79200 29456 80000 29568 0 FreeSans 448 0 0 0 io_wbs_datwr_0[4]
port 256 nsew signal tristate
flabel metal3 s 79200 30128 80000 30240 0 FreeSans 448 0 0 0 io_wbs_datwr_0[5]
port 257 nsew signal tristate
flabel metal3 s 79200 30800 80000 30912 0 FreeSans 448 0 0 0 io_wbs_datwr_0[6]
port 258 nsew signal tristate
flabel metal3 s 79200 31472 80000 31584 0 FreeSans 448 0 0 0 io_wbs_datwr_0[7]
port 259 nsew signal tristate
flabel metal3 s 79200 32144 80000 32256 0 FreeSans 448 0 0 0 io_wbs_datwr_0[8]
port 260 nsew signal tristate
flabel metal3 s 79200 32816 80000 32928 0 FreeSans 448 0 0 0 io_wbs_datwr_0[9]
port 261 nsew signal tristate
flabel metal3 s 0 26768 800 26880 0 FreeSans 448 0 0 0 io_wbs_datwr_1[0]
port 262 nsew signal tristate
flabel metal3 s 0 33488 800 33600 0 FreeSans 448 0 0 0 io_wbs_datwr_1[10]
port 263 nsew signal tristate
flabel metal3 s 0 34160 800 34272 0 FreeSans 448 0 0 0 io_wbs_datwr_1[11]
port 264 nsew signal tristate
flabel metal3 s 0 34832 800 34944 0 FreeSans 448 0 0 0 io_wbs_datwr_1[12]
port 265 nsew signal tristate
flabel metal3 s 0 35504 800 35616 0 FreeSans 448 0 0 0 io_wbs_datwr_1[13]
port 266 nsew signal tristate
flabel metal3 s 0 36176 800 36288 0 FreeSans 448 0 0 0 io_wbs_datwr_1[14]
port 267 nsew signal tristate
flabel metal3 s 0 36848 800 36960 0 FreeSans 448 0 0 0 io_wbs_datwr_1[15]
port 268 nsew signal tristate
flabel metal3 s 0 37520 800 37632 0 FreeSans 448 0 0 0 io_wbs_datwr_1[16]
port 269 nsew signal tristate
flabel metal3 s 0 38192 800 38304 0 FreeSans 448 0 0 0 io_wbs_datwr_1[17]
port 270 nsew signal tristate
flabel metal3 s 0 38864 800 38976 0 FreeSans 448 0 0 0 io_wbs_datwr_1[18]
port 271 nsew signal tristate
flabel metal3 s 0 39536 800 39648 0 FreeSans 448 0 0 0 io_wbs_datwr_1[19]
port 272 nsew signal tristate
flabel metal3 s 0 27440 800 27552 0 FreeSans 448 0 0 0 io_wbs_datwr_1[1]
port 273 nsew signal tristate
flabel metal3 s 0 40208 800 40320 0 FreeSans 448 0 0 0 io_wbs_datwr_1[20]
port 274 nsew signal tristate
flabel metal3 s 0 40880 800 40992 0 FreeSans 448 0 0 0 io_wbs_datwr_1[21]
port 275 nsew signal tristate
flabel metal3 s 0 41552 800 41664 0 FreeSans 448 0 0 0 io_wbs_datwr_1[22]
port 276 nsew signal tristate
flabel metal3 s 0 42224 800 42336 0 FreeSans 448 0 0 0 io_wbs_datwr_1[23]
port 277 nsew signal tristate
flabel metal3 s 0 42896 800 43008 0 FreeSans 448 0 0 0 io_wbs_datwr_1[24]
port 278 nsew signal tristate
flabel metal3 s 0 43568 800 43680 0 FreeSans 448 0 0 0 io_wbs_datwr_1[25]
port 279 nsew signal tristate
flabel metal3 s 0 44240 800 44352 0 FreeSans 448 0 0 0 io_wbs_datwr_1[26]
port 280 nsew signal tristate
flabel metal3 s 0 44912 800 45024 0 FreeSans 448 0 0 0 io_wbs_datwr_1[27]
port 281 nsew signal tristate
flabel metal3 s 0 45584 800 45696 0 FreeSans 448 0 0 0 io_wbs_datwr_1[28]
port 282 nsew signal tristate
flabel metal3 s 0 46256 800 46368 0 FreeSans 448 0 0 0 io_wbs_datwr_1[29]
port 283 nsew signal tristate
flabel metal3 s 0 28112 800 28224 0 FreeSans 448 0 0 0 io_wbs_datwr_1[2]
port 284 nsew signal tristate
flabel metal3 s 0 46928 800 47040 0 FreeSans 448 0 0 0 io_wbs_datwr_1[30]
port 285 nsew signal tristate
flabel metal3 s 0 47600 800 47712 0 FreeSans 448 0 0 0 io_wbs_datwr_1[31]
port 286 nsew signal tristate
flabel metal3 s 0 28784 800 28896 0 FreeSans 448 0 0 0 io_wbs_datwr_1[3]
port 287 nsew signal tristate
flabel metal3 s 0 29456 800 29568 0 FreeSans 448 0 0 0 io_wbs_datwr_1[4]
port 288 nsew signal tristate
flabel metal3 s 0 30128 800 30240 0 FreeSans 448 0 0 0 io_wbs_datwr_1[5]
port 289 nsew signal tristate
flabel metal3 s 0 30800 800 30912 0 FreeSans 448 0 0 0 io_wbs_datwr_1[6]
port 290 nsew signal tristate
flabel metal3 s 0 31472 800 31584 0 FreeSans 448 0 0 0 io_wbs_datwr_1[7]
port 291 nsew signal tristate
flabel metal3 s 0 32144 800 32256 0 FreeSans 448 0 0 0 io_wbs_datwr_1[8]
port 292 nsew signal tristate
flabel metal3 s 0 32816 800 32928 0 FreeSans 448 0 0 0 io_wbs_datwr_1[9]
port 293 nsew signal tristate
flabel metal2 s 70448 0 70560 800 0 FreeSans 448 90 0 0 io_wbs_sel[0]
port 294 nsew signal input
flabel metal2 s 71120 0 71232 800 0 FreeSans 448 90 0 0 io_wbs_sel[1]
port 295 nsew signal input
flabel metal2 s 71792 0 71904 800 0 FreeSans 448 90 0 0 io_wbs_sel[2]
port 296 nsew signal input
flabel metal2 s 72464 0 72576 800 0 FreeSans 448 90 0 0 io_wbs_sel[3]
port 297 nsew signal input
flabel metal3 s 79200 70448 80000 70560 0 FreeSans 448 0 0 0 io_wbs_sel_0[0]
port 298 nsew signal tristate
flabel metal3 s 79200 71120 80000 71232 0 FreeSans 448 0 0 0 io_wbs_sel_0[1]
port 299 nsew signal tristate
flabel metal3 s 79200 71792 80000 71904 0 FreeSans 448 0 0 0 io_wbs_sel_0[2]
port 300 nsew signal tristate
flabel metal3 s 79200 72464 80000 72576 0 FreeSans 448 0 0 0 io_wbs_sel_0[3]
port 301 nsew signal tristate
flabel metal3 s 0 70448 800 70560 0 FreeSans 448 0 0 0 io_wbs_sel_1[0]
port 302 nsew signal tristate
flabel metal3 s 0 71120 800 71232 0 FreeSans 448 0 0 0 io_wbs_sel_1[1]
port 303 nsew signal tristate
flabel metal3 s 0 71792 800 71904 0 FreeSans 448 0 0 0 io_wbs_sel_1[2]
port 304 nsew signal tristate
flabel metal3 s 0 72464 800 72576 0 FreeSans 448 0 0 0 io_wbs_sel_1[3]
port 305 nsew signal tristate
flabel metal2 s 73136 0 73248 800 0 FreeSans 448 90 0 0 io_wbs_stb
port 306 nsew signal input
flabel metal3 s 79200 73136 80000 73248 0 FreeSans 448 0 0 0 io_wbs_stb_0
port 307 nsew signal tristate
flabel metal3 s 0 73136 800 73248 0 FreeSans 448 0 0 0 io_wbs_stb_1
port 308 nsew signal tristate
flabel metal2 s 69776 0 69888 800 0 FreeSans 448 90 0 0 io_wbs_we
port 309 nsew signal input
flabel metal3 s 79200 69776 80000 69888 0 FreeSans 448 0 0 0 io_wbs_we_0
port 310 nsew signal tristate
flabel metal3 s 0 69776 800 69888 0 FreeSans 448 0 0 0 io_wbs_we_1
port 311 nsew signal tristate
flabel metal4 s 4448 3076 4768 76892 0 FreeSans 1280 90 0 0 vdd
port 312 nsew power bidirectional
flabel metal4 s 35168 3076 35488 76892 0 FreeSans 1280 90 0 0 vdd
port 312 nsew power bidirectional
flabel metal4 s 65888 3076 66208 76892 0 FreeSans 1280 90 0 0 vdd
port 312 nsew power bidirectional
flabel metal4 s 19808 3076 20128 76892 0 FreeSans 1280 90 0 0 vss
port 313 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 76892 0 FreeSans 1280 90 0 0 vss
port 313 nsew ground bidirectional
rlabel metal1 39984 76048 39984 76048 0 vdd
rlabel metal1 39984 76832 39984 76832 0 vss
rlabel metal3 73304 50008 73304 50008 0 _000_
rlabel metal2 20888 17472 20888 17472 0 _001_
rlabel metal2 26264 17304 26264 17304 0 _002_
rlabel metal2 55384 17136 55384 17136 0 _003_
rlabel metal3 20776 16072 20776 16072 0 _004_
rlabel metal2 22904 16464 22904 16464 0 _005_
rlabel metal2 23296 16296 23296 16296 0 _006_
rlabel metal2 55048 15960 55048 15960 0 _007_
rlabel metal3 56000 51352 56000 51352 0 _008_
rlabel metal2 57232 52024 57232 52024 0 _009_
rlabel metal3 68544 64120 68544 64120 0 _010_
rlabel metal2 67928 48720 67928 48720 0 _011_
rlabel metal2 56280 18144 56280 18144 0 _012_
rlabel metal2 55888 51912 55888 51912 0 _013_
rlabel metal2 59416 60648 59416 60648 0 _014_
rlabel metal2 68152 66528 68152 66528 0 _015_
rlabel metal3 69216 48888 69216 48888 0 _016_
rlabel metal2 73416 50064 73416 50064 0 _017_
rlabel metal3 67704 48776 67704 48776 0 _018_
rlabel metal3 68992 49000 68992 49000 0 _019_
rlabel metal2 48552 48608 48552 48608 0 _020_
rlabel metal2 53704 51520 53704 51520 0 _021_
rlabel metal2 50456 50400 50456 50400 0 _022_
rlabel metal3 54432 55272 54432 55272 0 _023_
rlabel metal2 50904 50792 50904 50792 0 _024_
rlabel metal2 49560 47880 49560 47880 0 _025_
rlabel metal3 49112 48216 49112 48216 0 _026_
rlabel metal2 50344 48496 50344 48496 0 _027_
rlabel metal3 48608 49896 48608 49896 0 _028_
rlabel metal2 51184 49560 51184 49560 0 _029_
rlabel metal3 50120 50456 50120 50456 0 _030_
rlabel metal2 51408 50568 51408 50568 0 _031_
rlabel metal2 52136 51408 52136 51408 0 _032_
rlabel metal2 51968 51912 51968 51912 0 _033_
rlabel metal2 52360 52584 52360 52584 0 _034_
rlabel metal2 52584 51744 52584 51744 0 _035_
rlabel metal3 50344 51912 50344 51912 0 _036_
rlabel metal3 57064 52360 57064 52360 0 _037_
rlabel metal2 53816 51688 53816 51688 0 _038_
rlabel metal3 56504 52472 56504 52472 0 _039_
rlabel metal3 51856 52920 51856 52920 0 _040_
rlabel metal2 53536 52920 53536 52920 0 _041_
rlabel metal3 53816 53704 53816 53704 0 _042_
rlabel metal2 54712 54208 54712 54208 0 _043_
rlabel metal2 54488 55272 54488 55272 0 _044_
rlabel metal2 54264 54096 54264 54096 0 _045_
rlabel metal3 53592 54600 53592 54600 0 _046_
rlabel metal3 55664 54264 55664 54264 0 _047_
rlabel metal3 53144 55160 53144 55160 0 _048_
rlabel metal2 56616 54992 56616 54992 0 _049_
rlabel metal3 54432 56056 54432 56056 0 _050_
rlabel metal2 56336 55832 56336 55832 0 _051_
rlabel metal3 57288 56280 57288 56280 0 _052_
rlabel metal2 57344 54824 57344 54824 0 _053_
rlabel metal3 57680 55160 57680 55160 0 _054_
rlabel metal3 58576 56056 58576 56056 0 _055_
rlabel metal2 55272 57120 55272 57120 0 _056_
rlabel metal2 58072 57232 58072 57232 0 _057_
rlabel metal3 57120 57624 57120 57624 0 _058_
rlabel metal3 58856 57624 58856 57624 0 _059_
rlabel metal3 57736 58408 57736 58408 0 _060_
rlabel metal2 58576 58632 58576 58632 0 _061_
rlabel metal2 59864 59584 59864 59584 0 _062_
rlabel metal3 61712 60872 61712 60872 0 _063_
rlabel metal3 61712 60648 61712 60648 0 _064_
rlabel metal2 60312 59472 60312 59472 0 _065_
rlabel metal3 59192 59864 59192 59864 0 _066_
rlabel metal3 63560 59976 63560 59976 0 _067_
rlabel metal3 59304 60760 59304 60760 0 _068_
rlabel metal3 62944 60536 62944 60536 0 _069_
rlabel metal3 61432 60984 61432 60984 0 _070_
rlabel metal2 61992 61040 61992 61040 0 _071_
rlabel metal2 61544 62720 61544 62720 0 _072_
rlabel metal2 63280 61320 63280 61320 0 _073_
rlabel metal3 63168 63784 63168 63784 0 _074_
rlabel metal3 62048 62216 62048 62216 0 _075_
rlabel metal3 61880 62328 61880 62328 0 _076_
rlabel metal3 66304 62216 66304 62216 0 _077_
rlabel metal3 61432 62888 61432 62888 0 _078_
rlabel metal2 63896 63896 63896 63896 0 _079_
rlabel metal3 62384 64008 62384 64008 0 _080_
rlabel metal2 64288 63672 64288 63672 0 _081_
rlabel metal3 63616 64456 63616 64456 0 _082_
rlabel metal2 65128 64344 65128 64344 0 _083_
rlabel metal2 65912 66360 65912 66360 0 _084_
rlabel metal2 66080 64680 66080 64680 0 _085_
rlabel metal2 62104 65520 62104 65520 0 _086_
rlabel metal2 65072 65240 65072 65240 0 _087_
rlabel metal3 64624 66024 64624 66024 0 _088_
rlabel metal2 66528 66248 66528 66248 0 _089_
rlabel metal3 64736 67032 64736 67032 0 _090_
rlabel metal2 66640 66808 66640 66808 0 _091_
rlabel metal2 67928 66528 67928 66528 0 _092_
rlabel metal3 68880 66472 68880 66472 0 _093_
rlabel metal2 68264 65968 68264 65968 0 _094_
rlabel metal2 68712 65520 68712 65520 0 _095_
rlabel metal2 68376 67816 68376 67816 0 _096_
rlabel metal2 68768 67032 68768 67032 0 _097_
rlabel metal2 73976 72128 73976 72128 0 _098_
rlabel metal2 74088 72128 74088 72128 0 _099_
rlabel metal2 73864 2198 73864 2198 0 io_wbs_ack
rlabel metal3 77336 73920 77336 73920 0 io_wbs_ack_0
rlabel metal3 3248 73976 3248 73976 0 io_wbs_ack_1
rlabel metal2 4200 5264 4200 5264 0 io_wbs_adr[0]
rlabel metal2 11872 3416 11872 3416 0 io_wbs_adr[10]
rlabel metal2 12712 2590 12712 2590 0 io_wbs_adr[11]
rlabel metal2 13720 4368 13720 4368 0 io_wbs_adr[12]
rlabel metal2 14224 4424 14224 4424 0 io_wbs_adr[13]
rlabel metal2 14728 2086 14728 2086 0 io_wbs_adr[14]
rlabel metal3 16520 3416 16520 3416 0 io_wbs_adr[15]
rlabel metal2 16016 5992 16016 5992 0 io_wbs_adr[16]
rlabel metal2 17976 5712 17976 5712 0 io_wbs_adr[17]
rlabel metal2 17528 4200 17528 4200 0 io_wbs_adr[18]
rlabel metal2 18424 6552 18424 6552 0 io_wbs_adr[19]
rlabel metal2 5768 3360 5768 3360 0 io_wbs_adr[1]
rlabel metal2 18816 4200 18816 4200 0 io_wbs_adr[20]
rlabel metal2 20496 5992 20496 5992 0 io_wbs_adr[21]
rlabel metal2 19544 3976 19544 3976 0 io_wbs_adr[22]
rlabel metal3 21336 5096 21336 5096 0 io_wbs_adr[23]
rlabel metal2 21336 4032 21336 4032 0 io_wbs_adr[24]
rlabel metal2 22008 6440 22008 6440 0 io_wbs_adr[25]
rlabel metal2 22792 2926 22792 2926 0 io_wbs_adr[26]
rlabel metal3 22960 3528 22960 3528 0 io_wbs_adr[27]
rlabel metal2 23968 4984 23968 4984 0 io_wbs_adr[28]
rlabel metal2 24808 2590 24808 2590 0 io_wbs_adr[29]
rlabel metal2 6776 3416 6776 3416 0 io_wbs_adr[2]
rlabel metal2 25424 3416 25424 3416 0 io_wbs_adr[30]
rlabel metal3 26488 4200 26488 4200 0 io_wbs_adr[31]
rlabel metal2 7336 3374 7336 3374 0 io_wbs_adr[3]
rlabel metal2 8120 3752 8120 3752 0 io_wbs_adr[4]
rlabel metal2 8008 4032 8008 4032 0 io_wbs_adr[5]
rlabel metal2 9352 2086 9352 2086 0 io_wbs_adr[6]
rlabel metal2 10304 4984 10304 4984 0 io_wbs_adr[7]
rlabel metal2 10976 4424 10976 4424 0 io_wbs_adr[8]
rlabel metal3 11928 4984 11928 4984 0 io_wbs_adr[9]
rlabel metal2 77896 5544 77896 5544 0 io_wbs_adr_0[0]
rlabel metal2 76104 11760 76104 11760 0 io_wbs_adr_0[10]
rlabel metal2 76104 12488 76104 12488 0 io_wbs_adr_0[11]
rlabel metal2 76104 13216 76104 13216 0 io_wbs_adr_0[12]
rlabel metal2 76104 13944 76104 13944 0 io_wbs_adr_0[13]
rlabel metal2 76104 14672 76104 14672 0 io_wbs_adr_0[14]
rlabel metal3 77658 15400 77658 15400 0 io_wbs_adr_0[15]
rlabel metal2 77896 16464 77896 16464 0 io_wbs_adr_0[16]
rlabel metal2 76104 16464 76104 16464 0 io_wbs_adr_0[17]
rlabel metal2 76104 17192 76104 17192 0 io_wbs_adr_0[18]
rlabel metal2 76104 17920 76104 17920 0 io_wbs_adr_0[19]
rlabel metal3 77658 5992 77658 5992 0 io_wbs_adr_0[1]
rlabel metal2 76104 18592 76104 18592 0 io_wbs_adr_0[20]
rlabel metal2 76104 19376 76104 19376 0 io_wbs_adr_0[21]
rlabel metal3 77658 20104 77658 20104 0 io_wbs_adr_0[22]
rlabel metal2 77896 21112 77896 21112 0 io_wbs_adr_0[23]
rlabel metal2 76104 21168 76104 21168 0 io_wbs_adr_0[24]
rlabel metal2 76104 21896 76104 21896 0 io_wbs_adr_0[25]
rlabel metal2 76104 22624 76104 22624 0 io_wbs_adr_0[26]
rlabel metal2 76104 23352 76104 23352 0 io_wbs_adr_0[27]
rlabel metal2 76104 24080 76104 24080 0 io_wbs_adr_0[28]
rlabel metal3 77658 24808 77658 24808 0 io_wbs_adr_0[29]
rlabel metal2 77896 7056 77896 7056 0 io_wbs_adr_0[2]
rlabel metal2 77896 25816 77896 25816 0 io_wbs_adr_0[30]
rlabel metal2 76104 25872 76104 25872 0 io_wbs_adr_0[31]
rlabel metal2 76104 7000 76104 7000 0 io_wbs_adr_0[3]
rlabel metal2 76104 7784 76104 7784 0 io_wbs_adr_0[4]
rlabel metal3 76328 8344 76328 8344 0 io_wbs_adr_0[5]
rlabel metal2 76104 9240 76104 9240 0 io_wbs_adr_0[6]
rlabel metal2 76104 9968 76104 9968 0 io_wbs_adr_0[7]
rlabel metal3 77658 10696 77658 10696 0 io_wbs_adr_0[8]
rlabel metal2 77896 11704 77896 11704 0 io_wbs_adr_0[9]
rlabel metal3 1358 5320 1358 5320 0 io_wbs_adr_1[0]
rlabel metal3 1358 12040 1358 12040 0 io_wbs_adr_1[10]
rlabel metal3 1358 12712 1358 12712 0 io_wbs_adr_1[11]
rlabel metal3 1358 13384 1358 13384 0 io_wbs_adr_1[12]
rlabel metal3 1358 14056 1358 14056 0 io_wbs_adr_1[13]
rlabel metal3 1358 14728 1358 14728 0 io_wbs_adr_1[14]
rlabel metal3 1358 15400 1358 15400 0 io_wbs_adr_1[15]
rlabel metal3 2254 16072 2254 16072 0 io_wbs_adr_1[16]
rlabel metal3 1358 16744 1358 16744 0 io_wbs_adr_1[17]
rlabel metal3 1358 17416 1358 17416 0 io_wbs_adr_1[18]
rlabel metal3 1358 18088 1358 18088 0 io_wbs_adr_1[19]
rlabel metal3 1358 5992 1358 5992 0 io_wbs_adr_1[1]
rlabel metal3 1358 18760 1358 18760 0 io_wbs_adr_1[20]
rlabel metal3 1358 19432 1358 19432 0 io_wbs_adr_1[21]
rlabel metal3 1358 20104 1358 20104 0 io_wbs_adr_1[22]
rlabel metal3 2254 20776 2254 20776 0 io_wbs_adr_1[23]
rlabel metal3 1358 21448 1358 21448 0 io_wbs_adr_1[24]
rlabel metal3 1358 22120 1358 22120 0 io_wbs_adr_1[25]
rlabel metal3 1358 22792 1358 22792 0 io_wbs_adr_1[26]
rlabel metal3 1358 23464 1358 23464 0 io_wbs_adr_1[27]
rlabel metal3 1358 24136 1358 24136 0 io_wbs_adr_1[28]
rlabel metal3 1358 24808 1358 24808 0 io_wbs_adr_1[29]
rlabel metal3 2254 6664 2254 6664 0 io_wbs_adr_1[2]
rlabel metal3 2254 25480 2254 25480 0 io_wbs_adr_1[30]
rlabel metal3 1358 26152 1358 26152 0 io_wbs_adr_1[31]
rlabel metal3 1358 7336 1358 7336 0 io_wbs_adr_1[3]
rlabel metal3 1358 8008 1358 8008 0 io_wbs_adr_1[4]
rlabel metal3 1358 8680 1358 8680 0 io_wbs_adr_1[5]
rlabel metal3 1358 9352 1358 9352 0 io_wbs_adr_1[6]
rlabel metal3 1358 10024 1358 10024 0 io_wbs_adr_1[7]
rlabel metal3 1358 10696 1358 10696 0 io_wbs_adr_1[8]
rlabel metal3 2254 11368 2254 11368 0 io_wbs_adr_1[9]
rlabel metal3 74816 3416 74816 3416 0 io_wbs_cyc
rlabel metal2 75600 75768 75600 75768 0 io_wbs_cyc_0
rlabel metal3 1414 74536 1414 74536 0 io_wbs_cyc_1
rlabel metal2 48328 2926 48328 2926 0 io_wbs_datrd[0]
rlabel metal2 55048 2982 55048 2982 0 io_wbs_datrd[10]
rlabel metal2 55720 1414 55720 1414 0 io_wbs_datrd[11]
rlabel metal2 56392 2086 56392 2086 0 io_wbs_datrd[12]
rlabel metal2 57064 2926 57064 2926 0 io_wbs_datrd[13]
rlabel metal2 57736 2478 57736 2478 0 io_wbs_datrd[14]
rlabel metal2 58408 2142 58408 2142 0 io_wbs_datrd[15]
rlabel metal2 59080 854 59080 854 0 io_wbs_datrd[16]
rlabel metal2 59752 2254 59752 2254 0 io_wbs_datrd[17]
rlabel metal2 60424 2198 60424 2198 0 io_wbs_datrd[18]
rlabel metal2 61096 1638 61096 1638 0 io_wbs_datrd[19]
rlabel metal2 49000 3262 49000 3262 0 io_wbs_datrd[1]
rlabel metal2 61768 1414 61768 1414 0 io_wbs_datrd[20]
rlabel metal2 62440 1246 62440 1246 0 io_wbs_datrd[21]
rlabel metal2 63112 854 63112 854 0 io_wbs_datrd[22]
rlabel metal2 63784 2422 63784 2422 0 io_wbs_datrd[23]
rlabel metal2 64456 2086 64456 2086 0 io_wbs_datrd[24]
rlabel metal2 65128 2870 65128 2870 0 io_wbs_datrd[25]
rlabel metal2 65800 2478 65800 2478 0 io_wbs_datrd[26]
rlabel metal2 66472 1694 66472 1694 0 io_wbs_datrd[27]
rlabel metal2 67256 5320 67256 5320 0 io_wbs_datrd[28]
rlabel metal2 67816 854 67816 854 0 io_wbs_datrd[29]
rlabel metal2 49672 2478 49672 2478 0 io_wbs_datrd[2]
rlabel metal2 68488 2926 68488 2926 0 io_wbs_datrd[30]
rlabel metal2 69160 2254 69160 2254 0 io_wbs_datrd[31]
rlabel metal2 50344 2198 50344 2198 0 io_wbs_datrd[3]
rlabel metal2 51016 2982 51016 2982 0 io_wbs_datrd[4]
rlabel metal2 51688 2142 51688 2142 0 io_wbs_datrd[5]
rlabel metal2 52360 2086 52360 2086 0 io_wbs_datrd[6]
rlabel metal2 53032 2870 53032 2870 0 io_wbs_datrd[7]
rlabel metal2 53704 2478 53704 2478 0 io_wbs_datrd[8]
rlabel metal2 54376 2198 54376 2198 0 io_wbs_datrd[9]
rlabel metal2 77336 48552 77336 48552 0 io_wbs_datrd_0[0]
rlabel metal3 79128 55384 79128 55384 0 io_wbs_datrd_0[10]
rlabel metal2 76944 57512 76944 57512 0 io_wbs_datrd_0[11]
rlabel metal2 77336 57848 77336 57848 0 io_wbs_datrd_0[12]
rlabel metal2 76832 59080 76832 59080 0 io_wbs_datrd_0[13]
rlabel metal2 77392 59752 77392 59752 0 io_wbs_datrd_0[14]
rlabel metal2 76888 60312 76888 60312 0 io_wbs_datrd_0[15]
rlabel metal2 77280 61320 77280 61320 0 io_wbs_datrd_0[16]
rlabel metal2 74312 59808 74312 59808 0 io_wbs_datrd_0[17]
rlabel metal2 76944 62216 76944 62216 0 io_wbs_datrd_0[18]
rlabel metal2 77336 62552 77336 62552 0 io_wbs_datrd_0[19]
rlabel metal2 76888 49336 76888 49336 0 io_wbs_datrd_0[1]
rlabel metal2 76888 63560 76888 63560 0 io_wbs_datrd_0[20]
rlabel metal2 77392 64456 77392 64456 0 io_wbs_datrd_0[21]
rlabel metal2 76832 65352 76832 65352 0 io_wbs_datrd_0[22]
rlabel metal2 77336 65800 77336 65800 0 io_wbs_datrd_0[23]
rlabel metal2 74312 64512 74312 64512 0 io_wbs_datrd_0[24]
rlabel metal2 76888 66248 76888 66248 0 io_wbs_datrd_0[25]
rlabel metal3 76832 67704 76832 67704 0 io_wbs_datrd_0[26]
rlabel metal2 76944 68488 76944 68488 0 io_wbs_datrd_0[27]
rlabel metal2 77392 69160 77392 69160 0 io_wbs_datrd_0[28]
rlabel metal2 76832 70056 76832 70056 0 io_wbs_datrd_0[29]
rlabel metal2 77336 50064 77336 50064 0 io_wbs_datrd_0[2]
rlabel metal2 77336 70672 77336 70672 0 io_wbs_datrd_0[30]
rlabel metal2 74312 69216 74312 69216 0 io_wbs_datrd_0[31]
rlabel metal2 76888 50792 76888 50792 0 io_wbs_datrd_0[3]
rlabel metal2 77336 51576 77336 51576 0 io_wbs_datrd_0[4]
rlabel metal2 76888 52248 76888 52248 0 io_wbs_datrd_0[5]
rlabel metal2 77336 52920 77336 52920 0 io_wbs_datrd_0[6]
rlabel metal2 76888 53816 76888 53816 0 io_wbs_datrd_0[7]
rlabel metal2 77336 54432 77336 54432 0 io_wbs_datrd_0[8]
rlabel metal3 78106 54376 78106 54376 0 io_wbs_datrd_0[9]
rlabel metal2 1960 48608 1960 48608 0 io_wbs_datrd_1[0]
rlabel metal3 910 55048 910 55048 0 io_wbs_datrd_1[10]
rlabel metal2 1960 56728 1960 56728 0 io_wbs_datrd_1[11]
rlabel metal2 2072 57344 2072 57344 0 io_wbs_datrd_1[12]
rlabel metal2 1904 59304 1904 59304 0 io_wbs_datrd_1[13]
rlabel metal2 2296 58800 2296 58800 0 io_wbs_datrd_1[14]
rlabel metal2 2184 59640 2184 59640 0 io_wbs_datrd_1[15]
rlabel metal2 3976 59192 3976 59192 0 io_wbs_datrd_1[16]
rlabel metal2 2072 60592 2072 60592 0 io_wbs_datrd_1[17]
rlabel metal2 1904 62440 1904 62440 0 io_wbs_datrd_1[18]
rlabel metal2 2184 62048 2184 62048 0 io_wbs_datrd_1[19]
rlabel metal2 2072 49448 2072 49448 0 io_wbs_datrd_1[1]
rlabel metal2 2072 62888 2072 62888 0 io_wbs_datrd_1[20]
rlabel metal2 1960 63616 1960 63616 0 io_wbs_datrd_1[21]
rlabel metal2 1904 65576 1904 65576 0 io_wbs_datrd_1[22]
rlabel metal2 3976 63896 3976 63896 0 io_wbs_datrd_1[23]
rlabel metal2 2072 65296 2072 65296 0 io_wbs_datrd_1[24]
rlabel metal2 2184 66136 2184 66136 0 io_wbs_datrd_1[25]
rlabel metal3 3248 67704 3248 67704 0 io_wbs_datrd_1[26]
rlabel metal3 3024 68712 3024 68712 0 io_wbs_datrd_1[27]
rlabel metal3 3248 69272 3248 69272 0 io_wbs_datrd_1[28]
rlabel metal2 1904 70280 1904 70280 0 io_wbs_datrd_1[29]
rlabel metal2 1960 50120 1960 50120 0 io_wbs_datrd_1[2]
rlabel metal2 3976 68600 3976 68600 0 io_wbs_datrd_1[30]
rlabel metal2 2184 70000 2184 70000 0 io_wbs_datrd_1[31]
rlabel metal2 2184 50960 2184 50960 0 io_wbs_datrd_1[3]
rlabel metal2 2072 51520 2072 51520 0 io_wbs_datrd_1[4]
rlabel metal2 1960 52360 1960 52360 0 io_wbs_datrd_1[5]
rlabel metal2 2072 52976 2072 52976 0 io_wbs_datrd_1[6]
rlabel metal2 2184 53816 2184 53816 0 io_wbs_datrd_1[7]
rlabel metal2 2072 54488 2072 54488 0 io_wbs_datrd_1[8]
rlabel metal3 1302 54376 1302 54376 0 io_wbs_datrd_1[9]
rlabel metal2 26600 5208 26600 5208 0 io_wbs_datwr[0]
rlabel metal2 33208 3360 33208 3360 0 io_wbs_datwr[10]
rlabel metal2 34384 4200 34384 4200 0 io_wbs_datwr[11]
rlabel metal2 34776 5768 34776 5768 0 io_wbs_datwr[12]
rlabel metal2 36344 5040 36344 5040 0 io_wbs_datwr[13]
rlabel metal3 36624 3528 36624 3528 0 io_wbs_datwr[14]
rlabel metal3 36064 3416 36064 3416 0 io_wbs_datwr[15]
rlabel metal2 38136 3920 38136 3920 0 io_wbs_datwr[16]
rlabel metal2 38024 4816 38024 4816 0 io_wbs_datwr[17]
rlabel metal3 39032 3640 39032 3640 0 io_wbs_datwr[18]
rlabel metal2 39704 3416 39704 3416 0 io_wbs_datwr[19]
rlabel metal3 28224 5992 28224 5992 0 io_wbs_datwr[1]
rlabel metal2 40264 3262 40264 3262 0 io_wbs_datwr[20]
rlabel metal2 41272 3024 41272 3024 0 io_wbs_datwr[21]
rlabel metal3 42224 3416 42224 3416 0 io_wbs_datwr[22]
rlabel metal2 42448 4984 42448 4984 0 io_wbs_datwr[23]
rlabel metal2 44296 4032 44296 4032 0 io_wbs_datwr[24]
rlabel metal2 45976 3528 45976 3528 0 io_wbs_datwr[25]
rlabel metal2 45752 4312 45752 4312 0 io_wbs_datwr[26]
rlabel metal2 44856 4200 44856 4200 0 io_wbs_datwr[27]
rlabel metal3 46928 3416 46928 3416 0 io_wbs_datwr[28]
rlabel metal3 46928 4200 46928 4200 0 io_wbs_datwr[29]
rlabel metal2 28280 4984 28280 4984 0 io_wbs_datwr[2]
rlabel metal2 46760 4872 46760 4872 0 io_wbs_datwr[30]
rlabel metal2 48776 4144 48776 4144 0 io_wbs_datwr[31]
rlabel metal2 29176 2968 29176 2968 0 io_wbs_datwr[3]
rlabel metal3 30016 5992 30016 5992 0 io_wbs_datwr[4]
rlabel metal2 29736 2800 29736 2800 0 io_wbs_datwr[5]
rlabel metal2 30856 2926 30856 2926 0 io_wbs_datwr[6]
rlabel metal2 31528 910 31528 910 0 io_wbs_datwr[7]
rlabel metal2 32312 4032 32312 4032 0 io_wbs_datwr[8]
rlabel metal2 32816 4424 32816 4424 0 io_wbs_datwr[9]
rlabel metal2 76104 26600 76104 26600 0 io_wbs_datwr_0[0]
rlabel metal2 76104 33488 76104 33488 0 io_wbs_datwr_0[10]
rlabel metal3 77658 34216 77658 34216 0 io_wbs_datwr_0[11]
rlabel metal2 77896 35224 77896 35224 0 io_wbs_datwr_0[12]
rlabel metal2 76104 35280 76104 35280 0 io_wbs_datwr_0[13]
rlabel metal2 76104 36008 76104 36008 0 io_wbs_datwr_0[14]
rlabel metal2 76104 36736 76104 36736 0 io_wbs_datwr_0[15]
rlabel metal2 76104 37464 76104 37464 0 io_wbs_datwr_0[16]
rlabel metal2 76104 38192 76104 38192 0 io_wbs_datwr_0[17]
rlabel metal3 77658 38920 77658 38920 0 io_wbs_datwr_0[18]
rlabel metal3 77658 39592 77658 39592 0 io_wbs_datwr_0[19]
rlabel metal2 76104 27328 76104 27328 0 io_wbs_datwr_0[1]
rlabel metal3 76104 40320 76104 40320 0 io_wbs_datwr_0[20]
rlabel metal2 76104 40992 76104 40992 0 io_wbs_datwr_0[21]
rlabel metal2 76104 41720 76104 41720 0 io_wbs_datwr_0[22]
rlabel metal2 76104 42448 76104 42448 0 io_wbs_datwr_0[23]
rlabel metal2 76104 43176 76104 43176 0 io_wbs_datwr_0[24]
rlabel metal2 76104 43960 76104 43960 0 io_wbs_datwr_0[25]
rlabel metal2 75992 44632 75992 44632 0 io_wbs_datwr_0[26]
rlabel metal2 76104 45360 76104 45360 0 io_wbs_datwr_0[27]
rlabel metal2 75992 46088 75992 46088 0 io_wbs_datwr_0[28]
rlabel metal2 76104 46816 76104 46816 0 io_wbs_datwr_0[29]
rlabel metal2 76104 28056 76104 28056 0 io_wbs_datwr_0[2]
rlabel metal2 75992 47600 75992 47600 0 io_wbs_datwr_0[30]
rlabel metal2 77896 47880 77896 47880 0 io_wbs_datwr_0[31]
rlabel metal2 76104 28784 76104 28784 0 io_wbs_datwr_0[3]
rlabel metal3 77658 29512 77658 29512 0 io_wbs_datwr_0[4]
rlabel metal2 77896 30576 77896 30576 0 io_wbs_datwr_0[5]
rlabel metal2 76104 30520 76104 30520 0 io_wbs_datwr_0[6]
rlabel metal2 76104 31304 76104 31304 0 io_wbs_datwr_0[7]
rlabel metal3 76328 31864 76328 31864 0 io_wbs_datwr_0[8]
rlabel metal2 76104 32760 76104 32760 0 io_wbs_datwr_0[9]
rlabel metal3 1358 26824 1358 26824 0 io_wbs_datwr_1[0]
rlabel metal3 1358 33544 1358 33544 0 io_wbs_datwr_1[10]
rlabel metal3 1358 34216 1358 34216 0 io_wbs_datwr_1[11]
rlabel metal3 2254 34888 2254 34888 0 io_wbs_datwr_1[12]
rlabel metal3 1358 35560 1358 35560 0 io_wbs_datwr_1[13]
rlabel metal3 1358 36232 1358 36232 0 io_wbs_datwr_1[14]
rlabel metal3 1358 36904 1358 36904 0 io_wbs_datwr_1[15]
rlabel metal3 1358 37576 1358 37576 0 io_wbs_datwr_1[16]
rlabel metal3 1358 38248 1358 38248 0 io_wbs_datwr_1[17]
rlabel metal3 1358 38920 1358 38920 0 io_wbs_datwr_1[18]
rlabel metal3 1358 39592 1358 39592 0 io_wbs_datwr_1[19]
rlabel metal3 1358 27496 1358 27496 0 io_wbs_datwr_1[1]
rlabel metal3 1358 40264 1358 40264 0 io_wbs_datwr_1[20]
rlabel metal3 1358 40936 1358 40936 0 io_wbs_datwr_1[21]
rlabel metal3 1358 41608 1358 41608 0 io_wbs_datwr_1[22]
rlabel metal3 1358 42280 1358 42280 0 io_wbs_datwr_1[23]
rlabel metal3 1358 42952 1358 42952 0 io_wbs_datwr_1[24]
rlabel metal3 1358 43624 1358 43624 0 io_wbs_datwr_1[25]
rlabel metal3 1414 44296 1414 44296 0 io_wbs_datwr_1[26]
rlabel metal3 1358 44968 1358 44968 0 io_wbs_datwr_1[27]
rlabel metal3 1414 45640 1414 45640 0 io_wbs_datwr_1[28]
rlabel metal3 1358 46312 1358 46312 0 io_wbs_datwr_1[29]
rlabel metal3 1358 28168 1358 28168 0 io_wbs_datwr_1[2]
rlabel metal3 1414 46984 1414 46984 0 io_wbs_datwr_1[30]
rlabel metal3 2254 47656 2254 47656 0 io_wbs_datwr_1[31]
rlabel metal3 1358 28840 1358 28840 0 io_wbs_datwr_1[3]
rlabel metal3 1358 29512 1358 29512 0 io_wbs_datwr_1[4]
rlabel metal3 2254 30184 2254 30184 0 io_wbs_datwr_1[5]
rlabel metal3 1358 30856 1358 30856 0 io_wbs_datwr_1[6]
rlabel metal3 1358 31528 1358 31528 0 io_wbs_datwr_1[7]
rlabel metal3 1358 32200 1358 32200 0 io_wbs_datwr_1[8]
rlabel metal3 1358 32872 1358 32872 0 io_wbs_datwr_1[9]
rlabel metal2 70392 4200 70392 4200 0 io_wbs_sel[0]
rlabel metal3 72296 3416 72296 3416 0 io_wbs_sel[1]
rlabel metal2 71736 5096 71736 5096 0 io_wbs_sel[2]
rlabel metal3 73472 4424 73472 4424 0 io_wbs_sel[3]
rlabel metal2 76104 71512 76104 71512 0 io_wbs_sel_0[0]
rlabel metal2 77896 71400 77896 71400 0 io_wbs_sel_0[1]
rlabel metal2 75992 72520 75992 72520 0 io_wbs_sel_0[2]
rlabel metal2 77896 72856 77896 72856 0 io_wbs_sel_0[3]
rlabel metal3 1302 70504 1302 70504 0 io_wbs_sel_1[0]
rlabel metal3 2254 71176 2254 71176 0 io_wbs_sel_1[1]
rlabel metal3 1414 71848 1414 71848 0 io_wbs_sel_1[2]
rlabel metal3 2254 72520 2254 72520 0 io_wbs_sel_1[3]
rlabel metal2 73864 5712 73864 5712 0 io_wbs_stb
rlabel metal2 75656 74368 75656 74368 0 io_wbs_stb_0
rlabel metal3 1358 73192 1358 73192 0 io_wbs_stb_1
rlabel metal2 69720 3416 69720 3416 0 io_wbs_we
rlabel metal2 75600 71624 75600 71624 0 io_wbs_we_0
rlabel metal3 1414 69832 1414 69832 0 io_wbs_we_1
rlabel metal2 74144 50680 74144 50680 0 net1
rlabel metal3 16912 5768 16912 5768 0 net10
rlabel metal2 27104 25368 27104 25368 0 net100
rlabel metal2 32200 6020 32200 6020 0 net101
rlabel metal2 34552 6804 34552 6804 0 net102
rlabel metal2 36288 20160 36288 20160 0 net103
rlabel metal2 35168 5208 35168 5208 0 net104
rlabel metal2 36624 4200 36624 4200 0 net105
rlabel metal2 36400 3640 36400 3640 0 net106
rlabel metal2 37464 4200 37464 4200 0 net107
rlabel metal3 39312 5208 39312 5208 0 net108
rlabel metal2 39536 37800 39536 37800 0 net109
rlabel metal2 16296 7588 16296 7588 0 net11
rlabel metal2 39144 3640 39144 3640 0 net110
rlabel metal2 27328 5768 27328 5768 0 net111
rlabel metal2 40432 38696 40432 38696 0 net112
rlabel metal3 42224 4984 42224 4984 0 net113
rlabel metal3 42112 40600 42112 40600 0 net114
rlabel metal3 43344 5208 43344 5208 0 net115
rlabel metal2 43568 20160 43568 20160 0 net116
rlabel metal3 44632 43512 44632 43512 0 net117
rlabel metal3 44352 44184 44352 44184 0 net118
rlabel metal2 46816 44072 46816 44072 0 net119
rlabel metal3 16968 5208 16968 5208 0 net12
rlabel metal3 48384 3640 48384 3640 0 net120
rlabel metal3 48272 5208 48272 5208 0 net121
rlabel metal2 27104 27720 27104 27720 0 net122
rlabel metal2 48328 46536 48328 46536 0 net123
rlabel metal3 48496 47320 48496 47320 0 net124
rlabel metal2 27776 28616 27776 28616 0 net125
rlabel metal3 29680 29400 29680 29400 0 net126
rlabel metal2 28560 3640 28560 3640 0 net127
rlabel metal2 31024 29400 31024 29400 0 net128
rlabel metal2 31640 7084 31640 7084 0 net129
rlabel metal2 19544 7588 19544 7588 0 net13
rlabel metal2 31192 30968 31192 30968 0 net130
rlabel metal2 31640 29512 31640 29512 0 net131
rlabel metal3 71456 4200 71456 4200 0 net132
rlabel metal2 72464 70728 72464 70728 0 net133
rlabel metal3 73080 70728 73080 70728 0 net134
rlabel metal2 73304 4200 73304 4200 0 net135
rlabel metal2 73920 5208 73920 5208 0 net136
rlabel metal3 70616 3640 70616 3640 0 net137
rlabel metal2 75656 3696 75656 3696 0 net138
rlabel metal2 76552 4984 76552 4984 0 net139
rlabel metal2 4984 5488 4984 5488 0 net14
rlabel metal2 74984 11312 74984 11312 0 net140
rlabel metal2 74984 12208 74984 12208 0 net141
rlabel metal2 74480 13048 74480 13048 0 net142
rlabel metal2 74984 13776 74984 13776 0 net143
rlabel metal2 74984 14392 74984 14392 0 net144
rlabel metal2 74984 15344 74984 15344 0 net145
rlabel metal2 76776 16352 76776 16352 0 net146
rlabel metal3 74760 16072 74760 16072 0 net147
rlabel metal2 74984 16912 74984 16912 0 net148
rlabel metal2 74984 17584 74984 17584 0 net149
rlabel metal2 20552 17360 20552 17360 0 net15
rlabel metal2 6776 4760 6776 4760 0 net150
rlabel metal2 21112 18480 21112 18480 0 net151
rlabel metal2 74984 19152 74984 19152 0 net152
rlabel metal2 74480 19880 74480 19880 0 net153
rlabel metal2 77224 20384 77224 20384 0 net154
rlabel metal2 74984 20664 74984 20664 0 net155
rlabel metal2 74984 21616 74984 21616 0 net156
rlabel metal2 74984 22232 74984 22232 0 net157
rlabel metal2 74984 23184 74984 23184 0 net158
rlabel metal2 74984 23800 74984 23800 0 net159
rlabel metal2 21616 18648 21616 18648 0 net16
rlabel metal2 24920 24752 24920 24752 0 net160
rlabel metal2 7336 6608 7336 6608 0 net161
rlabel metal2 77224 25088 77224 25088 0 net162
rlabel metal2 74984 25368 74984 25368 0 net163
rlabel metal2 8232 6272 8232 6272 0 net164
rlabel metal2 74984 7504 74984 7504 0 net165
rlabel metal2 74984 8120 74984 8120 0 net166
rlabel metal2 74984 9072 74984 9072 0 net167
rlabel metal2 74984 9688 74984 9688 0 net168
rlabel metal2 74984 10640 74984 10640 0 net169
rlabel metal2 20216 17472 20216 17472 0 net17
rlabel metal2 76776 11648 76776 11648 0 net170
rlabel metal3 3864 4536 3864 4536 0 net171
rlabel metal2 3080 11424 3080 11424 0 net172
rlabel metal2 3080 12208 3080 12208 0 net173
rlabel metal2 3080 12824 3080 12824 0 net174
rlabel metal2 3080 13664 3080 13664 0 net175
rlabel metal2 3080 14392 3080 14392 0 net176
rlabel metal2 3080 15232 3080 15232 0 net177
rlabel metal3 5152 16856 5152 16856 0 net178
rlabel metal2 3080 15960 3080 15960 0 net179
rlabel metal2 21000 7084 21000 7084 0 net18
rlabel metal2 3080 16912 3080 16912 0 net180
rlabel metal2 3640 17360 3640 17360 0 net181
rlabel metal2 3080 5936 3080 5936 0 net182
rlabel metal2 3080 18368 3080 18368 0 net183
rlabel metal2 3640 18928 3640 18928 0 net184
rlabel metal2 3080 19936 3080 19936 0 net185
rlabel metal2 4872 21504 4872 21504 0 net186
rlabel metal2 3080 20720 3080 20720 0 net187
rlabel metal2 2968 21224 2968 21224 0 net188
rlabel metal2 3080 22232 3080 22232 0 net189
rlabel metal3 21448 20776 21448 20776 0 net19
rlabel metal2 3080 23072 3080 23072 0 net190
rlabel metal2 3080 23800 3080 23800 0 net191
rlabel metal2 3640 24528 3640 24528 0 net192
rlabel metal3 5488 6552 5488 6552 0 net193
rlabel metal2 4872 26208 4872 26208 0 net194
rlabel metal2 3080 25424 3080 25424 0 net195
rlabel metal2 3080 6720 3080 6720 0 net196
rlabel metal2 3080 7504 3080 7504 0 net197
rlabel metal3 5600 8120 5600 8120 0 net198
rlabel metal2 3080 9072 3080 9072 0 net199
rlabel metal2 3360 74200 3360 74200 0 net2
rlabel metal3 22624 21560 22624 21560 0 net20
rlabel metal2 3080 9744 3080 9744 0 net200
rlabel metal2 3080 10640 3080 10640 0 net201
rlabel metal2 4872 11704 4872 11704 0 net202
rlabel metal3 74368 75096 74368 75096 0 net203
rlabel metal2 3528 74592 3528 74592 0 net204
rlabel metal2 51688 5544 51688 5544 0 net205
rlabel metal2 55160 6104 55160 6104 0 net206
rlabel metal2 55272 55048 55272 55048 0 net207
rlabel metal2 58184 6160 58184 6160 0 net208
rlabel metal2 58688 6104 58688 6104 0 net209
rlabel metal2 24304 22120 24304 22120 0 net21
rlabel metal2 59640 6216 59640 6216 0 net210
rlabel metal2 60312 6384 60312 6384 0 net211
rlabel metal2 59192 6272 59192 6272 0 net212
rlabel metal2 61544 6160 61544 6160 0 net213
rlabel metal2 62104 6216 62104 6216 0 net214
rlabel metal2 61320 5096 61320 5096 0 net215
rlabel metal3 50288 5880 50288 5880 0 net216
rlabel metal3 63560 4312 63560 4312 0 net217
rlabel metal2 64232 6160 64232 6160 0 net218
rlabel metal2 64960 5096 64960 5096 0 net219
rlabel metal2 23744 23128 23744 23128 0 net22
rlabel metal2 65800 6216 65800 6216 0 net220
rlabel metal2 67480 3976 67480 3976 0 net221
rlabel metal2 66360 6160 66360 6160 0 net222
rlabel metal3 68600 4312 68600 4312 0 net223
rlabel metal2 66752 6552 66752 6552 0 net224
rlabel metal2 67368 6048 67368 6048 0 net225
rlabel metal2 69384 5320 69384 5320 0 net226
rlabel metal3 50736 4312 50736 4312 0 net227
rlabel metal3 69496 5880 69496 5880 0 net228
rlabel metal3 68208 6664 68208 6664 0 net229
rlabel metal2 24360 22960 24360 22960 0 net23
rlabel metal2 52136 3696 52136 3696 0 net230
rlabel metal2 51240 3640 51240 3640 0 net231
rlabel metal2 53032 6160 53032 6160 0 net232
rlabel metal2 54264 6328 54264 6328 0 net233
rlabel metal2 55384 6216 55384 6216 0 net234
rlabel metal2 53032 29624 53032 29624 0 net235
rlabel metal2 54376 53480 54376 53480 0 net236
rlabel metal2 74984 26320 74984 26320 0 net237
rlabel metal2 74984 33208 74984 33208 0 net238
rlabel metal2 74984 34160 74984 34160 0 net239
rlabel metal2 23408 4200 23408 4200 0 net24
rlabel metal2 76776 35168 76776 35168 0 net240
rlabel metal2 74984 34832 74984 34832 0 net241
rlabel metal2 74984 35728 74984 35728 0 net242
rlabel metal2 74984 36344 74984 36344 0 net243
rlabel metal2 74984 37296 74984 37296 0 net244
rlabel metal2 74984 37912 74984 37912 0 net245
rlabel metal2 74984 38864 74984 38864 0 net246
rlabel metal2 74984 39480 74984 39480 0 net247
rlabel metal2 74536 26880 74536 26880 0 net248
rlabel metal2 74536 39984 74536 39984 0 net249
rlabel metal3 6048 6664 6048 6664 0 net25
rlabel metal2 74424 40712 74424 40712 0 net250
rlabel metal2 74536 41384 74536 41384 0 net251
rlabel metal2 74424 42280 74424 42280 0 net252
rlabel metal2 74536 42952 74536 42952 0 net253
rlabel metal2 74424 43904 74424 43904 0 net254
rlabel metal2 74536 44520 74536 44520 0 net255
rlabel metal2 45640 45416 45640 45416 0 net256
rlabel metal2 74536 45920 74536 45920 0 net257
rlabel metal2 74368 47208 74368 47208 0 net258
rlabel metal2 74984 27888 74984 27888 0 net259
rlabel metal2 26096 23688 26096 23688 0 net26
rlabel metal2 74536 47488 74536 47488 0 net260
rlabel metal2 76776 47712 76776 47712 0 net261
rlabel metal2 74536 28504 74536 28504 0 net262
rlabel metal2 74984 29456 74984 29456 0 net263
rlabel metal2 76776 30464 76776 30464 0 net264
rlabel metal2 74984 30128 74984 30128 0 net265
rlabel metal2 74984 31024 74984 31024 0 net266
rlabel metal2 74984 31640 74984 31640 0 net267
rlabel metal2 74984 32592 74984 32592 0 net268
rlabel metal2 2968 25760 2968 25760 0 net269
rlabel metal2 26544 25480 26544 25480 0 net27
rlabel metal2 3080 33264 3080 33264 0 net270
rlabel metal2 3080 34048 3080 34048 0 net271
rlabel metal2 4872 35616 4872 35616 0 net272
rlabel metal2 3080 34776 3080 34776 0 net273
rlabel metal2 3080 35728 3080 35728 0 net274
rlabel metal2 3080 36344 3080 36344 0 net275
rlabel metal2 3640 37072 3640 37072 0 net276
rlabel metal2 3080 37912 3080 37912 0 net277
rlabel metal3 3360 38808 3360 38808 0 net278
rlabel metal2 3080 39536 3080 39536 0 net279
rlabel metal2 7896 6720 7896 6720 0 net28
rlabel metal3 3360 27048 3360 27048 0 net280
rlabel metal3 3360 40376 3360 40376 0 net281
rlabel metal2 3080 41048 3080 41048 0 net282
rlabel metal2 3080 41888 3080 41888 0 net283
rlabel metal2 3080 42672 3080 42672 0 net284
rlabel metal2 3080 43456 3080 43456 0 net285
rlabel metal2 3080 44184 3080 44184 0 net286
rlabel metal2 3080 45024 3080 45024 0 net287
rlabel metal2 3528 45472 3528 45472 0 net288
rlabel metal2 3640 45864 3640 45864 0 net289
rlabel metal2 7672 6328 7672 6328 0 net29
rlabel metal2 3640 47208 3640 47208 0 net290
rlabel metal2 3080 27776 3080 27776 0 net291
rlabel metal2 3864 47768 3864 47768 0 net292
rlabel metal2 4872 48160 4872 48160 0 net293
rlabel metal3 3360 28616 3360 28616 0 net294
rlabel metal2 3080 29344 3080 29344 0 net295
rlabel metal2 4872 30912 4872 30912 0 net296
rlabel metal2 3080 30072 3080 30072 0 net297
rlabel metal2 3080 31024 3080 31024 0 net298
rlabel metal2 3080 31640 3080 31640 0 net299
rlabel metal2 4648 5096 4648 5096 0 net3
rlabel metal2 9072 8120 9072 8120 0 net30
rlabel metal2 3640 32368 3640 32368 0 net300
rlabel metal2 75096 71568 75096 71568 0 net301
rlabel metal2 71960 71288 71960 71288 0 net302
rlabel metal2 72520 72632 72520 72632 0 net303
rlabel metal2 76776 72856 76776 72856 0 net304
rlabel metal2 3976 71288 3976 71288 0 net305
rlabel metal2 4872 71680 4872 71680 0 net306
rlabel metal2 3864 73080 3864 73080 0 net307
rlabel metal2 4872 73248 4872 73248 0 net308
rlabel metal2 74088 72856 74088 72856 0 net309
rlabel metal2 8904 6020 8904 6020 0 net31
rlabel metal2 3640 73696 3640 73696 0 net310
rlabel metal2 74984 71512 74984 71512 0 net311
rlabel metal2 3080 70448 3080 70448 0 net312
rlabel metal3 10136 9688 10136 9688 0 net32
rlabel metal2 10528 4200 10528 4200 0 net33
rlabel metal2 11312 11256 11312 11256 0 net34
rlabel metal3 74928 70728 74928 70728 0 net35
rlabel metal3 72240 49112 72240 49112 0 net36
rlabel metal2 56504 53872 56504 53872 0 net37
rlabel metal2 74928 57512 74928 57512 0 net38
rlabel metal2 75096 57400 75096 57400 0 net39
rlabel metal3 13104 11368 13104 11368 0 net4
rlabel metal2 75208 57904 75208 57904 0 net40
rlabel metal2 63336 58968 63336 58968 0 net41
rlabel metal2 74872 59248 74872 59248 0 net42
rlabel metal2 74760 60424 74760 60424 0 net43
rlabel metal2 72968 59976 72968 59976 0 net44
rlabel metal2 75096 61208 75096 61208 0 net45
rlabel metal2 74648 61936 74648 61936 0 net46
rlabel metal3 49952 47320 49952 47320 0 net47
rlabel metal2 75208 62552 75208 62552 0 net48
rlabel metal2 74984 64568 74984 64568 0 net49
rlabel metal2 13608 6300 13608 6300 0 net5
rlabel metal2 74984 65184 74984 65184 0 net50
rlabel metal2 75096 65520 75096 65520 0 net51
rlabel metal2 64680 64400 64680 64400 0 net52
rlabel metal2 75208 66024 75208 66024 0 net53
rlabel metal2 64904 67144 64904 67144 0 net54
rlabel metal2 75208 67816 75208 67816 0 net55
rlabel metal2 74984 69440 74984 69440 0 net56
rlabel metal2 75096 69160 75096 69160 0 net57
rlabel metal2 51240 49168 51240 49168 0 net58
rlabel metal2 74984 70560 74984 70560 0 net59
rlabel metal2 12824 13608 12824 13608 0 net6
rlabel metal2 68600 69104 68600 69104 0 net60
rlabel metal3 51800 49672 51800 49672 0 net61
rlabel metal3 52080 50568 52080 50568 0 net62
rlabel metal2 75096 52472 75096 52472 0 net63
rlabel metal2 61432 53032 61432 53032 0 net64
rlabel metal2 75096 54152 75096 54152 0 net65
rlabel metal2 53648 53592 53648 53592 0 net66
rlabel metal2 53928 54656 53928 54656 0 net67
rlabel metal3 66920 49112 66920 49112 0 net68
rlabel metal3 51856 54488 51856 54488 0 net69
rlabel metal3 54992 13720 54992 13720 0 net7
rlabel metal2 50680 55104 50680 55104 0 net70
rlabel metal2 3304 58352 3304 58352 0 net71
rlabel metal2 3360 59080 3360 59080 0 net72
rlabel metal2 3304 59920 3304 59920 0 net73
rlabel metal2 3472 60648 3472 60648 0 net74
rlabel metal2 5320 58632 5320 58632 0 net75
rlabel metal2 58520 61320 58520 61320 0 net76
rlabel metal2 3360 62216 3360 62216 0 net77
rlabel metal2 3416 63224 3416 63224 0 net78
rlabel metal2 3360 49672 3360 49672 0 net79
rlabel metal2 55160 14392 55160 14392 0 net8
rlabel metal2 3304 63616 3304 63616 0 net80
rlabel metal2 3360 64792 3360 64792 0 net81
rlabel metal2 3304 65296 3304 65296 0 net82
rlabel metal2 59304 63504 59304 63504 0 net83
rlabel metal2 3304 66136 3304 66136 0 net84
rlabel metal2 3416 66920 3416 66920 0 net85
rlabel metal2 3416 67928 3416 67928 0 net86
rlabel metal2 3192 68096 3192 68096 0 net87
rlabel metal2 3304 69440 3304 69440 0 net88
rlabel metal2 3304 70000 3304 70000 0 net89
rlabel metal2 55384 14952 55384 14952 0 net9
rlabel metal2 3416 50680 3416 50680 0 net90
rlabel metal2 5320 68432 5320 68432 0 net91
rlabel metal2 3304 71008 3304 71008 0 net92
rlabel metal2 3472 51240 3472 51240 0 net93
rlabel metal2 3360 52248 3360 52248 0 net94
rlabel metal2 3360 52808 3360 52808 0 net95
rlabel metal2 3360 53816 3360 53816 0 net96
rlabel metal2 3416 54376 3416 54376 0 net97
rlabel metal3 3640 55384 3640 55384 0 net98
rlabel metal3 3416 54488 3416 54488 0 net99
<< properties >>
string FIXED_BBOX 0 0 80000 80000
<< end >>
