VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_mux
  CLASS BLOCK ;
  FOREIGN wb_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN io_wbs_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.040 0.000 369.600 4.000 ;
    END
  END io_wbs_ack
  PIN io_wbs_ack_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 369.040 400.000 369.600 ;
    END
  END io_wbs_ack_0
  PIN io_wbs_ack_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 369.040 4.000 369.600 ;
    END
  END io_wbs_ack_1
  PIN io_wbs_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.320 0.000 26.880 4.000 ;
    END
  END io_wbs_adr[0]
  PIN io_wbs_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.920 0.000 60.480 4.000 ;
    END
  END io_wbs_adr[10]
  PIN io_wbs_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.280 0.000 63.840 4.000 ;
    END
  END io_wbs_adr[11]
  PIN io_wbs_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.640 0.000 67.200 4.000 ;
    END
  END io_wbs_adr[12]
  PIN io_wbs_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.000 0.000 70.560 4.000 ;
    END
  END io_wbs_adr[13]
  PIN io_wbs_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.360 0.000 73.920 4.000 ;
    END
  END io_wbs_adr[14]
  PIN io_wbs_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 76.720 0.000 77.280 4.000 ;
    END
  END io_wbs_adr[15]
  PIN io_wbs_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.080 0.000 80.640 4.000 ;
    END
  END io_wbs_adr[16]
  PIN io_wbs_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.440 0.000 84.000 4.000 ;
    END
  END io_wbs_adr[17]
  PIN io_wbs_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.800 0.000 87.360 4.000 ;
    END
  END io_wbs_adr[18]
  PIN io_wbs_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.160 0.000 90.720 4.000 ;
    END
  END io_wbs_adr[19]
  PIN io_wbs_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.680 0.000 30.240 4.000 ;
    END
  END io_wbs_adr[1]
  PIN io_wbs_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.520 0.000 94.080 4.000 ;
    END
  END io_wbs_adr[20]
  PIN io_wbs_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 96.880 0.000 97.440 4.000 ;
    END
  END io_wbs_adr[21]
  PIN io_wbs_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.240 0.000 100.800 4.000 ;
    END
  END io_wbs_adr[22]
  PIN io_wbs_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.600 0.000 104.160 4.000 ;
    END
  END io_wbs_adr[23]
  PIN io_wbs_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.960 0.000 107.520 4.000 ;
    END
  END io_wbs_adr[24]
  PIN io_wbs_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.320 0.000 110.880 4.000 ;
    END
  END io_wbs_adr[25]
  PIN io_wbs_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.680 0.000 114.240 4.000 ;
    END
  END io_wbs_adr[26]
  PIN io_wbs_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.040 0.000 117.600 4.000 ;
    END
  END io_wbs_adr[27]
  PIN io_wbs_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.400 0.000 120.960 4.000 ;
    END
  END io_wbs_adr[28]
  PIN io_wbs_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.760 0.000 124.320 4.000 ;
    END
  END io_wbs_adr[29]
  PIN io_wbs_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.040 0.000 33.600 4.000 ;
    END
  END io_wbs_adr[2]
  PIN io_wbs_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.120 0.000 127.680 4.000 ;
    END
  END io_wbs_adr[30]
  PIN io_wbs_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.480 0.000 131.040 4.000 ;
    END
  END io_wbs_adr[31]
  PIN io_wbs_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.400 0.000 36.960 4.000 ;
    END
  END io_wbs_adr[3]
  PIN io_wbs_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 39.760 0.000 40.320 4.000 ;
    END
  END io_wbs_adr[4]
  PIN io_wbs_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.120 0.000 43.680 4.000 ;
    END
  END io_wbs_adr[5]
  PIN io_wbs_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.480 0.000 47.040 4.000 ;
    END
  END io_wbs_adr[6]
  PIN io_wbs_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.840 0.000 50.400 4.000 ;
    END
  END io_wbs_adr[7]
  PIN io_wbs_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.200 0.000 53.760 4.000 ;
    END
  END io_wbs_adr[8]
  PIN io_wbs_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.560 0.000 57.120 4.000 ;
    END
  END io_wbs_adr[9]
  PIN io_wbs_adr_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 26.320 400.000 26.880 ;
    END
  END io_wbs_adr_0[0]
  PIN io_wbs_adr_0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 59.920 400.000 60.480 ;
    END
  END io_wbs_adr_0[10]
  PIN io_wbs_adr_0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 63.280 400.000 63.840 ;
    END
  END io_wbs_adr_0[11]
  PIN io_wbs_adr_0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 66.640 400.000 67.200 ;
    END
  END io_wbs_adr_0[12]
  PIN io_wbs_adr_0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 70.000 400.000 70.560 ;
    END
  END io_wbs_adr_0[13]
  PIN io_wbs_adr_0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 73.360 400.000 73.920 ;
    END
  END io_wbs_adr_0[14]
  PIN io_wbs_adr_0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 76.720 400.000 77.280 ;
    END
  END io_wbs_adr_0[15]
  PIN io_wbs_adr_0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 80.080 400.000 80.640 ;
    END
  END io_wbs_adr_0[16]
  PIN io_wbs_adr_0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 83.440 400.000 84.000 ;
    END
  END io_wbs_adr_0[17]
  PIN io_wbs_adr_0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 86.800 400.000 87.360 ;
    END
  END io_wbs_adr_0[18]
  PIN io_wbs_adr_0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 90.160 400.000 90.720 ;
    END
  END io_wbs_adr_0[19]
  PIN io_wbs_adr_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 29.680 400.000 30.240 ;
    END
  END io_wbs_adr_0[1]
  PIN io_wbs_adr_0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 93.520 400.000 94.080 ;
    END
  END io_wbs_adr_0[20]
  PIN io_wbs_adr_0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 96.880 400.000 97.440 ;
    END
  END io_wbs_adr_0[21]
  PIN io_wbs_adr_0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 100.240 400.000 100.800 ;
    END
  END io_wbs_adr_0[22]
  PIN io_wbs_adr_0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 103.600 400.000 104.160 ;
    END
  END io_wbs_adr_0[23]
  PIN io_wbs_adr_0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 106.960 400.000 107.520 ;
    END
  END io_wbs_adr_0[24]
  PIN io_wbs_adr_0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 110.320 400.000 110.880 ;
    END
  END io_wbs_adr_0[25]
  PIN io_wbs_adr_0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 113.680 400.000 114.240 ;
    END
  END io_wbs_adr_0[26]
  PIN io_wbs_adr_0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 117.040 400.000 117.600 ;
    END
  END io_wbs_adr_0[27]
  PIN io_wbs_adr_0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 120.400 400.000 120.960 ;
    END
  END io_wbs_adr_0[28]
  PIN io_wbs_adr_0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 123.760 400.000 124.320 ;
    END
  END io_wbs_adr_0[29]
  PIN io_wbs_adr_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 33.040 400.000 33.600 ;
    END
  END io_wbs_adr_0[2]
  PIN io_wbs_adr_0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 127.120 400.000 127.680 ;
    END
  END io_wbs_adr_0[30]
  PIN io_wbs_adr_0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 130.480 400.000 131.040 ;
    END
  END io_wbs_adr_0[31]
  PIN io_wbs_adr_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 36.400 400.000 36.960 ;
    END
  END io_wbs_adr_0[3]
  PIN io_wbs_adr_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 39.760 400.000 40.320 ;
    END
  END io_wbs_adr_0[4]
  PIN io_wbs_adr_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 43.120 400.000 43.680 ;
    END
  END io_wbs_adr_0[5]
  PIN io_wbs_adr_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 46.480 400.000 47.040 ;
    END
  END io_wbs_adr_0[6]
  PIN io_wbs_adr_0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 49.840 400.000 50.400 ;
    END
  END io_wbs_adr_0[7]
  PIN io_wbs_adr_0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 53.200 400.000 53.760 ;
    END
  END io_wbs_adr_0[8]
  PIN io_wbs_adr_0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 56.560 400.000 57.120 ;
    END
  END io_wbs_adr_0[9]
  PIN io_wbs_adr_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.320 4.000 26.880 ;
    END
  END io_wbs_adr_1[0]
  PIN io_wbs_adr_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.920 4.000 60.480 ;
    END
  END io_wbs_adr_1[10]
  PIN io_wbs_adr_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.280 4.000 63.840 ;
    END
  END io_wbs_adr_1[11]
  PIN io_wbs_adr_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.640 4.000 67.200 ;
    END
  END io_wbs_adr_1[12]
  PIN io_wbs_adr_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 4.000 70.560 ;
    END
  END io_wbs_adr_1[13]
  PIN io_wbs_adr_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.360 4.000 73.920 ;
    END
  END io_wbs_adr_1[14]
  PIN io_wbs_adr_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 76.720 4.000 77.280 ;
    END
  END io_wbs_adr_1[15]
  PIN io_wbs_adr_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.080 4.000 80.640 ;
    END
  END io_wbs_adr_1[16]
  PIN io_wbs_adr_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 83.440 4.000 84.000 ;
    END
  END io_wbs_adr_1[17]
  PIN io_wbs_adr_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.800 4.000 87.360 ;
    END
  END io_wbs_adr_1[18]
  PIN io_wbs_adr_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.160 4.000 90.720 ;
    END
  END io_wbs_adr_1[19]
  PIN io_wbs_adr_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.680 4.000 30.240 ;
    END
  END io_wbs_adr_1[1]
  PIN io_wbs_adr_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 93.520 4.000 94.080 ;
    END
  END io_wbs_adr_1[20]
  PIN io_wbs_adr_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.880 4.000 97.440 ;
    END
  END io_wbs_adr_1[21]
  PIN io_wbs_adr_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.240 4.000 100.800 ;
    END
  END io_wbs_adr_1[22]
  PIN io_wbs_adr_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 103.600 4.000 104.160 ;
    END
  END io_wbs_adr_1[23]
  PIN io_wbs_adr_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.960 4.000 107.520 ;
    END
  END io_wbs_adr_1[24]
  PIN io_wbs_adr_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.320 4.000 110.880 ;
    END
  END io_wbs_adr_1[25]
  PIN io_wbs_adr_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 113.680 4.000 114.240 ;
    END
  END io_wbs_adr_1[26]
  PIN io_wbs_adr_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.040 4.000 117.600 ;
    END
  END io_wbs_adr_1[27]
  PIN io_wbs_adr_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.400 4.000 120.960 ;
    END
  END io_wbs_adr_1[28]
  PIN io_wbs_adr_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.760 4.000 124.320 ;
    END
  END io_wbs_adr_1[29]
  PIN io_wbs_adr_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.040 4.000 33.600 ;
    END
  END io_wbs_adr_1[2]
  PIN io_wbs_adr_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.120 4.000 127.680 ;
    END
  END io_wbs_adr_1[30]
  PIN io_wbs_adr_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 130.480 4.000 131.040 ;
    END
  END io_wbs_adr_1[31]
  PIN io_wbs_adr_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.400 4.000 36.960 ;
    END
  END io_wbs_adr_1[3]
  PIN io_wbs_adr_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.760 4.000 40.320 ;
    END
  END io_wbs_adr_1[4]
  PIN io_wbs_adr_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.120 4.000 43.680 ;
    END
  END io_wbs_adr_1[5]
  PIN io_wbs_adr_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 46.480 4.000 47.040 ;
    END
  END io_wbs_adr_1[6]
  PIN io_wbs_adr_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 49.840 4.000 50.400 ;
    END
  END io_wbs_adr_1[7]
  PIN io_wbs_adr_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.200 4.000 53.760 ;
    END
  END io_wbs_adr_1[8]
  PIN io_wbs_adr_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.560 4.000 57.120 ;
    END
  END io_wbs_adr_1[9]
  PIN io_wbs_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.400 0.000 372.960 4.000 ;
    END
  END io_wbs_cyc
  PIN io_wbs_cyc_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 372.400 400.000 372.960 ;
    END
  END io_wbs_cyc_0
  PIN io_wbs_cyc_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 372.400 4.000 372.960 ;
    END
  END io_wbs_cyc_1
  PIN io_wbs_datrd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.360 0.000 241.920 4.000 ;
    END
  END io_wbs_datrd[0]
  PIN io_wbs_datrd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 274.960 0.000 275.520 4.000 ;
    END
  END io_wbs_datrd[10]
  PIN io_wbs_datrd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.320 0.000 278.880 4.000 ;
    END
  END io_wbs_datrd[11]
  PIN io_wbs_datrd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.680 0.000 282.240 4.000 ;
    END
  END io_wbs_datrd[12]
  PIN io_wbs_datrd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.040 0.000 285.600 4.000 ;
    END
  END io_wbs_datrd[13]
  PIN io_wbs_datrd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.400 0.000 288.960 4.000 ;
    END
  END io_wbs_datrd[14]
  PIN io_wbs_datrd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.760 0.000 292.320 4.000 ;
    END
  END io_wbs_datrd[15]
  PIN io_wbs_datrd[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.120 0.000 295.680 4.000 ;
    END
  END io_wbs_datrd[16]
  PIN io_wbs_datrd[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 298.480 0.000 299.040 4.000 ;
    END
  END io_wbs_datrd[17]
  PIN io_wbs_datrd[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 301.840 0.000 302.400 4.000 ;
    END
  END io_wbs_datrd[18]
  PIN io_wbs_datrd[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.200 0.000 305.760 4.000 ;
    END
  END io_wbs_datrd[19]
  PIN io_wbs_datrd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 244.720 0.000 245.280 4.000 ;
    END
  END io_wbs_datrd[1]
  PIN io_wbs_datrd[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 308.560 0.000 309.120 4.000 ;
    END
  END io_wbs_datrd[20]
  PIN io_wbs_datrd[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 311.920 0.000 312.480 4.000 ;
    END
  END io_wbs_datrd[21]
  PIN io_wbs_datrd[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.280 0.000 315.840 4.000 ;
    END
  END io_wbs_datrd[22]
  PIN io_wbs_datrd[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.640 0.000 319.200 4.000 ;
    END
  END io_wbs_datrd[23]
  PIN io_wbs_datrd[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.000 0.000 322.560 4.000 ;
    END
  END io_wbs_datrd[24]
  PIN io_wbs_datrd[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.360 0.000 325.920 4.000 ;
    END
  END io_wbs_datrd[25]
  PIN io_wbs_datrd[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.720 0.000 329.280 4.000 ;
    END
  END io_wbs_datrd[26]
  PIN io_wbs_datrd[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.080 0.000 332.640 4.000 ;
    END
  END io_wbs_datrd[27]
  PIN io_wbs_datrd[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 335.440 0.000 336.000 4.000 ;
    END
  END io_wbs_datrd[28]
  PIN io_wbs_datrd[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.800 0.000 339.360 4.000 ;
    END
  END io_wbs_datrd[29]
  PIN io_wbs_datrd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.080 0.000 248.640 4.000 ;
    END
  END io_wbs_datrd[2]
  PIN io_wbs_datrd[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.160 0.000 342.720 4.000 ;
    END
  END io_wbs_datrd[30]
  PIN io_wbs_datrd[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 345.520 0.000 346.080 4.000 ;
    END
  END io_wbs_datrd[31]
  PIN io_wbs_datrd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 251.440 0.000 252.000 4.000 ;
    END
  END io_wbs_datrd[3]
  PIN io_wbs_datrd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.800 0.000 255.360 4.000 ;
    END
  END io_wbs_datrd[4]
  PIN io_wbs_datrd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.160 0.000 258.720 4.000 ;
    END
  END io_wbs_datrd[5]
  PIN io_wbs_datrd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 261.520 0.000 262.080 4.000 ;
    END
  END io_wbs_datrd[6]
  PIN io_wbs_datrd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 264.880 0.000 265.440 4.000 ;
    END
  END io_wbs_datrd[7]
  PIN io_wbs_datrd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.240 0.000 268.800 4.000 ;
    END
  END io_wbs_datrd[8]
  PIN io_wbs_datrd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.600 0.000 272.160 4.000 ;
    END
  END io_wbs_datrd[9]
  PIN io_wbs_datrd_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 241.360 400.000 241.920 ;
    END
  END io_wbs_datrd_0[0]
  PIN io_wbs_datrd_0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 274.960 400.000 275.520 ;
    END
  END io_wbs_datrd_0[10]
  PIN io_wbs_datrd_0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 278.320 400.000 278.880 ;
    END
  END io_wbs_datrd_0[11]
  PIN io_wbs_datrd_0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 281.680 400.000 282.240 ;
    END
  END io_wbs_datrd_0[12]
  PIN io_wbs_datrd_0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 285.040 400.000 285.600 ;
    END
  END io_wbs_datrd_0[13]
  PIN io_wbs_datrd_0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 288.400 400.000 288.960 ;
    END
  END io_wbs_datrd_0[14]
  PIN io_wbs_datrd_0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 291.760 400.000 292.320 ;
    END
  END io_wbs_datrd_0[15]
  PIN io_wbs_datrd_0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 295.120 400.000 295.680 ;
    END
  END io_wbs_datrd_0[16]
  PIN io_wbs_datrd_0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 298.480 400.000 299.040 ;
    END
  END io_wbs_datrd_0[17]
  PIN io_wbs_datrd_0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 301.840 400.000 302.400 ;
    END
  END io_wbs_datrd_0[18]
  PIN io_wbs_datrd_0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 305.200 400.000 305.760 ;
    END
  END io_wbs_datrd_0[19]
  PIN io_wbs_datrd_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 244.720 400.000 245.280 ;
    END
  END io_wbs_datrd_0[1]
  PIN io_wbs_datrd_0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 308.560 400.000 309.120 ;
    END
  END io_wbs_datrd_0[20]
  PIN io_wbs_datrd_0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 311.920 400.000 312.480 ;
    END
  END io_wbs_datrd_0[21]
  PIN io_wbs_datrd_0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 315.280 400.000 315.840 ;
    END
  END io_wbs_datrd_0[22]
  PIN io_wbs_datrd_0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 318.640 400.000 319.200 ;
    END
  END io_wbs_datrd_0[23]
  PIN io_wbs_datrd_0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 322.000 400.000 322.560 ;
    END
  END io_wbs_datrd_0[24]
  PIN io_wbs_datrd_0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 325.360 400.000 325.920 ;
    END
  END io_wbs_datrd_0[25]
  PIN io_wbs_datrd_0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 328.720 400.000 329.280 ;
    END
  END io_wbs_datrd_0[26]
  PIN io_wbs_datrd_0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 332.080 400.000 332.640 ;
    END
  END io_wbs_datrd_0[27]
  PIN io_wbs_datrd_0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 335.440 400.000 336.000 ;
    END
  END io_wbs_datrd_0[28]
  PIN io_wbs_datrd_0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 338.800 400.000 339.360 ;
    END
  END io_wbs_datrd_0[29]
  PIN io_wbs_datrd_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 248.080 400.000 248.640 ;
    END
  END io_wbs_datrd_0[2]
  PIN io_wbs_datrd_0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 342.160 400.000 342.720 ;
    END
  END io_wbs_datrd_0[30]
  PIN io_wbs_datrd_0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 345.520 400.000 346.080 ;
    END
  END io_wbs_datrd_0[31]
  PIN io_wbs_datrd_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 251.440 400.000 252.000 ;
    END
  END io_wbs_datrd_0[3]
  PIN io_wbs_datrd_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 254.800 400.000 255.360 ;
    END
  END io_wbs_datrd_0[4]
  PIN io_wbs_datrd_0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 258.160 400.000 258.720 ;
    END
  END io_wbs_datrd_0[5]
  PIN io_wbs_datrd_0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 261.520 400.000 262.080 ;
    END
  END io_wbs_datrd_0[6]
  PIN io_wbs_datrd_0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 264.880 400.000 265.440 ;
    END
  END io_wbs_datrd_0[7]
  PIN io_wbs_datrd_0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 268.240 400.000 268.800 ;
    END
  END io_wbs_datrd_0[8]
  PIN io_wbs_datrd_0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 271.600 400.000 272.160 ;
    END
  END io_wbs_datrd_0[9]
  PIN io_wbs_datrd_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.360 4.000 241.920 ;
    END
  END io_wbs_datrd_1[0]
  PIN io_wbs_datrd_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 274.960 4.000 275.520 ;
    END
  END io_wbs_datrd_1[10]
  PIN io_wbs_datrd_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.320 4.000 278.880 ;
    END
  END io_wbs_datrd_1[11]
  PIN io_wbs_datrd_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 281.680 4.000 282.240 ;
    END
  END io_wbs_datrd_1[12]
  PIN io_wbs_datrd_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.040 4.000 285.600 ;
    END
  END io_wbs_datrd_1[13]
  PIN io_wbs_datrd_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 288.400 4.000 288.960 ;
    END
  END io_wbs_datrd_1[14]
  PIN io_wbs_datrd_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 291.760 4.000 292.320 ;
    END
  END io_wbs_datrd_1[15]
  PIN io_wbs_datrd_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 295.120 4.000 295.680 ;
    END
  END io_wbs_datrd_1[16]
  PIN io_wbs_datrd_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 298.480 4.000 299.040 ;
    END
  END io_wbs_datrd_1[17]
  PIN io_wbs_datrd_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 301.840 4.000 302.400 ;
    END
  END io_wbs_datrd_1[18]
  PIN io_wbs_datrd_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 305.200 4.000 305.760 ;
    END
  END io_wbs_datrd_1[19]
  PIN io_wbs_datrd_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 244.720 4.000 245.280 ;
    END
  END io_wbs_datrd_1[1]
  PIN io_wbs_datrd_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 308.560 4.000 309.120 ;
    END
  END io_wbs_datrd_1[20]
  PIN io_wbs_datrd_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 311.920 4.000 312.480 ;
    END
  END io_wbs_datrd_1[21]
  PIN io_wbs_datrd_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 315.280 4.000 315.840 ;
    END
  END io_wbs_datrd_1[22]
  PIN io_wbs_datrd_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.640 4.000 319.200 ;
    END
  END io_wbs_datrd_1[23]
  PIN io_wbs_datrd_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 322.000 4.000 322.560 ;
    END
  END io_wbs_datrd_1[24]
  PIN io_wbs_datrd_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 325.360 4.000 325.920 ;
    END
  END io_wbs_datrd_1[25]
  PIN io_wbs_datrd_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 328.720 4.000 329.280 ;
    END
  END io_wbs_datrd_1[26]
  PIN io_wbs_datrd_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 332.080 4.000 332.640 ;
    END
  END io_wbs_datrd_1[27]
  PIN io_wbs_datrd_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 335.440 4.000 336.000 ;
    END
  END io_wbs_datrd_1[28]
  PIN io_wbs_datrd_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 338.800 4.000 339.360 ;
    END
  END io_wbs_datrd_1[29]
  PIN io_wbs_datrd_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 248.080 4.000 248.640 ;
    END
  END io_wbs_datrd_1[2]
  PIN io_wbs_datrd_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.160 4.000 342.720 ;
    END
  END io_wbs_datrd_1[30]
  PIN io_wbs_datrd_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 345.520 4.000 346.080 ;
    END
  END io_wbs_datrd_1[31]
  PIN io_wbs_datrd_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 251.440 4.000 252.000 ;
    END
  END io_wbs_datrd_1[3]
  PIN io_wbs_datrd_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.800 4.000 255.360 ;
    END
  END io_wbs_datrd_1[4]
  PIN io_wbs_datrd_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.160 4.000 258.720 ;
    END
  END io_wbs_datrd_1[5]
  PIN io_wbs_datrd_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 261.520 4.000 262.080 ;
    END
  END io_wbs_datrd_1[6]
  PIN io_wbs_datrd_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 264.880 4.000 265.440 ;
    END
  END io_wbs_datrd_1[7]
  PIN io_wbs_datrd_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 268.240 4.000 268.800 ;
    END
  END io_wbs_datrd_1[8]
  PIN io_wbs_datrd_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 271.600 4.000 272.160 ;
    END
  END io_wbs_datrd_1[9]
  PIN io_wbs_datwr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.840 0.000 134.400 4.000 ;
    END
  END io_wbs_datwr[0]
  PIN io_wbs_datwr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.440 0.000 168.000 4.000 ;
    END
  END io_wbs_datwr[10]
  PIN io_wbs_datwr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.800 0.000 171.360 4.000 ;
    END
  END io_wbs_datwr[11]
  PIN io_wbs_datwr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.160 0.000 174.720 4.000 ;
    END
  END io_wbs_datwr[12]
  PIN io_wbs_datwr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 177.520 0.000 178.080 4.000 ;
    END
  END io_wbs_datwr[13]
  PIN io_wbs_datwr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.880 0.000 181.440 4.000 ;
    END
  END io_wbs_datwr[14]
  PIN io_wbs_datwr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.240 0.000 184.800 4.000 ;
    END
  END io_wbs_datwr[15]
  PIN io_wbs_datwr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.600 0.000 188.160 4.000 ;
    END
  END io_wbs_datwr[16]
  PIN io_wbs_datwr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 190.960 0.000 191.520 4.000 ;
    END
  END io_wbs_datwr[17]
  PIN io_wbs_datwr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.320 0.000 194.880 4.000 ;
    END
  END io_wbs_datwr[18]
  PIN io_wbs_datwr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.680 0.000 198.240 4.000 ;
    END
  END io_wbs_datwr[19]
  PIN io_wbs_datwr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.200 0.000 137.760 4.000 ;
    END
  END io_wbs_datwr[1]
  PIN io_wbs_datwr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.040 0.000 201.600 4.000 ;
    END
  END io_wbs_datwr[20]
  PIN io_wbs_datwr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.400 0.000 204.960 4.000 ;
    END
  END io_wbs_datwr[21]
  PIN io_wbs_datwr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 207.760 0.000 208.320 4.000 ;
    END
  END io_wbs_datwr[22]
  PIN io_wbs_datwr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.120 0.000 211.680 4.000 ;
    END
  END io_wbs_datwr[23]
  PIN io_wbs_datwr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 214.480 0.000 215.040 4.000 ;
    END
  END io_wbs_datwr[24]
  PIN io_wbs_datwr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 217.840 0.000 218.400 4.000 ;
    END
  END io_wbs_datwr[25]
  PIN io_wbs_datwr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.200 0.000 221.760 4.000 ;
    END
  END io_wbs_datwr[26]
  PIN io_wbs_datwr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 224.560 0.000 225.120 4.000 ;
    END
  END io_wbs_datwr[27]
  PIN io_wbs_datwr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 227.920 0.000 228.480 4.000 ;
    END
  END io_wbs_datwr[28]
  PIN io_wbs_datwr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.280 0.000 231.840 4.000 ;
    END
  END io_wbs_datwr[29]
  PIN io_wbs_datwr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.560 0.000 141.120 4.000 ;
    END
  END io_wbs_datwr[2]
  PIN io_wbs_datwr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.640 0.000 235.200 4.000 ;
    END
  END io_wbs_datwr[30]
  PIN io_wbs_datwr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.000 0.000 238.560 4.000 ;
    END
  END io_wbs_datwr[31]
  PIN io_wbs_datwr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 143.920 0.000 144.480 4.000 ;
    END
  END io_wbs_datwr[3]
  PIN io_wbs_datwr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.280 0.000 147.840 4.000 ;
    END
  END io_wbs_datwr[4]
  PIN io_wbs_datwr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.640 0.000 151.200 4.000 ;
    END
  END io_wbs_datwr[5]
  PIN io_wbs_datwr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.000 0.000 154.560 4.000 ;
    END
  END io_wbs_datwr[6]
  PIN io_wbs_datwr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.360 0.000 157.920 4.000 ;
    END
  END io_wbs_datwr[7]
  PIN io_wbs_datwr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 160.720 0.000 161.280 4.000 ;
    END
  END io_wbs_datwr[8]
  PIN io_wbs_datwr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.080 0.000 164.640 4.000 ;
    END
  END io_wbs_datwr[9]
  PIN io_wbs_datwr_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 133.840 400.000 134.400 ;
    END
  END io_wbs_datwr_0[0]
  PIN io_wbs_datwr_0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 167.440 400.000 168.000 ;
    END
  END io_wbs_datwr_0[10]
  PIN io_wbs_datwr_0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 170.800 400.000 171.360 ;
    END
  END io_wbs_datwr_0[11]
  PIN io_wbs_datwr_0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 174.160 400.000 174.720 ;
    END
  END io_wbs_datwr_0[12]
  PIN io_wbs_datwr_0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 177.520 400.000 178.080 ;
    END
  END io_wbs_datwr_0[13]
  PIN io_wbs_datwr_0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 180.880 400.000 181.440 ;
    END
  END io_wbs_datwr_0[14]
  PIN io_wbs_datwr_0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 184.240 400.000 184.800 ;
    END
  END io_wbs_datwr_0[15]
  PIN io_wbs_datwr_0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 187.600 400.000 188.160 ;
    END
  END io_wbs_datwr_0[16]
  PIN io_wbs_datwr_0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 190.960 400.000 191.520 ;
    END
  END io_wbs_datwr_0[17]
  PIN io_wbs_datwr_0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 194.320 400.000 194.880 ;
    END
  END io_wbs_datwr_0[18]
  PIN io_wbs_datwr_0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 197.680 400.000 198.240 ;
    END
  END io_wbs_datwr_0[19]
  PIN io_wbs_datwr_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 137.200 400.000 137.760 ;
    END
  END io_wbs_datwr_0[1]
  PIN io_wbs_datwr_0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 201.040 400.000 201.600 ;
    END
  END io_wbs_datwr_0[20]
  PIN io_wbs_datwr_0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 204.400 400.000 204.960 ;
    END
  END io_wbs_datwr_0[21]
  PIN io_wbs_datwr_0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 207.760 400.000 208.320 ;
    END
  END io_wbs_datwr_0[22]
  PIN io_wbs_datwr_0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 211.120 400.000 211.680 ;
    END
  END io_wbs_datwr_0[23]
  PIN io_wbs_datwr_0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 214.480 400.000 215.040 ;
    END
  END io_wbs_datwr_0[24]
  PIN io_wbs_datwr_0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 217.840 400.000 218.400 ;
    END
  END io_wbs_datwr_0[25]
  PIN io_wbs_datwr_0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 221.200 400.000 221.760 ;
    END
  END io_wbs_datwr_0[26]
  PIN io_wbs_datwr_0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 224.560 400.000 225.120 ;
    END
  END io_wbs_datwr_0[27]
  PIN io_wbs_datwr_0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 227.920 400.000 228.480 ;
    END
  END io_wbs_datwr_0[28]
  PIN io_wbs_datwr_0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 231.280 400.000 231.840 ;
    END
  END io_wbs_datwr_0[29]
  PIN io_wbs_datwr_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 140.560 400.000 141.120 ;
    END
  END io_wbs_datwr_0[2]
  PIN io_wbs_datwr_0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 234.640 400.000 235.200 ;
    END
  END io_wbs_datwr_0[30]
  PIN io_wbs_datwr_0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 238.000 400.000 238.560 ;
    END
  END io_wbs_datwr_0[31]
  PIN io_wbs_datwr_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 143.920 400.000 144.480 ;
    END
  END io_wbs_datwr_0[3]
  PIN io_wbs_datwr_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 147.280 400.000 147.840 ;
    END
  END io_wbs_datwr_0[4]
  PIN io_wbs_datwr_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 150.640 400.000 151.200 ;
    END
  END io_wbs_datwr_0[5]
  PIN io_wbs_datwr_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 154.000 400.000 154.560 ;
    END
  END io_wbs_datwr_0[6]
  PIN io_wbs_datwr_0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 157.360 400.000 157.920 ;
    END
  END io_wbs_datwr_0[7]
  PIN io_wbs_datwr_0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 160.720 400.000 161.280 ;
    END
  END io_wbs_datwr_0[8]
  PIN io_wbs_datwr_0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 164.080 400.000 164.640 ;
    END
  END io_wbs_datwr_0[9]
  PIN io_wbs_datwr_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.840 4.000 134.400 ;
    END
  END io_wbs_datwr_1[0]
  PIN io_wbs_datwr_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 167.440 4.000 168.000 ;
    END
  END io_wbs_datwr_1[10]
  PIN io_wbs_datwr_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.800 4.000 171.360 ;
    END
  END io_wbs_datwr_1[11]
  PIN io_wbs_datwr_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.160 4.000 174.720 ;
    END
  END io_wbs_datwr_1[12]
  PIN io_wbs_datwr_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 177.520 4.000 178.080 ;
    END
  END io_wbs_datwr_1[13]
  PIN io_wbs_datwr_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 180.880 4.000 181.440 ;
    END
  END io_wbs_datwr_1[14]
  PIN io_wbs_datwr_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.240 4.000 184.800 ;
    END
  END io_wbs_datwr_1[15]
  PIN io_wbs_datwr_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.600 4.000 188.160 ;
    END
  END io_wbs_datwr_1[16]
  PIN io_wbs_datwr_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.960 4.000 191.520 ;
    END
  END io_wbs_datwr_1[17]
  PIN io_wbs_datwr_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.320 4.000 194.880 ;
    END
  END io_wbs_datwr_1[18]
  PIN io_wbs_datwr_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 197.680 4.000 198.240 ;
    END
  END io_wbs_datwr_1[19]
  PIN io_wbs_datwr_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.200 4.000 137.760 ;
    END
  END io_wbs_datwr_1[1]
  PIN io_wbs_datwr_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.040 4.000 201.600 ;
    END
  END io_wbs_datwr_1[20]
  PIN io_wbs_datwr_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.400 4.000 204.960 ;
    END
  END io_wbs_datwr_1[21]
  PIN io_wbs_datwr_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.760 4.000 208.320 ;
    END
  END io_wbs_datwr_1[22]
  PIN io_wbs_datwr_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.120 4.000 211.680 ;
    END
  END io_wbs_datwr_1[23]
  PIN io_wbs_datwr_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.480 4.000 215.040 ;
    END
  END io_wbs_datwr_1[24]
  PIN io_wbs_datwr_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 217.840 4.000 218.400 ;
    END
  END io_wbs_datwr_1[25]
  PIN io_wbs_datwr_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.200 4.000 221.760 ;
    END
  END io_wbs_datwr_1[26]
  PIN io_wbs_datwr_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 224.560 4.000 225.120 ;
    END
  END io_wbs_datwr_1[27]
  PIN io_wbs_datwr_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 227.920 4.000 228.480 ;
    END
  END io_wbs_datwr_1[28]
  PIN io_wbs_datwr_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 231.280 4.000 231.840 ;
    END
  END io_wbs_datwr_1[29]
  PIN io_wbs_datwr_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.560 4.000 141.120 ;
    END
  END io_wbs_datwr_1[2]
  PIN io_wbs_datwr_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.640 4.000 235.200 ;
    END
  END io_wbs_datwr_1[30]
  PIN io_wbs_datwr_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.000 4.000 238.560 ;
    END
  END io_wbs_datwr_1[31]
  PIN io_wbs_datwr_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 143.920 4.000 144.480 ;
    END
  END io_wbs_datwr_1[3]
  PIN io_wbs_datwr_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.280 4.000 147.840 ;
    END
  END io_wbs_datwr_1[4]
  PIN io_wbs_datwr_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.640 4.000 151.200 ;
    END
  END io_wbs_datwr_1[5]
  PIN io_wbs_datwr_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.000 4.000 154.560 ;
    END
  END io_wbs_datwr_1[6]
  PIN io_wbs_datwr_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.360 4.000 157.920 ;
    END
  END io_wbs_datwr_1[7]
  PIN io_wbs_datwr_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 160.720 4.000 161.280 ;
    END
  END io_wbs_datwr_1[8]
  PIN io_wbs_datwr_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.080 4.000 164.640 ;
    END
  END io_wbs_datwr_1[9]
  PIN io_wbs_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.240 0.000 352.800 4.000 ;
    END
  END io_wbs_sel[0]
  PIN io_wbs_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.600 0.000 356.160 4.000 ;
    END
  END io_wbs_sel[1]
  PIN io_wbs_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 358.960 0.000 359.520 4.000 ;
    END
  END io_wbs_sel[2]
  PIN io_wbs_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.320 0.000 362.880 4.000 ;
    END
  END io_wbs_sel[3]
  PIN io_wbs_sel_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 352.240 400.000 352.800 ;
    END
  END io_wbs_sel_0[0]
  PIN io_wbs_sel_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 355.600 400.000 356.160 ;
    END
  END io_wbs_sel_0[1]
  PIN io_wbs_sel_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 358.960 400.000 359.520 ;
    END
  END io_wbs_sel_0[2]
  PIN io_wbs_sel_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 362.320 400.000 362.880 ;
    END
  END io_wbs_sel_0[3]
  PIN io_wbs_sel_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.240 4.000 352.800 ;
    END
  END io_wbs_sel_1[0]
  PIN io_wbs_sel_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 355.600 4.000 356.160 ;
    END
  END io_wbs_sel_1[1]
  PIN io_wbs_sel_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.960 4.000 359.520 ;
    END
  END io_wbs_sel_1[2]
  PIN io_wbs_sel_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.320 4.000 362.880 ;
    END
  END io_wbs_sel_1[3]
  PIN io_wbs_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.680 0.000 366.240 4.000 ;
    END
  END io_wbs_stb
  PIN io_wbs_stb_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 365.680 400.000 366.240 ;
    END
  END io_wbs_stb_0
  PIN io_wbs_stb_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 365.680 4.000 366.240 ;
    END
  END io_wbs_stb_1
  PIN io_wbs_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.880 0.000 349.440 4.000 ;
    END
  END io_wbs_we
  PIN io_wbs_we_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 348.880 400.000 349.440 ;
    END
  END io_wbs_we_0
  PIN io_wbs_we_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 348.880 4.000 349.440 ;
    END
  END io_wbs_we_1
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 384.460 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 384.460 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 393.120 384.460 ;
      LAYER Metal2 ;
        RECT 8.540 4.300 391.300 384.350 ;
        RECT 8.540 3.500 26.020 4.300 ;
        RECT 27.180 3.500 29.380 4.300 ;
        RECT 30.540 3.500 32.740 4.300 ;
        RECT 33.900 3.500 36.100 4.300 ;
        RECT 37.260 3.500 39.460 4.300 ;
        RECT 40.620 3.500 42.820 4.300 ;
        RECT 43.980 3.500 46.180 4.300 ;
        RECT 47.340 3.500 49.540 4.300 ;
        RECT 50.700 3.500 52.900 4.300 ;
        RECT 54.060 3.500 56.260 4.300 ;
        RECT 57.420 3.500 59.620 4.300 ;
        RECT 60.780 3.500 62.980 4.300 ;
        RECT 64.140 3.500 66.340 4.300 ;
        RECT 67.500 3.500 69.700 4.300 ;
        RECT 70.860 3.500 73.060 4.300 ;
        RECT 74.220 3.500 76.420 4.300 ;
        RECT 77.580 3.500 79.780 4.300 ;
        RECT 80.940 3.500 83.140 4.300 ;
        RECT 84.300 3.500 86.500 4.300 ;
        RECT 87.660 3.500 89.860 4.300 ;
        RECT 91.020 3.500 93.220 4.300 ;
        RECT 94.380 3.500 96.580 4.300 ;
        RECT 97.740 3.500 99.940 4.300 ;
        RECT 101.100 3.500 103.300 4.300 ;
        RECT 104.460 3.500 106.660 4.300 ;
        RECT 107.820 3.500 110.020 4.300 ;
        RECT 111.180 3.500 113.380 4.300 ;
        RECT 114.540 3.500 116.740 4.300 ;
        RECT 117.900 3.500 120.100 4.300 ;
        RECT 121.260 3.500 123.460 4.300 ;
        RECT 124.620 3.500 126.820 4.300 ;
        RECT 127.980 3.500 130.180 4.300 ;
        RECT 131.340 3.500 133.540 4.300 ;
        RECT 134.700 3.500 136.900 4.300 ;
        RECT 138.060 3.500 140.260 4.300 ;
        RECT 141.420 3.500 143.620 4.300 ;
        RECT 144.780 3.500 146.980 4.300 ;
        RECT 148.140 3.500 150.340 4.300 ;
        RECT 151.500 3.500 153.700 4.300 ;
        RECT 154.860 3.500 157.060 4.300 ;
        RECT 158.220 3.500 160.420 4.300 ;
        RECT 161.580 3.500 163.780 4.300 ;
        RECT 164.940 3.500 167.140 4.300 ;
        RECT 168.300 3.500 170.500 4.300 ;
        RECT 171.660 3.500 173.860 4.300 ;
        RECT 175.020 3.500 177.220 4.300 ;
        RECT 178.380 3.500 180.580 4.300 ;
        RECT 181.740 3.500 183.940 4.300 ;
        RECT 185.100 3.500 187.300 4.300 ;
        RECT 188.460 3.500 190.660 4.300 ;
        RECT 191.820 3.500 194.020 4.300 ;
        RECT 195.180 3.500 197.380 4.300 ;
        RECT 198.540 3.500 200.740 4.300 ;
        RECT 201.900 3.500 204.100 4.300 ;
        RECT 205.260 3.500 207.460 4.300 ;
        RECT 208.620 3.500 210.820 4.300 ;
        RECT 211.980 3.500 214.180 4.300 ;
        RECT 215.340 3.500 217.540 4.300 ;
        RECT 218.700 3.500 220.900 4.300 ;
        RECT 222.060 3.500 224.260 4.300 ;
        RECT 225.420 3.500 227.620 4.300 ;
        RECT 228.780 3.500 230.980 4.300 ;
        RECT 232.140 3.500 234.340 4.300 ;
        RECT 235.500 3.500 237.700 4.300 ;
        RECT 238.860 3.500 241.060 4.300 ;
        RECT 242.220 3.500 244.420 4.300 ;
        RECT 245.580 3.500 247.780 4.300 ;
        RECT 248.940 3.500 251.140 4.300 ;
        RECT 252.300 3.500 254.500 4.300 ;
        RECT 255.660 3.500 257.860 4.300 ;
        RECT 259.020 3.500 261.220 4.300 ;
        RECT 262.380 3.500 264.580 4.300 ;
        RECT 265.740 3.500 267.940 4.300 ;
        RECT 269.100 3.500 271.300 4.300 ;
        RECT 272.460 3.500 274.660 4.300 ;
        RECT 275.820 3.500 278.020 4.300 ;
        RECT 279.180 3.500 281.380 4.300 ;
        RECT 282.540 3.500 284.740 4.300 ;
        RECT 285.900 3.500 288.100 4.300 ;
        RECT 289.260 3.500 291.460 4.300 ;
        RECT 292.620 3.500 294.820 4.300 ;
        RECT 295.980 3.500 298.180 4.300 ;
        RECT 299.340 3.500 301.540 4.300 ;
        RECT 302.700 3.500 304.900 4.300 ;
        RECT 306.060 3.500 308.260 4.300 ;
        RECT 309.420 3.500 311.620 4.300 ;
        RECT 312.780 3.500 314.980 4.300 ;
        RECT 316.140 3.500 318.340 4.300 ;
        RECT 319.500 3.500 321.700 4.300 ;
        RECT 322.860 3.500 325.060 4.300 ;
        RECT 326.220 3.500 328.420 4.300 ;
        RECT 329.580 3.500 331.780 4.300 ;
        RECT 332.940 3.500 335.140 4.300 ;
        RECT 336.300 3.500 338.500 4.300 ;
        RECT 339.660 3.500 341.860 4.300 ;
        RECT 343.020 3.500 345.220 4.300 ;
        RECT 346.380 3.500 348.580 4.300 ;
        RECT 349.740 3.500 351.940 4.300 ;
        RECT 353.100 3.500 355.300 4.300 ;
        RECT 356.460 3.500 358.660 4.300 ;
        RECT 359.820 3.500 362.020 4.300 ;
        RECT 363.180 3.500 365.380 4.300 ;
        RECT 366.540 3.500 368.740 4.300 ;
        RECT 369.900 3.500 372.100 4.300 ;
        RECT 373.260 3.500 391.300 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 373.260 396.340 384.300 ;
        RECT 4.300 372.100 395.700 373.260 ;
        RECT 4.000 369.900 396.340 372.100 ;
        RECT 4.300 368.740 395.700 369.900 ;
        RECT 4.000 366.540 396.340 368.740 ;
        RECT 4.300 365.380 395.700 366.540 ;
        RECT 4.000 363.180 396.340 365.380 ;
        RECT 4.300 362.020 395.700 363.180 ;
        RECT 4.000 359.820 396.340 362.020 ;
        RECT 4.300 358.660 395.700 359.820 ;
        RECT 4.000 356.460 396.340 358.660 ;
        RECT 4.300 355.300 395.700 356.460 ;
        RECT 4.000 353.100 396.340 355.300 ;
        RECT 4.300 351.940 395.700 353.100 ;
        RECT 4.000 349.740 396.340 351.940 ;
        RECT 4.300 348.580 395.700 349.740 ;
        RECT 4.000 346.380 396.340 348.580 ;
        RECT 4.300 345.220 395.700 346.380 ;
        RECT 4.000 343.020 396.340 345.220 ;
        RECT 4.300 341.860 395.700 343.020 ;
        RECT 4.000 339.660 396.340 341.860 ;
        RECT 4.300 338.500 395.700 339.660 ;
        RECT 4.000 336.300 396.340 338.500 ;
        RECT 4.300 335.140 395.700 336.300 ;
        RECT 4.000 332.940 396.340 335.140 ;
        RECT 4.300 331.780 395.700 332.940 ;
        RECT 4.000 329.580 396.340 331.780 ;
        RECT 4.300 328.420 395.700 329.580 ;
        RECT 4.000 326.220 396.340 328.420 ;
        RECT 4.300 325.060 395.700 326.220 ;
        RECT 4.000 322.860 396.340 325.060 ;
        RECT 4.300 321.700 395.700 322.860 ;
        RECT 4.000 319.500 396.340 321.700 ;
        RECT 4.300 318.340 395.700 319.500 ;
        RECT 4.000 316.140 396.340 318.340 ;
        RECT 4.300 314.980 395.700 316.140 ;
        RECT 4.000 312.780 396.340 314.980 ;
        RECT 4.300 311.620 395.700 312.780 ;
        RECT 4.000 309.420 396.340 311.620 ;
        RECT 4.300 308.260 395.700 309.420 ;
        RECT 4.000 306.060 396.340 308.260 ;
        RECT 4.300 304.900 395.700 306.060 ;
        RECT 4.000 302.700 396.340 304.900 ;
        RECT 4.300 301.540 395.700 302.700 ;
        RECT 4.000 299.340 396.340 301.540 ;
        RECT 4.300 298.180 395.700 299.340 ;
        RECT 4.000 295.980 396.340 298.180 ;
        RECT 4.300 294.820 395.700 295.980 ;
        RECT 4.000 292.620 396.340 294.820 ;
        RECT 4.300 291.460 395.700 292.620 ;
        RECT 4.000 289.260 396.340 291.460 ;
        RECT 4.300 288.100 395.700 289.260 ;
        RECT 4.000 285.900 396.340 288.100 ;
        RECT 4.300 284.740 395.700 285.900 ;
        RECT 4.000 282.540 396.340 284.740 ;
        RECT 4.300 281.380 395.700 282.540 ;
        RECT 4.000 279.180 396.340 281.380 ;
        RECT 4.300 278.020 395.700 279.180 ;
        RECT 4.000 275.820 396.340 278.020 ;
        RECT 4.300 274.660 395.700 275.820 ;
        RECT 4.000 272.460 396.340 274.660 ;
        RECT 4.300 271.300 395.700 272.460 ;
        RECT 4.000 269.100 396.340 271.300 ;
        RECT 4.300 267.940 395.700 269.100 ;
        RECT 4.000 265.740 396.340 267.940 ;
        RECT 4.300 264.580 395.700 265.740 ;
        RECT 4.000 262.380 396.340 264.580 ;
        RECT 4.300 261.220 395.700 262.380 ;
        RECT 4.000 259.020 396.340 261.220 ;
        RECT 4.300 257.860 395.700 259.020 ;
        RECT 4.000 255.660 396.340 257.860 ;
        RECT 4.300 254.500 395.700 255.660 ;
        RECT 4.000 252.300 396.340 254.500 ;
        RECT 4.300 251.140 395.700 252.300 ;
        RECT 4.000 248.940 396.340 251.140 ;
        RECT 4.300 247.780 395.700 248.940 ;
        RECT 4.000 245.580 396.340 247.780 ;
        RECT 4.300 244.420 395.700 245.580 ;
        RECT 4.000 242.220 396.340 244.420 ;
        RECT 4.300 241.060 395.700 242.220 ;
        RECT 4.000 238.860 396.340 241.060 ;
        RECT 4.300 237.700 395.700 238.860 ;
        RECT 4.000 235.500 396.340 237.700 ;
        RECT 4.300 234.340 395.700 235.500 ;
        RECT 4.000 232.140 396.340 234.340 ;
        RECT 4.300 230.980 395.700 232.140 ;
        RECT 4.000 228.780 396.340 230.980 ;
        RECT 4.300 227.620 395.700 228.780 ;
        RECT 4.000 225.420 396.340 227.620 ;
        RECT 4.300 224.260 395.700 225.420 ;
        RECT 4.000 222.060 396.340 224.260 ;
        RECT 4.300 220.900 395.700 222.060 ;
        RECT 4.000 218.700 396.340 220.900 ;
        RECT 4.300 217.540 395.700 218.700 ;
        RECT 4.000 215.340 396.340 217.540 ;
        RECT 4.300 214.180 395.700 215.340 ;
        RECT 4.000 211.980 396.340 214.180 ;
        RECT 4.300 210.820 395.700 211.980 ;
        RECT 4.000 208.620 396.340 210.820 ;
        RECT 4.300 207.460 395.700 208.620 ;
        RECT 4.000 205.260 396.340 207.460 ;
        RECT 4.300 204.100 395.700 205.260 ;
        RECT 4.000 201.900 396.340 204.100 ;
        RECT 4.300 200.740 395.700 201.900 ;
        RECT 4.000 198.540 396.340 200.740 ;
        RECT 4.300 197.380 395.700 198.540 ;
        RECT 4.000 195.180 396.340 197.380 ;
        RECT 4.300 194.020 395.700 195.180 ;
        RECT 4.000 191.820 396.340 194.020 ;
        RECT 4.300 190.660 395.700 191.820 ;
        RECT 4.000 188.460 396.340 190.660 ;
        RECT 4.300 187.300 395.700 188.460 ;
        RECT 4.000 185.100 396.340 187.300 ;
        RECT 4.300 183.940 395.700 185.100 ;
        RECT 4.000 181.740 396.340 183.940 ;
        RECT 4.300 180.580 395.700 181.740 ;
        RECT 4.000 178.380 396.340 180.580 ;
        RECT 4.300 177.220 395.700 178.380 ;
        RECT 4.000 175.020 396.340 177.220 ;
        RECT 4.300 173.860 395.700 175.020 ;
        RECT 4.000 171.660 396.340 173.860 ;
        RECT 4.300 170.500 395.700 171.660 ;
        RECT 4.000 168.300 396.340 170.500 ;
        RECT 4.300 167.140 395.700 168.300 ;
        RECT 4.000 164.940 396.340 167.140 ;
        RECT 4.300 163.780 395.700 164.940 ;
        RECT 4.000 161.580 396.340 163.780 ;
        RECT 4.300 160.420 395.700 161.580 ;
        RECT 4.000 158.220 396.340 160.420 ;
        RECT 4.300 157.060 395.700 158.220 ;
        RECT 4.000 154.860 396.340 157.060 ;
        RECT 4.300 153.700 395.700 154.860 ;
        RECT 4.000 151.500 396.340 153.700 ;
        RECT 4.300 150.340 395.700 151.500 ;
        RECT 4.000 148.140 396.340 150.340 ;
        RECT 4.300 146.980 395.700 148.140 ;
        RECT 4.000 144.780 396.340 146.980 ;
        RECT 4.300 143.620 395.700 144.780 ;
        RECT 4.000 141.420 396.340 143.620 ;
        RECT 4.300 140.260 395.700 141.420 ;
        RECT 4.000 138.060 396.340 140.260 ;
        RECT 4.300 136.900 395.700 138.060 ;
        RECT 4.000 134.700 396.340 136.900 ;
        RECT 4.300 133.540 395.700 134.700 ;
        RECT 4.000 131.340 396.340 133.540 ;
        RECT 4.300 130.180 395.700 131.340 ;
        RECT 4.000 127.980 396.340 130.180 ;
        RECT 4.300 126.820 395.700 127.980 ;
        RECT 4.000 124.620 396.340 126.820 ;
        RECT 4.300 123.460 395.700 124.620 ;
        RECT 4.000 121.260 396.340 123.460 ;
        RECT 4.300 120.100 395.700 121.260 ;
        RECT 4.000 117.900 396.340 120.100 ;
        RECT 4.300 116.740 395.700 117.900 ;
        RECT 4.000 114.540 396.340 116.740 ;
        RECT 4.300 113.380 395.700 114.540 ;
        RECT 4.000 111.180 396.340 113.380 ;
        RECT 4.300 110.020 395.700 111.180 ;
        RECT 4.000 107.820 396.340 110.020 ;
        RECT 4.300 106.660 395.700 107.820 ;
        RECT 4.000 104.460 396.340 106.660 ;
        RECT 4.300 103.300 395.700 104.460 ;
        RECT 4.000 101.100 396.340 103.300 ;
        RECT 4.300 99.940 395.700 101.100 ;
        RECT 4.000 97.740 396.340 99.940 ;
        RECT 4.300 96.580 395.700 97.740 ;
        RECT 4.000 94.380 396.340 96.580 ;
        RECT 4.300 93.220 395.700 94.380 ;
        RECT 4.000 91.020 396.340 93.220 ;
        RECT 4.300 89.860 395.700 91.020 ;
        RECT 4.000 87.660 396.340 89.860 ;
        RECT 4.300 86.500 395.700 87.660 ;
        RECT 4.000 84.300 396.340 86.500 ;
        RECT 4.300 83.140 395.700 84.300 ;
        RECT 4.000 80.940 396.340 83.140 ;
        RECT 4.300 79.780 395.700 80.940 ;
        RECT 4.000 77.580 396.340 79.780 ;
        RECT 4.300 76.420 395.700 77.580 ;
        RECT 4.000 74.220 396.340 76.420 ;
        RECT 4.300 73.060 395.700 74.220 ;
        RECT 4.000 70.860 396.340 73.060 ;
        RECT 4.300 69.700 395.700 70.860 ;
        RECT 4.000 67.500 396.340 69.700 ;
        RECT 4.300 66.340 395.700 67.500 ;
        RECT 4.000 64.140 396.340 66.340 ;
        RECT 4.300 62.980 395.700 64.140 ;
        RECT 4.000 60.780 396.340 62.980 ;
        RECT 4.300 59.620 395.700 60.780 ;
        RECT 4.000 57.420 396.340 59.620 ;
        RECT 4.300 56.260 395.700 57.420 ;
        RECT 4.000 54.060 396.340 56.260 ;
        RECT 4.300 52.900 395.700 54.060 ;
        RECT 4.000 50.700 396.340 52.900 ;
        RECT 4.300 49.540 395.700 50.700 ;
        RECT 4.000 47.340 396.340 49.540 ;
        RECT 4.300 46.180 395.700 47.340 ;
        RECT 4.000 43.980 396.340 46.180 ;
        RECT 4.300 42.820 395.700 43.980 ;
        RECT 4.000 40.620 396.340 42.820 ;
        RECT 4.300 39.460 395.700 40.620 ;
        RECT 4.000 37.260 396.340 39.460 ;
        RECT 4.300 36.100 395.700 37.260 ;
        RECT 4.000 33.900 396.340 36.100 ;
        RECT 4.300 32.740 395.700 33.900 ;
        RECT 4.000 30.540 396.340 32.740 ;
        RECT 4.300 29.380 395.700 30.540 ;
        RECT 4.000 27.180 396.340 29.380 ;
        RECT 4.300 26.020 395.700 27.180 ;
        RECT 4.000 15.540 396.340 26.020 ;
      LAYER Metal4 ;
        RECT 259.980 247.050 329.140 333.670 ;
        RECT 331.340 247.050 342.020 333.670 ;
  END
END wb_mux
END LIBRARY

