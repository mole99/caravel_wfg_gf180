magic
tech gf180mcuC
magscale 1 5
timestamp 1670254938
<< obsm1 >>
rect 672 1538 74392 18454
<< metal2 >>
rect 2576 0 2632 400
rect 3416 0 3472 400
rect 4256 0 4312 400
rect 5096 0 5152 400
rect 5936 0 5992 400
rect 6776 0 6832 400
rect 7616 0 7672 400
rect 8456 0 8512 400
rect 9296 0 9352 400
rect 10136 0 10192 400
rect 10976 0 11032 400
rect 11816 0 11872 400
rect 12656 0 12712 400
rect 13496 0 13552 400
rect 14336 0 14392 400
rect 15176 0 15232 400
rect 16016 0 16072 400
rect 16856 0 16912 400
rect 17696 0 17752 400
rect 18536 0 18592 400
rect 19376 0 19432 400
rect 20216 0 20272 400
rect 21056 0 21112 400
rect 21896 0 21952 400
rect 22736 0 22792 400
rect 23576 0 23632 400
rect 24416 0 24472 400
rect 25256 0 25312 400
rect 26096 0 26152 400
rect 26936 0 26992 400
rect 27776 0 27832 400
rect 28616 0 28672 400
rect 29456 0 29512 400
rect 30296 0 30352 400
rect 31136 0 31192 400
rect 31976 0 32032 400
rect 32816 0 32872 400
rect 33656 0 33712 400
rect 34496 0 34552 400
rect 35336 0 35392 400
rect 36176 0 36232 400
rect 37016 0 37072 400
rect 37856 0 37912 400
rect 38696 0 38752 400
rect 39536 0 39592 400
rect 40376 0 40432 400
rect 41216 0 41272 400
rect 42056 0 42112 400
rect 42896 0 42952 400
rect 43736 0 43792 400
rect 44576 0 44632 400
rect 45416 0 45472 400
rect 46256 0 46312 400
rect 47096 0 47152 400
rect 47936 0 47992 400
rect 48776 0 48832 400
rect 49616 0 49672 400
rect 50456 0 50512 400
rect 51296 0 51352 400
rect 52136 0 52192 400
rect 52976 0 53032 400
rect 53816 0 53872 400
rect 54656 0 54712 400
rect 55496 0 55552 400
rect 56336 0 56392 400
rect 57176 0 57232 400
rect 58016 0 58072 400
rect 58856 0 58912 400
rect 59696 0 59752 400
rect 60536 0 60592 400
rect 61376 0 61432 400
rect 62216 0 62272 400
rect 63056 0 63112 400
rect 63896 0 63952 400
rect 64736 0 64792 400
rect 65576 0 65632 400
rect 66416 0 66472 400
rect 67256 0 67312 400
rect 68096 0 68152 400
rect 68936 0 68992 400
rect 69776 0 69832 400
rect 70616 0 70672 400
rect 71456 0 71512 400
rect 72296 0 72352 400
<< obsm2 >>
rect 2590 430 74378 19423
rect 2662 350 3386 430
rect 3502 350 4226 430
rect 4342 350 5066 430
rect 5182 350 5906 430
rect 6022 350 6746 430
rect 6862 350 7586 430
rect 7702 350 8426 430
rect 8542 350 9266 430
rect 9382 350 10106 430
rect 10222 350 10946 430
rect 11062 350 11786 430
rect 11902 350 12626 430
rect 12742 350 13466 430
rect 13582 350 14306 430
rect 14422 350 15146 430
rect 15262 350 15986 430
rect 16102 350 16826 430
rect 16942 350 17666 430
rect 17782 350 18506 430
rect 18622 350 19346 430
rect 19462 350 20186 430
rect 20302 350 21026 430
rect 21142 350 21866 430
rect 21982 350 22706 430
rect 22822 350 23546 430
rect 23662 350 24386 430
rect 24502 350 25226 430
rect 25342 350 26066 430
rect 26182 350 26906 430
rect 27022 350 27746 430
rect 27862 350 28586 430
rect 28702 350 29426 430
rect 29542 350 30266 430
rect 30382 350 31106 430
rect 31222 350 31946 430
rect 32062 350 32786 430
rect 32902 350 33626 430
rect 33742 350 34466 430
rect 34582 350 35306 430
rect 35422 350 36146 430
rect 36262 350 36986 430
rect 37102 350 37826 430
rect 37942 350 38666 430
rect 38782 350 39506 430
rect 39622 350 40346 430
rect 40462 350 41186 430
rect 41302 350 42026 430
rect 42142 350 42866 430
rect 42982 350 43706 430
rect 43822 350 44546 430
rect 44662 350 45386 430
rect 45502 350 46226 430
rect 46342 350 47066 430
rect 47182 350 47906 430
rect 48022 350 48746 430
rect 48862 350 49586 430
rect 49702 350 50426 430
rect 50542 350 51266 430
rect 51382 350 52106 430
rect 52222 350 52946 430
rect 53062 350 53786 430
rect 53902 350 54626 430
rect 54742 350 55466 430
rect 55582 350 56306 430
rect 56422 350 57146 430
rect 57262 350 57986 430
rect 58102 350 58826 430
rect 58942 350 59666 430
rect 59782 350 60506 430
rect 60622 350 61346 430
rect 61462 350 62186 430
rect 62302 350 63026 430
rect 63142 350 63866 430
rect 63982 350 64706 430
rect 64822 350 65546 430
rect 65662 350 66386 430
rect 66502 350 67226 430
rect 67342 350 68066 430
rect 68182 350 68906 430
rect 69022 350 69746 430
rect 69862 350 70586 430
rect 70702 350 71426 430
rect 71542 350 72266 430
rect 72382 350 74378 430
<< metal3 >>
rect 74600 19376 75000 19432
rect 74600 18928 75000 18984
rect 74600 18480 75000 18536
rect 74600 18032 75000 18088
rect 74600 17584 75000 17640
rect 74600 17136 75000 17192
rect 74600 16688 75000 16744
rect 74600 16240 75000 16296
rect 74600 15792 75000 15848
rect 74600 15344 75000 15400
rect 74600 14896 75000 14952
rect 74600 14448 75000 14504
rect 74600 14000 75000 14056
rect 74600 13552 75000 13608
rect 74600 13104 75000 13160
rect 74600 12656 75000 12712
rect 74600 12208 75000 12264
rect 74600 11760 75000 11816
rect 74600 11312 75000 11368
rect 74600 10864 75000 10920
rect 74600 10416 75000 10472
rect 74600 9968 75000 10024
rect 74600 9520 75000 9576
rect 74600 9072 75000 9128
rect 74600 8624 75000 8680
rect 74600 8176 75000 8232
rect 74600 7728 75000 7784
rect 74600 7280 75000 7336
rect 74600 6832 75000 6888
rect 74600 6384 75000 6440
rect 74600 5936 75000 5992
rect 74600 5488 75000 5544
rect 74600 5040 75000 5096
rect 74600 4592 75000 4648
rect 74600 4144 75000 4200
rect 74600 3696 75000 3752
rect 74600 3248 75000 3304
rect 74600 2800 75000 2856
rect 74600 2352 75000 2408
rect 74600 1904 75000 1960
rect 74600 1456 75000 1512
rect 74600 1008 75000 1064
rect 74600 560 75000 616
<< obsm3 >>
rect 2585 19346 74570 19418
rect 2585 19014 74600 19346
rect 2585 18898 74570 19014
rect 2585 18566 74600 18898
rect 2585 18450 74570 18566
rect 2585 18118 74600 18450
rect 2585 18002 74570 18118
rect 2585 17670 74600 18002
rect 2585 17554 74570 17670
rect 2585 17222 74600 17554
rect 2585 17106 74570 17222
rect 2585 16774 74600 17106
rect 2585 16658 74570 16774
rect 2585 16326 74600 16658
rect 2585 16210 74570 16326
rect 2585 15878 74600 16210
rect 2585 15762 74570 15878
rect 2585 15430 74600 15762
rect 2585 15314 74570 15430
rect 2585 14982 74600 15314
rect 2585 14866 74570 14982
rect 2585 14534 74600 14866
rect 2585 14418 74570 14534
rect 2585 14086 74600 14418
rect 2585 13970 74570 14086
rect 2585 13638 74600 13970
rect 2585 13522 74570 13638
rect 2585 13190 74600 13522
rect 2585 13074 74570 13190
rect 2585 12742 74600 13074
rect 2585 12626 74570 12742
rect 2585 12294 74600 12626
rect 2585 12178 74570 12294
rect 2585 11846 74600 12178
rect 2585 11730 74570 11846
rect 2585 11398 74600 11730
rect 2585 11282 74570 11398
rect 2585 10950 74600 11282
rect 2585 10834 74570 10950
rect 2585 10502 74600 10834
rect 2585 10386 74570 10502
rect 2585 10054 74600 10386
rect 2585 9938 74570 10054
rect 2585 9606 74600 9938
rect 2585 9490 74570 9606
rect 2585 9158 74600 9490
rect 2585 9042 74570 9158
rect 2585 8710 74600 9042
rect 2585 8594 74570 8710
rect 2585 8262 74600 8594
rect 2585 8146 74570 8262
rect 2585 7814 74600 8146
rect 2585 7698 74570 7814
rect 2585 7366 74600 7698
rect 2585 7250 74570 7366
rect 2585 6918 74600 7250
rect 2585 6802 74570 6918
rect 2585 6470 74600 6802
rect 2585 6354 74570 6470
rect 2585 6022 74600 6354
rect 2585 5906 74570 6022
rect 2585 5574 74600 5906
rect 2585 5458 74570 5574
rect 2585 5126 74600 5458
rect 2585 5010 74570 5126
rect 2585 4678 74600 5010
rect 2585 4562 74570 4678
rect 2585 4230 74600 4562
rect 2585 4114 74570 4230
rect 2585 3782 74600 4114
rect 2585 3666 74570 3782
rect 2585 3334 74600 3666
rect 2585 3218 74570 3334
rect 2585 2886 74600 3218
rect 2585 2770 74570 2886
rect 2585 2438 74600 2770
rect 2585 2322 74570 2438
rect 2585 1990 74600 2322
rect 2585 1874 74570 1990
rect 2585 1542 74600 1874
rect 2585 1426 74570 1542
rect 2585 1094 74600 1426
rect 2585 978 74570 1094
rect 2585 646 74600 978
rect 2585 530 74570 646
rect 2585 406 74600 530
<< metal4 >>
rect 9797 1538 9957 18454
rect 19002 1538 19162 18454
rect 28207 1538 28367 18454
rect 37412 1538 37572 18454
rect 46617 1538 46777 18454
rect 55822 1538 55982 18454
rect 65027 1538 65187 18454
rect 74232 1538 74392 18454
<< obsm4 >>
rect 15246 1689 18972 3015
rect 19192 1689 28177 3015
rect 28397 1689 37382 3015
rect 37602 1689 46587 3015
rect 46807 1689 55792 3015
rect 56012 1689 64997 3015
rect 65217 1689 65506 3015
<< labels >>
rlabel metal3 s 74600 1008 75000 1064 6 addr[0]
port 1 nsew signal input
rlabel metal3 s 74600 1456 75000 1512 6 addr[1]
port 2 nsew signal input
rlabel metal3 s 74600 1904 75000 1960 6 addr[2]
port 3 nsew signal input
rlabel metal3 s 74600 2352 75000 2408 6 addr[3]
port 4 nsew signal input
rlabel metal3 s 74600 2800 75000 2856 6 addr[4]
port 5 nsew signal input
rlabel metal3 s 74600 3248 75000 3304 6 addr[5]
port 6 nsew signal input
rlabel metal3 s 74600 3696 75000 3752 6 addr[6]
port 7 nsew signal input
rlabel metal3 s 74600 4144 75000 4200 6 addr[7]
port 8 nsew signal input
rlabel metal3 s 74600 4592 75000 4648 6 addr[8]
port 9 nsew signal input
rlabel metal3 s 74600 5040 75000 5096 6 addr[9]
port 10 nsew signal input
rlabel metal2 s 3416 0 3472 400 6 addr_mem0[0]
port 11 nsew signal output
rlabel metal2 s 4256 0 4312 400 6 addr_mem0[1]
port 12 nsew signal output
rlabel metal2 s 5096 0 5152 400 6 addr_mem0[2]
port 13 nsew signal output
rlabel metal2 s 5936 0 5992 400 6 addr_mem0[3]
port 14 nsew signal output
rlabel metal2 s 6776 0 6832 400 6 addr_mem0[4]
port 15 nsew signal output
rlabel metal2 s 7616 0 7672 400 6 addr_mem0[5]
port 16 nsew signal output
rlabel metal2 s 8456 0 8512 400 6 addr_mem0[6]
port 17 nsew signal output
rlabel metal2 s 9296 0 9352 400 6 addr_mem0[7]
port 18 nsew signal output
rlabel metal2 s 10136 0 10192 400 6 addr_mem0[8]
port 19 nsew signal output
rlabel metal2 s 38696 0 38752 400 6 addr_mem1[0]
port 20 nsew signal output
rlabel metal2 s 39536 0 39592 400 6 addr_mem1[1]
port 21 nsew signal output
rlabel metal2 s 40376 0 40432 400 6 addr_mem1[2]
port 22 nsew signal output
rlabel metal2 s 41216 0 41272 400 6 addr_mem1[3]
port 23 nsew signal output
rlabel metal2 s 42056 0 42112 400 6 addr_mem1[4]
port 24 nsew signal output
rlabel metal2 s 42896 0 42952 400 6 addr_mem1[5]
port 25 nsew signal output
rlabel metal2 s 43736 0 43792 400 6 addr_mem1[6]
port 26 nsew signal output
rlabel metal2 s 44576 0 44632 400 6 addr_mem1[7]
port 27 nsew signal output
rlabel metal2 s 45416 0 45472 400 6 addr_mem1[8]
port 28 nsew signal output
rlabel metal3 s 74600 560 75000 616 6 csb
port 29 nsew signal input
rlabel metal2 s 2576 0 2632 400 6 csb_mem0
port 30 nsew signal output
rlabel metal2 s 37856 0 37912 400 6 csb_mem1
port 31 nsew signal output
rlabel metal3 s 74600 5488 75000 5544 6 dout[0]
port 32 nsew signal output
rlabel metal3 s 74600 9968 75000 10024 6 dout[10]
port 33 nsew signal output
rlabel metal3 s 74600 10416 75000 10472 6 dout[11]
port 34 nsew signal output
rlabel metal3 s 74600 10864 75000 10920 6 dout[12]
port 35 nsew signal output
rlabel metal3 s 74600 11312 75000 11368 6 dout[13]
port 36 nsew signal output
rlabel metal3 s 74600 11760 75000 11816 6 dout[14]
port 37 nsew signal output
rlabel metal3 s 74600 12208 75000 12264 6 dout[15]
port 38 nsew signal output
rlabel metal3 s 74600 12656 75000 12712 6 dout[16]
port 39 nsew signal output
rlabel metal3 s 74600 13104 75000 13160 6 dout[17]
port 40 nsew signal output
rlabel metal3 s 74600 13552 75000 13608 6 dout[18]
port 41 nsew signal output
rlabel metal3 s 74600 14000 75000 14056 6 dout[19]
port 42 nsew signal output
rlabel metal3 s 74600 5936 75000 5992 6 dout[1]
port 43 nsew signal output
rlabel metal3 s 74600 14448 75000 14504 6 dout[20]
port 44 nsew signal output
rlabel metal3 s 74600 14896 75000 14952 6 dout[21]
port 45 nsew signal output
rlabel metal3 s 74600 15344 75000 15400 6 dout[22]
port 46 nsew signal output
rlabel metal3 s 74600 15792 75000 15848 6 dout[23]
port 47 nsew signal output
rlabel metal3 s 74600 16240 75000 16296 6 dout[24]
port 48 nsew signal output
rlabel metal3 s 74600 16688 75000 16744 6 dout[25]
port 49 nsew signal output
rlabel metal3 s 74600 17136 75000 17192 6 dout[26]
port 50 nsew signal output
rlabel metal3 s 74600 17584 75000 17640 6 dout[27]
port 51 nsew signal output
rlabel metal3 s 74600 18032 75000 18088 6 dout[28]
port 52 nsew signal output
rlabel metal3 s 74600 18480 75000 18536 6 dout[29]
port 53 nsew signal output
rlabel metal3 s 74600 6384 75000 6440 6 dout[2]
port 54 nsew signal output
rlabel metal3 s 74600 18928 75000 18984 6 dout[30]
port 55 nsew signal output
rlabel metal3 s 74600 19376 75000 19432 6 dout[31]
port 56 nsew signal output
rlabel metal3 s 74600 6832 75000 6888 6 dout[3]
port 57 nsew signal output
rlabel metal3 s 74600 7280 75000 7336 6 dout[4]
port 58 nsew signal output
rlabel metal3 s 74600 7728 75000 7784 6 dout[5]
port 59 nsew signal output
rlabel metal3 s 74600 8176 75000 8232 6 dout[6]
port 60 nsew signal output
rlabel metal3 s 74600 8624 75000 8680 6 dout[7]
port 61 nsew signal output
rlabel metal3 s 74600 9072 75000 9128 6 dout[8]
port 62 nsew signal output
rlabel metal3 s 74600 9520 75000 9576 6 dout[9]
port 63 nsew signal output
rlabel metal2 s 10976 0 11032 400 6 dout_mem0[0]
port 64 nsew signal input
rlabel metal2 s 19376 0 19432 400 6 dout_mem0[10]
port 65 nsew signal input
rlabel metal2 s 20216 0 20272 400 6 dout_mem0[11]
port 66 nsew signal input
rlabel metal2 s 21056 0 21112 400 6 dout_mem0[12]
port 67 nsew signal input
rlabel metal2 s 21896 0 21952 400 6 dout_mem0[13]
port 68 nsew signal input
rlabel metal2 s 22736 0 22792 400 6 dout_mem0[14]
port 69 nsew signal input
rlabel metal2 s 23576 0 23632 400 6 dout_mem0[15]
port 70 nsew signal input
rlabel metal2 s 24416 0 24472 400 6 dout_mem0[16]
port 71 nsew signal input
rlabel metal2 s 25256 0 25312 400 6 dout_mem0[17]
port 72 nsew signal input
rlabel metal2 s 26096 0 26152 400 6 dout_mem0[18]
port 73 nsew signal input
rlabel metal2 s 26936 0 26992 400 6 dout_mem0[19]
port 74 nsew signal input
rlabel metal2 s 11816 0 11872 400 6 dout_mem0[1]
port 75 nsew signal input
rlabel metal2 s 27776 0 27832 400 6 dout_mem0[20]
port 76 nsew signal input
rlabel metal2 s 28616 0 28672 400 6 dout_mem0[21]
port 77 nsew signal input
rlabel metal2 s 29456 0 29512 400 6 dout_mem0[22]
port 78 nsew signal input
rlabel metal2 s 30296 0 30352 400 6 dout_mem0[23]
port 79 nsew signal input
rlabel metal2 s 31136 0 31192 400 6 dout_mem0[24]
port 80 nsew signal input
rlabel metal2 s 31976 0 32032 400 6 dout_mem0[25]
port 81 nsew signal input
rlabel metal2 s 32816 0 32872 400 6 dout_mem0[26]
port 82 nsew signal input
rlabel metal2 s 33656 0 33712 400 6 dout_mem0[27]
port 83 nsew signal input
rlabel metal2 s 34496 0 34552 400 6 dout_mem0[28]
port 84 nsew signal input
rlabel metal2 s 35336 0 35392 400 6 dout_mem0[29]
port 85 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 dout_mem0[2]
port 86 nsew signal input
rlabel metal2 s 36176 0 36232 400 6 dout_mem0[30]
port 87 nsew signal input
rlabel metal2 s 37016 0 37072 400 6 dout_mem0[31]
port 88 nsew signal input
rlabel metal2 s 13496 0 13552 400 6 dout_mem0[3]
port 89 nsew signal input
rlabel metal2 s 14336 0 14392 400 6 dout_mem0[4]
port 90 nsew signal input
rlabel metal2 s 15176 0 15232 400 6 dout_mem0[5]
port 91 nsew signal input
rlabel metal2 s 16016 0 16072 400 6 dout_mem0[6]
port 92 nsew signal input
rlabel metal2 s 16856 0 16912 400 6 dout_mem0[7]
port 93 nsew signal input
rlabel metal2 s 17696 0 17752 400 6 dout_mem0[8]
port 94 nsew signal input
rlabel metal2 s 18536 0 18592 400 6 dout_mem0[9]
port 95 nsew signal input
rlabel metal2 s 46256 0 46312 400 6 dout_mem1[0]
port 96 nsew signal input
rlabel metal2 s 54656 0 54712 400 6 dout_mem1[10]
port 97 nsew signal input
rlabel metal2 s 55496 0 55552 400 6 dout_mem1[11]
port 98 nsew signal input
rlabel metal2 s 56336 0 56392 400 6 dout_mem1[12]
port 99 nsew signal input
rlabel metal2 s 57176 0 57232 400 6 dout_mem1[13]
port 100 nsew signal input
rlabel metal2 s 58016 0 58072 400 6 dout_mem1[14]
port 101 nsew signal input
rlabel metal2 s 58856 0 58912 400 6 dout_mem1[15]
port 102 nsew signal input
rlabel metal2 s 59696 0 59752 400 6 dout_mem1[16]
port 103 nsew signal input
rlabel metal2 s 60536 0 60592 400 6 dout_mem1[17]
port 104 nsew signal input
rlabel metal2 s 61376 0 61432 400 6 dout_mem1[18]
port 105 nsew signal input
rlabel metal2 s 62216 0 62272 400 6 dout_mem1[19]
port 106 nsew signal input
rlabel metal2 s 47096 0 47152 400 6 dout_mem1[1]
port 107 nsew signal input
rlabel metal2 s 63056 0 63112 400 6 dout_mem1[20]
port 108 nsew signal input
rlabel metal2 s 63896 0 63952 400 6 dout_mem1[21]
port 109 nsew signal input
rlabel metal2 s 64736 0 64792 400 6 dout_mem1[22]
port 110 nsew signal input
rlabel metal2 s 65576 0 65632 400 6 dout_mem1[23]
port 111 nsew signal input
rlabel metal2 s 66416 0 66472 400 6 dout_mem1[24]
port 112 nsew signal input
rlabel metal2 s 67256 0 67312 400 6 dout_mem1[25]
port 113 nsew signal input
rlabel metal2 s 68096 0 68152 400 6 dout_mem1[26]
port 114 nsew signal input
rlabel metal2 s 68936 0 68992 400 6 dout_mem1[27]
port 115 nsew signal input
rlabel metal2 s 69776 0 69832 400 6 dout_mem1[28]
port 116 nsew signal input
rlabel metal2 s 70616 0 70672 400 6 dout_mem1[29]
port 117 nsew signal input
rlabel metal2 s 47936 0 47992 400 6 dout_mem1[2]
port 118 nsew signal input
rlabel metal2 s 71456 0 71512 400 6 dout_mem1[30]
port 119 nsew signal input
rlabel metal2 s 72296 0 72352 400 6 dout_mem1[31]
port 120 nsew signal input
rlabel metal2 s 48776 0 48832 400 6 dout_mem1[3]
port 121 nsew signal input
rlabel metal2 s 49616 0 49672 400 6 dout_mem1[4]
port 122 nsew signal input
rlabel metal2 s 50456 0 50512 400 6 dout_mem1[5]
port 123 nsew signal input
rlabel metal2 s 51296 0 51352 400 6 dout_mem1[6]
port 124 nsew signal input
rlabel metal2 s 52136 0 52192 400 6 dout_mem1[7]
port 125 nsew signal input
rlabel metal2 s 52976 0 53032 400 6 dout_mem1[8]
port 126 nsew signal input
rlabel metal2 s 53816 0 53872 400 6 dout_mem1[9]
port 127 nsew signal input
rlabel metal4 s 9797 1538 9957 18454 6 vdd
port 128 nsew power bidirectional
rlabel metal4 s 28207 1538 28367 18454 6 vdd
port 128 nsew power bidirectional
rlabel metal4 s 46617 1538 46777 18454 6 vdd
port 128 nsew power bidirectional
rlabel metal4 s 65027 1538 65187 18454 6 vdd
port 128 nsew power bidirectional
rlabel metal4 s 19002 1538 19162 18454 6 vss
port 129 nsew ground bidirectional
rlabel metal4 s 37412 1538 37572 18454 6 vss
port 129 nsew ground bidirectional
rlabel metal4 s 55822 1538 55982 18454 6 vss
port 129 nsew ground bidirectional
rlabel metal4 s 74232 1538 74392 18454 6 vss
port 129 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 75000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 825798
string GDS_FILE /home/leo/Dokumente/the-final-workspace/caravel_user_project/openlane/merge_memory/runs/22_12_05_16_41/results/signoff/merge_memory.magic.gds
string GDS_START 65398
<< end >>

