magic
tech gf180mcuC
magscale 1 10
timestamp 1669805783
<< metal1 >>
rect 1344 36874 148624 36908
rect 1344 36822 19624 36874
rect 19676 36822 19728 36874
rect 19780 36822 19832 36874
rect 19884 36822 56444 36874
rect 56496 36822 56548 36874
rect 56600 36822 56652 36874
rect 56704 36822 93264 36874
rect 93316 36822 93368 36874
rect 93420 36822 93472 36874
rect 93524 36822 130084 36874
rect 130136 36822 130188 36874
rect 130240 36822 130292 36874
rect 130344 36822 148624 36874
rect 1344 36788 148624 36822
rect 145842 36542 145854 36594
rect 145906 36542 145918 36594
rect 144834 36430 144846 36482
rect 144898 36430 144910 36482
rect 146850 36430 146862 36482
rect 146914 36430 146926 36482
rect 147746 36318 147758 36370
rect 147810 36318 147822 36370
rect 143838 36258 143890 36270
rect 143838 36194 143890 36206
rect 144286 36258 144338 36270
rect 144286 36194 144338 36206
rect 1344 36090 148784 36124
rect 1344 36038 38034 36090
rect 38086 36038 38138 36090
rect 38190 36038 38242 36090
rect 38294 36038 74854 36090
rect 74906 36038 74958 36090
rect 75010 36038 75062 36090
rect 75114 36038 111674 36090
rect 111726 36038 111778 36090
rect 111830 36038 111882 36090
rect 111934 36038 148494 36090
rect 148546 36038 148598 36090
rect 148650 36038 148702 36090
rect 148754 36038 148784 36090
rect 1344 36004 148784 36038
rect 145954 35758 145966 35810
rect 146018 35758 146030 35810
rect 145058 35646 145070 35698
rect 145122 35646 145134 35698
rect 146962 35646 146974 35698
rect 147026 35646 147038 35698
rect 144286 35586 144338 35598
rect 147746 35534 147758 35586
rect 147810 35534 147822 35586
rect 144286 35522 144338 35534
rect 1344 35306 148624 35340
rect 1344 35254 19624 35306
rect 19676 35254 19728 35306
rect 19780 35254 19832 35306
rect 19884 35254 56444 35306
rect 56496 35254 56548 35306
rect 56600 35254 56652 35306
rect 56704 35254 93264 35306
rect 93316 35254 93368 35306
rect 93420 35254 93472 35306
rect 93524 35254 130084 35306
rect 130136 35254 130188 35306
rect 130240 35254 130292 35306
rect 130344 35254 148624 35306
rect 1344 35220 148624 35254
rect 146066 34974 146078 35026
rect 146130 34974 146142 35026
rect 145058 34862 145070 34914
rect 145122 34862 145134 34914
rect 146850 34862 146862 34914
rect 146914 34862 146926 34914
rect 147746 34750 147758 34802
rect 147810 34750 147822 34802
rect 144510 34690 144562 34702
rect 144510 34626 144562 34638
rect 1344 34522 148784 34556
rect 1344 34470 38034 34522
rect 38086 34470 38138 34522
rect 38190 34470 38242 34522
rect 38294 34470 74854 34522
rect 74906 34470 74958 34522
rect 75010 34470 75062 34522
rect 75114 34470 111674 34522
rect 111726 34470 111778 34522
rect 111830 34470 111882 34522
rect 111934 34470 148494 34522
rect 148546 34470 148598 34522
rect 148650 34470 148702 34522
rect 148754 34470 148784 34522
rect 1344 34436 148784 34470
rect 146414 34130 146466 34142
rect 147074 34078 147086 34130
rect 147138 34078 147150 34130
rect 146414 34066 146466 34078
rect 145406 34018 145458 34030
rect 145406 33954 145458 33966
rect 145854 34018 145906 34030
rect 147746 33966 147758 34018
rect 147810 33966 147822 34018
rect 145854 33954 145906 33966
rect 1344 33738 148624 33772
rect 1344 33686 19624 33738
rect 19676 33686 19728 33738
rect 19780 33686 19832 33738
rect 19884 33686 56444 33738
rect 56496 33686 56548 33738
rect 56600 33686 56652 33738
rect 56704 33686 93264 33738
rect 93316 33686 93368 33738
rect 93420 33686 93472 33738
rect 93524 33686 130084 33738
rect 130136 33686 130188 33738
rect 130240 33686 130292 33738
rect 130344 33686 148624 33738
rect 1344 33652 148624 33686
rect 146302 33346 146354 33358
rect 146850 33294 146862 33346
rect 146914 33294 146926 33346
rect 146302 33282 146354 33294
rect 147746 33182 147758 33234
rect 147810 33182 147822 33234
rect 1344 32954 148784 32988
rect 1344 32902 38034 32954
rect 38086 32902 38138 32954
rect 38190 32902 38242 32954
rect 38294 32902 74854 32954
rect 74906 32902 74958 32954
rect 75010 32902 75062 32954
rect 75114 32902 111674 32954
rect 111726 32902 111778 32954
rect 111830 32902 111882 32954
rect 111934 32902 148494 32954
rect 148546 32902 148598 32954
rect 148650 32902 148702 32954
rect 148754 32902 148784 32954
rect 1344 32868 148784 32902
rect 1344 32170 148624 32204
rect 1344 32118 19624 32170
rect 19676 32118 19728 32170
rect 19780 32118 19832 32170
rect 19884 32118 56444 32170
rect 56496 32118 56548 32170
rect 56600 32118 56652 32170
rect 56704 32118 93264 32170
rect 93316 32118 93368 32170
rect 93420 32118 93472 32170
rect 93524 32118 130084 32170
rect 130136 32118 130188 32170
rect 130240 32118 130292 32170
rect 130344 32118 148624 32170
rect 1344 32084 148624 32118
rect 146850 31726 146862 31778
rect 146914 31726 146926 31778
rect 147746 31614 147758 31666
rect 147810 31614 147822 31666
rect 146302 31554 146354 31566
rect 146302 31490 146354 31502
rect 1344 31386 148784 31420
rect 1344 31334 38034 31386
rect 38086 31334 38138 31386
rect 38190 31334 38242 31386
rect 38294 31334 74854 31386
rect 74906 31334 74958 31386
rect 75010 31334 75062 31386
rect 75114 31334 111674 31386
rect 111726 31334 111778 31386
rect 111830 31334 111882 31386
rect 111934 31334 148494 31386
rect 148546 31334 148598 31386
rect 148650 31334 148702 31386
rect 148754 31334 148784 31386
rect 1344 31300 148784 31334
rect 146414 30994 146466 31006
rect 146850 30942 146862 30994
rect 146914 30942 146926 30994
rect 146414 30930 146466 30942
rect 147746 30830 147758 30882
rect 147810 30830 147822 30882
rect 1344 30602 148624 30636
rect 1344 30550 19624 30602
rect 19676 30550 19728 30602
rect 19780 30550 19832 30602
rect 19884 30550 56444 30602
rect 56496 30550 56548 30602
rect 56600 30550 56652 30602
rect 56704 30550 93264 30602
rect 93316 30550 93368 30602
rect 93420 30550 93472 30602
rect 93524 30550 130084 30602
rect 130136 30550 130188 30602
rect 130240 30550 130292 30602
rect 130344 30550 148624 30602
rect 1344 30516 148624 30550
rect 146302 30210 146354 30222
rect 147074 30158 147086 30210
rect 147138 30158 147150 30210
rect 146302 30146 146354 30158
rect 147746 30046 147758 30098
rect 147810 30046 147822 30098
rect 1344 29818 148784 29852
rect 1344 29766 38034 29818
rect 38086 29766 38138 29818
rect 38190 29766 38242 29818
rect 38294 29766 74854 29818
rect 74906 29766 74958 29818
rect 75010 29766 75062 29818
rect 75114 29766 111674 29818
rect 111726 29766 111778 29818
rect 111830 29766 111882 29818
rect 111934 29766 148494 29818
rect 148546 29766 148598 29818
rect 148650 29766 148702 29818
rect 148754 29766 148784 29818
rect 1344 29732 148784 29766
rect 146414 29426 146466 29438
rect 146850 29374 146862 29426
rect 146914 29374 146926 29426
rect 146414 29362 146466 29374
rect 147746 29262 147758 29314
rect 147810 29262 147822 29314
rect 1344 29034 148624 29068
rect 1344 28982 19624 29034
rect 19676 28982 19728 29034
rect 19780 28982 19832 29034
rect 19884 28982 56444 29034
rect 56496 28982 56548 29034
rect 56600 28982 56652 29034
rect 56704 28982 93264 29034
rect 93316 28982 93368 29034
rect 93420 28982 93472 29034
rect 93524 28982 130084 29034
rect 130136 28982 130188 29034
rect 130240 28982 130292 29034
rect 130344 28982 148624 29034
rect 1344 28948 148624 28982
rect 146302 28642 146354 28654
rect 146850 28590 146862 28642
rect 146914 28590 146926 28642
rect 147746 28590 147758 28642
rect 147810 28590 147822 28642
rect 146302 28578 146354 28590
rect 1344 28250 148784 28284
rect 1344 28198 38034 28250
rect 38086 28198 38138 28250
rect 38190 28198 38242 28250
rect 38294 28198 74854 28250
rect 74906 28198 74958 28250
rect 75010 28198 75062 28250
rect 75114 28198 111674 28250
rect 111726 28198 111778 28250
rect 111830 28198 111882 28250
rect 111934 28198 148494 28250
rect 148546 28198 148598 28250
rect 148650 28198 148702 28250
rect 148754 28198 148784 28250
rect 1344 28164 148784 28198
rect 146414 27858 146466 27870
rect 147074 27806 147086 27858
rect 147138 27806 147150 27858
rect 146414 27794 146466 27806
rect 147746 27694 147758 27746
rect 147810 27694 147822 27746
rect 1344 27466 148624 27500
rect 1344 27414 19624 27466
rect 19676 27414 19728 27466
rect 19780 27414 19832 27466
rect 19884 27414 56444 27466
rect 56496 27414 56548 27466
rect 56600 27414 56652 27466
rect 56704 27414 93264 27466
rect 93316 27414 93368 27466
rect 93420 27414 93472 27466
rect 93524 27414 130084 27466
rect 130136 27414 130188 27466
rect 130240 27414 130292 27466
rect 130344 27414 148624 27466
rect 1344 27380 148624 27414
rect 146302 27186 146354 27198
rect 146302 27122 146354 27134
rect 146850 27022 146862 27074
rect 146914 27022 146926 27074
rect 147746 26910 147758 26962
rect 147810 26910 147822 26962
rect 1344 26682 148784 26716
rect 1344 26630 38034 26682
rect 38086 26630 38138 26682
rect 38190 26630 38242 26682
rect 38294 26630 74854 26682
rect 74906 26630 74958 26682
rect 75010 26630 75062 26682
rect 75114 26630 111674 26682
rect 111726 26630 111778 26682
rect 111830 26630 111882 26682
rect 111934 26630 148494 26682
rect 148546 26630 148598 26682
rect 148650 26630 148702 26682
rect 148754 26630 148784 26682
rect 1344 26596 148784 26630
rect 1344 25898 148624 25932
rect 1344 25846 19624 25898
rect 19676 25846 19728 25898
rect 19780 25846 19832 25898
rect 19884 25846 56444 25898
rect 56496 25846 56548 25898
rect 56600 25846 56652 25898
rect 56704 25846 93264 25898
rect 93316 25846 93368 25898
rect 93420 25846 93472 25898
rect 93524 25846 130084 25898
rect 130136 25846 130188 25898
rect 130240 25846 130292 25898
rect 130344 25846 148624 25898
rect 1344 25812 148624 25846
rect 146850 25454 146862 25506
rect 146914 25454 146926 25506
rect 147746 25342 147758 25394
rect 147810 25342 147822 25394
rect 146302 25282 146354 25294
rect 146302 25218 146354 25230
rect 1344 25114 148784 25148
rect 1344 25062 38034 25114
rect 38086 25062 38138 25114
rect 38190 25062 38242 25114
rect 38294 25062 74854 25114
rect 74906 25062 74958 25114
rect 75010 25062 75062 25114
rect 75114 25062 111674 25114
rect 111726 25062 111778 25114
rect 111830 25062 111882 25114
rect 111934 25062 148494 25114
rect 148546 25062 148598 25114
rect 148650 25062 148702 25114
rect 148754 25062 148784 25114
rect 1344 25028 148784 25062
rect 146850 24670 146862 24722
rect 146914 24670 146926 24722
rect 146414 24610 146466 24622
rect 147746 24558 147758 24610
rect 147810 24558 147822 24610
rect 146414 24546 146466 24558
rect 1344 24330 148624 24364
rect 1344 24278 19624 24330
rect 19676 24278 19728 24330
rect 19780 24278 19832 24330
rect 19884 24278 56444 24330
rect 56496 24278 56548 24330
rect 56600 24278 56652 24330
rect 56704 24278 93264 24330
rect 93316 24278 93368 24330
rect 93420 24278 93472 24330
rect 93524 24278 130084 24330
rect 130136 24278 130188 24330
rect 130240 24278 130292 24330
rect 130344 24278 148624 24330
rect 1344 24244 148624 24278
rect 146850 23886 146862 23938
rect 146914 23886 146926 23938
rect 147746 23774 147758 23826
rect 147810 23774 147822 23826
rect 146302 23714 146354 23726
rect 146302 23650 146354 23662
rect 1344 23546 148784 23580
rect 1344 23494 38034 23546
rect 38086 23494 38138 23546
rect 38190 23494 38242 23546
rect 38294 23494 74854 23546
rect 74906 23494 74958 23546
rect 75010 23494 75062 23546
rect 75114 23494 111674 23546
rect 111726 23494 111778 23546
rect 111830 23494 111882 23546
rect 111934 23494 148494 23546
rect 148546 23494 148598 23546
rect 148650 23494 148702 23546
rect 148754 23494 148784 23546
rect 1344 23460 148784 23494
rect 146414 23154 146466 23166
rect 146850 23102 146862 23154
rect 146914 23102 146926 23154
rect 146414 23090 146466 23102
rect 147746 22990 147758 23042
rect 147810 22990 147822 23042
rect 1344 22762 148624 22796
rect 1344 22710 19624 22762
rect 19676 22710 19728 22762
rect 19780 22710 19832 22762
rect 19884 22710 56444 22762
rect 56496 22710 56548 22762
rect 56600 22710 56652 22762
rect 56704 22710 93264 22762
rect 93316 22710 93368 22762
rect 93420 22710 93472 22762
rect 93524 22710 130084 22762
rect 130136 22710 130188 22762
rect 130240 22710 130292 22762
rect 130344 22710 148624 22762
rect 1344 22676 148624 22710
rect 146302 22370 146354 22382
rect 146850 22318 146862 22370
rect 146914 22318 146926 22370
rect 146302 22306 146354 22318
rect 147746 22206 147758 22258
rect 147810 22206 147822 22258
rect 1344 21978 148784 22012
rect 1344 21926 38034 21978
rect 38086 21926 38138 21978
rect 38190 21926 38242 21978
rect 38294 21926 74854 21978
rect 74906 21926 74958 21978
rect 75010 21926 75062 21978
rect 75114 21926 111674 21978
rect 111726 21926 111778 21978
rect 111830 21926 111882 21978
rect 111934 21926 148494 21978
rect 148546 21926 148598 21978
rect 148650 21926 148702 21978
rect 148754 21926 148784 21978
rect 1344 21892 148784 21926
rect 146850 21534 146862 21586
rect 146914 21534 146926 21586
rect 146414 21474 146466 21486
rect 147746 21422 147758 21474
rect 147810 21422 147822 21474
rect 146414 21410 146466 21422
rect 1344 21194 148624 21228
rect 1344 21142 19624 21194
rect 19676 21142 19728 21194
rect 19780 21142 19832 21194
rect 19884 21142 56444 21194
rect 56496 21142 56548 21194
rect 56600 21142 56652 21194
rect 56704 21142 93264 21194
rect 93316 21142 93368 21194
rect 93420 21142 93472 21194
rect 93524 21142 130084 21194
rect 130136 21142 130188 21194
rect 130240 21142 130292 21194
rect 130344 21142 148624 21194
rect 1344 21108 148624 21142
rect 146302 20802 146354 20814
rect 146850 20750 146862 20802
rect 146914 20750 146926 20802
rect 146302 20738 146354 20750
rect 147746 20638 147758 20690
rect 147810 20638 147822 20690
rect 1344 20410 148784 20444
rect 1344 20358 38034 20410
rect 38086 20358 38138 20410
rect 38190 20358 38242 20410
rect 38294 20358 74854 20410
rect 74906 20358 74958 20410
rect 75010 20358 75062 20410
rect 75114 20358 111674 20410
rect 111726 20358 111778 20410
rect 111830 20358 111882 20410
rect 111934 20358 148494 20410
rect 148546 20358 148598 20410
rect 148650 20358 148702 20410
rect 148754 20358 148784 20410
rect 1344 20324 148784 20358
rect 1344 19626 148624 19660
rect 1344 19574 19624 19626
rect 19676 19574 19728 19626
rect 19780 19574 19832 19626
rect 19884 19574 56444 19626
rect 56496 19574 56548 19626
rect 56600 19574 56652 19626
rect 56704 19574 93264 19626
rect 93316 19574 93368 19626
rect 93420 19574 93472 19626
rect 93524 19574 130084 19626
rect 130136 19574 130188 19626
rect 130240 19574 130292 19626
rect 130344 19574 148624 19626
rect 1344 19540 148624 19574
rect 146302 19234 146354 19246
rect 146850 19182 146862 19234
rect 146914 19182 146926 19234
rect 146302 19170 146354 19182
rect 147746 19070 147758 19122
rect 147810 19070 147822 19122
rect 1344 18842 148784 18876
rect 1344 18790 38034 18842
rect 38086 18790 38138 18842
rect 38190 18790 38242 18842
rect 38294 18790 74854 18842
rect 74906 18790 74958 18842
rect 75010 18790 75062 18842
rect 75114 18790 111674 18842
rect 111726 18790 111778 18842
rect 111830 18790 111882 18842
rect 111934 18790 148494 18842
rect 148546 18790 148598 18842
rect 148650 18790 148702 18842
rect 148754 18790 148784 18842
rect 1344 18756 148784 18790
rect 114046 18674 114098 18686
rect 114046 18610 114098 18622
rect 113710 18450 113762 18462
rect 146850 18398 146862 18450
rect 146914 18398 146926 18450
rect 113710 18386 113762 18398
rect 113150 18338 113202 18350
rect 113150 18274 113202 18286
rect 146414 18338 146466 18350
rect 147746 18286 147758 18338
rect 147810 18286 147822 18338
rect 146414 18274 146466 18286
rect 1344 18058 148624 18092
rect 1344 18006 19624 18058
rect 19676 18006 19728 18058
rect 19780 18006 19832 18058
rect 19884 18006 56444 18058
rect 56496 18006 56548 18058
rect 56600 18006 56652 18058
rect 56704 18006 93264 18058
rect 93316 18006 93368 18058
rect 93420 18006 93472 18058
rect 93524 18006 130084 18058
rect 130136 18006 130188 18058
rect 130240 18006 130292 18058
rect 130344 18006 148624 18058
rect 1344 17972 148624 18006
rect 146850 17614 146862 17666
rect 146914 17614 146926 17666
rect 147746 17502 147758 17554
rect 147810 17502 147822 17554
rect 146302 17442 146354 17454
rect 146302 17378 146354 17390
rect 1344 17274 148784 17308
rect 1344 17222 38034 17274
rect 38086 17222 38138 17274
rect 38190 17222 38242 17274
rect 38294 17222 74854 17274
rect 74906 17222 74958 17274
rect 75010 17222 75062 17274
rect 75114 17222 111674 17274
rect 111726 17222 111778 17274
rect 111830 17222 111882 17274
rect 111934 17222 148494 17274
rect 148546 17222 148598 17274
rect 148650 17222 148702 17274
rect 148754 17222 148784 17274
rect 1344 17188 148784 17222
rect 146414 16994 146466 17006
rect 146414 16930 146466 16942
rect 146850 16830 146862 16882
rect 146914 16830 146926 16882
rect 147746 16830 147758 16882
rect 147810 16830 147822 16882
rect 1344 16490 148624 16524
rect 1344 16438 19624 16490
rect 19676 16438 19728 16490
rect 19780 16438 19832 16490
rect 19884 16438 56444 16490
rect 56496 16438 56548 16490
rect 56600 16438 56652 16490
rect 56704 16438 93264 16490
rect 93316 16438 93368 16490
rect 93420 16438 93472 16490
rect 93524 16438 130084 16490
rect 130136 16438 130188 16490
rect 130240 16438 130292 16490
rect 130344 16438 148624 16490
rect 1344 16404 148624 16438
rect 146850 16046 146862 16098
rect 146914 16046 146926 16098
rect 147746 15934 147758 15986
rect 147810 15934 147822 15986
rect 146302 15874 146354 15886
rect 146302 15810 146354 15822
rect 1344 15706 148784 15740
rect 1344 15654 38034 15706
rect 38086 15654 38138 15706
rect 38190 15654 38242 15706
rect 38294 15654 74854 15706
rect 74906 15654 74958 15706
rect 75010 15654 75062 15706
rect 75114 15654 111674 15706
rect 111726 15654 111778 15706
rect 111830 15654 111882 15706
rect 111934 15654 148494 15706
rect 148546 15654 148598 15706
rect 148650 15654 148702 15706
rect 148754 15654 148784 15706
rect 1344 15620 148784 15654
rect 146414 15426 146466 15438
rect 146414 15362 146466 15374
rect 146850 15262 146862 15314
rect 146914 15262 146926 15314
rect 147746 15150 147758 15202
rect 147810 15150 147822 15202
rect 1344 14922 148624 14956
rect 1344 14870 19624 14922
rect 19676 14870 19728 14922
rect 19780 14870 19832 14922
rect 19884 14870 56444 14922
rect 56496 14870 56548 14922
rect 56600 14870 56652 14922
rect 56704 14870 93264 14922
rect 93316 14870 93368 14922
rect 93420 14870 93472 14922
rect 93524 14870 130084 14922
rect 130136 14870 130188 14922
rect 130240 14870 130292 14922
rect 130344 14870 148624 14922
rect 1344 14836 148624 14870
rect 146302 14530 146354 14542
rect 146850 14478 146862 14530
rect 146914 14478 146926 14530
rect 146302 14466 146354 14478
rect 147746 14366 147758 14418
rect 147810 14366 147822 14418
rect 1344 14138 148784 14172
rect 1344 14086 38034 14138
rect 38086 14086 38138 14138
rect 38190 14086 38242 14138
rect 38294 14086 74854 14138
rect 74906 14086 74958 14138
rect 75010 14086 75062 14138
rect 75114 14086 111674 14138
rect 111726 14086 111778 14138
rect 111830 14086 111882 14138
rect 111934 14086 148494 14138
rect 148546 14086 148598 14138
rect 148650 14086 148702 14138
rect 148754 14086 148784 14138
rect 1344 14052 148784 14086
rect 1344 13354 148624 13388
rect 1344 13302 19624 13354
rect 19676 13302 19728 13354
rect 19780 13302 19832 13354
rect 19884 13302 56444 13354
rect 56496 13302 56548 13354
rect 56600 13302 56652 13354
rect 56704 13302 93264 13354
rect 93316 13302 93368 13354
rect 93420 13302 93472 13354
rect 93524 13302 130084 13354
rect 130136 13302 130188 13354
rect 130240 13302 130292 13354
rect 130344 13302 148624 13354
rect 1344 13268 148624 13302
rect 146302 12962 146354 12974
rect 146850 12910 146862 12962
rect 146914 12910 146926 12962
rect 146302 12898 146354 12910
rect 101502 12850 101554 12862
rect 101502 12786 101554 12798
rect 101838 12850 101890 12862
rect 147746 12798 147758 12850
rect 147810 12798 147822 12850
rect 101838 12786 101890 12798
rect 1344 12570 148784 12604
rect 1344 12518 38034 12570
rect 38086 12518 38138 12570
rect 38190 12518 38242 12570
rect 38294 12518 74854 12570
rect 74906 12518 74958 12570
rect 75010 12518 75062 12570
rect 75114 12518 111674 12570
rect 111726 12518 111778 12570
rect 111830 12518 111882 12570
rect 111934 12518 148494 12570
rect 148546 12518 148598 12570
rect 148650 12518 148702 12570
rect 148754 12518 148784 12570
rect 1344 12484 148784 12518
rect 100718 12402 100770 12414
rect 100718 12338 100770 12350
rect 100482 12126 100494 12178
rect 100546 12126 100558 12178
rect 146850 12126 146862 12178
rect 146914 12126 146926 12178
rect 101166 12066 101218 12078
rect 101166 12002 101218 12014
rect 146414 12066 146466 12078
rect 147746 12014 147758 12066
rect 147810 12014 147822 12066
rect 146414 12002 146466 12014
rect 1344 11786 148624 11820
rect 1344 11734 19624 11786
rect 19676 11734 19728 11786
rect 19780 11734 19832 11786
rect 19884 11734 56444 11786
rect 56496 11734 56548 11786
rect 56600 11734 56652 11786
rect 56704 11734 93264 11786
rect 93316 11734 93368 11786
rect 93420 11734 93472 11786
rect 93524 11734 130084 11786
rect 130136 11734 130188 11786
rect 130240 11734 130292 11786
rect 130344 11734 148624 11786
rect 1344 11700 148624 11734
rect 146302 11394 146354 11406
rect 146850 11342 146862 11394
rect 146914 11342 146926 11394
rect 146302 11330 146354 11342
rect 99486 11282 99538 11294
rect 99486 11218 99538 11230
rect 99822 11282 99874 11294
rect 147746 11230 147758 11282
rect 147810 11230 147822 11282
rect 99822 11218 99874 11230
rect 1344 11002 148784 11036
rect 1344 10950 38034 11002
rect 38086 10950 38138 11002
rect 38190 10950 38242 11002
rect 38294 10950 74854 11002
rect 74906 10950 74958 11002
rect 75010 10950 75062 11002
rect 75114 10950 111674 11002
rect 111726 10950 111778 11002
rect 111830 10950 111882 11002
rect 111934 10950 148494 11002
rect 148546 10950 148598 11002
rect 148650 10950 148702 11002
rect 148754 10950 148784 11002
rect 1344 10916 148784 10950
rect 147758 10722 147810 10734
rect 147758 10658 147810 10670
rect 148094 10610 148146 10622
rect 148094 10546 148146 10558
rect 147310 10498 147362 10510
rect 147310 10434 147362 10446
rect 1344 10218 148624 10252
rect 1344 10166 19624 10218
rect 19676 10166 19728 10218
rect 19780 10166 19832 10218
rect 19884 10166 56444 10218
rect 56496 10166 56548 10218
rect 56600 10166 56652 10218
rect 56704 10166 93264 10218
rect 93316 10166 93368 10218
rect 93420 10166 93472 10218
rect 93524 10166 130084 10218
rect 130136 10166 130188 10218
rect 130240 10166 130292 10218
rect 130344 10166 148624 10218
rect 1344 10132 148624 10166
rect 148094 9714 148146 9726
rect 148094 9650 148146 9662
rect 147310 9602 147362 9614
rect 147310 9538 147362 9550
rect 147758 9602 147810 9614
rect 147758 9538 147810 9550
rect 1344 9434 148784 9468
rect 1344 9382 38034 9434
rect 38086 9382 38138 9434
rect 38190 9382 38242 9434
rect 38294 9382 74854 9434
rect 74906 9382 74958 9434
rect 75010 9382 75062 9434
rect 75114 9382 111674 9434
rect 111726 9382 111778 9434
rect 111830 9382 111882 9434
rect 111934 9382 148494 9434
rect 148546 9382 148598 9434
rect 148650 9382 148702 9434
rect 148754 9382 148784 9434
rect 1344 9348 148784 9382
rect 147758 9154 147810 9166
rect 147758 9090 147810 9102
rect 147310 9042 147362 9054
rect 147310 8978 147362 8990
rect 148094 9042 148146 9054
rect 148094 8978 148146 8990
rect 1344 8650 148624 8684
rect 1344 8598 19624 8650
rect 19676 8598 19728 8650
rect 19780 8598 19832 8650
rect 19884 8598 56444 8650
rect 56496 8598 56548 8650
rect 56600 8598 56652 8650
rect 56704 8598 93264 8650
rect 93316 8598 93368 8650
rect 93420 8598 93472 8650
rect 93524 8598 130084 8650
rect 130136 8598 130188 8650
rect 130240 8598 130292 8650
rect 130344 8598 148624 8650
rect 1344 8564 148624 8598
rect 134878 8146 134930 8158
rect 134878 8082 134930 8094
rect 135326 8146 135378 8158
rect 135326 8082 135378 8094
rect 148094 8146 148146 8158
rect 148094 8082 148146 8094
rect 134542 8034 134594 8046
rect 134542 7970 134594 7982
rect 147310 8034 147362 8046
rect 147310 7970 147362 7982
rect 147758 8034 147810 8046
rect 147758 7970 147810 7982
rect 1344 7866 148784 7900
rect 1344 7814 38034 7866
rect 38086 7814 38138 7866
rect 38190 7814 38242 7866
rect 38294 7814 74854 7866
rect 74906 7814 74958 7866
rect 75010 7814 75062 7866
rect 75114 7814 111674 7866
rect 111726 7814 111778 7866
rect 111830 7814 111882 7866
rect 111934 7814 148494 7866
rect 148546 7814 148598 7866
rect 148650 7814 148702 7866
rect 148754 7814 148784 7866
rect 1344 7780 148784 7814
rect 99598 7698 99650 7710
rect 99598 7634 99650 7646
rect 113486 7698 113538 7710
rect 113486 7634 113538 7646
rect 113150 7474 113202 7486
rect 99362 7422 99374 7474
rect 99426 7422 99438 7474
rect 113150 7410 113202 7422
rect 1344 7082 148624 7116
rect 1344 7030 19624 7082
rect 19676 7030 19728 7082
rect 19780 7030 19832 7082
rect 19884 7030 56444 7082
rect 56496 7030 56548 7082
rect 56600 7030 56652 7082
rect 56704 7030 93264 7082
rect 93316 7030 93368 7082
rect 93420 7030 93472 7082
rect 93524 7030 130084 7082
rect 130136 7030 130188 7082
rect 130240 7030 130292 7082
rect 130344 7030 148624 7082
rect 1344 6996 148624 7030
rect 129278 6578 129330 6590
rect 129278 6514 129330 6526
rect 147310 6578 147362 6590
rect 147310 6514 147362 6526
rect 148094 6578 148146 6590
rect 148094 6514 148146 6526
rect 103518 6466 103570 6478
rect 103518 6402 103570 6414
rect 111582 6466 111634 6478
rect 111582 6402 111634 6414
rect 128606 6466 128658 6478
rect 128606 6402 128658 6414
rect 130958 6466 131010 6478
rect 130958 6402 131010 6414
rect 140926 6466 140978 6478
rect 140926 6402 140978 6414
rect 141262 6466 141314 6478
rect 141262 6402 141314 6414
rect 147758 6466 147810 6478
rect 147758 6402 147810 6414
rect 1344 6298 148784 6332
rect 1344 6246 38034 6298
rect 38086 6246 38138 6298
rect 38190 6246 38242 6298
rect 38294 6246 74854 6298
rect 74906 6246 74958 6298
rect 75010 6246 75062 6298
rect 75114 6246 111674 6298
rect 111726 6246 111778 6298
rect 111830 6246 111882 6298
rect 111934 6246 148494 6298
rect 148546 6246 148598 6298
rect 148650 6246 148702 6298
rect 148754 6246 148784 6298
rect 1344 6212 148784 6246
rect 84478 6130 84530 6142
rect 84478 6066 84530 6078
rect 88398 6130 88450 6142
rect 88398 6066 88450 6078
rect 105534 6130 105586 6142
rect 105534 6066 105586 6078
rect 112142 6130 112194 6142
rect 112142 6066 112194 6078
rect 131406 6130 131458 6142
rect 131406 6066 131458 6078
rect 140814 6130 140866 6142
rect 140814 6066 140866 6078
rect 141710 6130 141762 6142
rect 141710 6066 141762 6078
rect 142606 6130 142658 6142
rect 142606 6066 142658 6078
rect 130062 6018 130114 6030
rect 130062 5954 130114 5966
rect 147758 6018 147810 6030
rect 147758 5954 147810 5966
rect 103966 5906 104018 5918
rect 103966 5842 104018 5854
rect 104414 5906 104466 5918
rect 104414 5842 104466 5854
rect 105198 5906 105250 5918
rect 105198 5842 105250 5854
rect 111246 5906 111298 5918
rect 129726 5906 129778 5918
rect 111906 5854 111918 5906
rect 111970 5854 111982 5906
rect 111246 5842 111298 5854
rect 129726 5842 129778 5854
rect 131070 5906 131122 5918
rect 131070 5842 131122 5854
rect 140478 5906 140530 5918
rect 140478 5842 140530 5854
rect 141374 5906 141426 5918
rect 141374 5842 141426 5854
rect 142270 5906 142322 5918
rect 142270 5842 142322 5854
rect 148094 5906 148146 5918
rect 148094 5842 148146 5854
rect 82686 5794 82738 5806
rect 82686 5730 82738 5742
rect 83582 5794 83634 5806
rect 83582 5730 83634 5742
rect 99598 5794 99650 5806
rect 99598 5730 99650 5742
rect 102510 5794 102562 5806
rect 102510 5730 102562 5742
rect 102958 5794 103010 5806
rect 110238 5794 110290 5806
rect 113262 5794 113314 5806
rect 103506 5742 103518 5794
rect 103570 5742 103582 5794
rect 110786 5742 110798 5794
rect 110850 5742 110862 5794
rect 102958 5730 103010 5742
rect 110238 5730 110290 5742
rect 113262 5730 113314 5742
rect 114158 5794 114210 5806
rect 114158 5730 114210 5742
rect 115614 5794 115666 5806
rect 115614 5730 115666 5742
rect 116062 5794 116114 5806
rect 116062 5730 116114 5742
rect 117070 5794 117122 5806
rect 117070 5730 117122 5742
rect 117518 5794 117570 5806
rect 117518 5730 117570 5742
rect 117854 5794 117906 5806
rect 117854 5730 117906 5742
rect 118302 5794 118354 5806
rect 118302 5730 118354 5742
rect 119198 5794 119250 5806
rect 119198 5730 119250 5742
rect 123902 5794 123954 5806
rect 123902 5730 123954 5742
rect 127598 5794 127650 5806
rect 127598 5730 127650 5742
rect 128270 5794 128322 5806
rect 128270 5730 128322 5742
rect 129278 5794 129330 5806
rect 129278 5730 129330 5742
rect 130510 5794 130562 5806
rect 130510 5730 130562 5742
rect 131966 5794 132018 5806
rect 131966 5730 132018 5742
rect 132862 5794 132914 5806
rect 132862 5730 132914 5742
rect 133758 5794 133810 5806
rect 133758 5730 133810 5742
rect 138798 5794 138850 5806
rect 138798 5730 138850 5742
rect 139582 5794 139634 5806
rect 139582 5730 139634 5742
rect 139918 5794 139970 5806
rect 139918 5730 139970 5742
rect 143054 5794 143106 5806
rect 143054 5730 143106 5742
rect 143502 5794 143554 5806
rect 143502 5730 143554 5742
rect 147310 5794 147362 5806
rect 147310 5730 147362 5742
rect 1344 5514 148624 5548
rect 1344 5462 19624 5514
rect 19676 5462 19728 5514
rect 19780 5462 19832 5514
rect 19884 5462 56444 5514
rect 56496 5462 56548 5514
rect 56600 5462 56652 5514
rect 56704 5462 93264 5514
rect 93316 5462 93368 5514
rect 93420 5462 93472 5514
rect 93524 5462 130084 5514
rect 130136 5462 130188 5514
rect 130240 5462 130292 5514
rect 130344 5462 148624 5514
rect 1344 5428 148624 5462
rect 104862 5346 104914 5358
rect 104862 5282 104914 5294
rect 142158 5346 142210 5358
rect 142158 5282 142210 5294
rect 77646 5234 77698 5246
rect 77646 5170 77698 5182
rect 88062 5234 88114 5246
rect 88062 5170 88114 5182
rect 90190 5234 90242 5246
rect 90190 5170 90242 5182
rect 103070 5234 103122 5246
rect 103070 5170 103122 5182
rect 109566 5234 109618 5246
rect 109566 5170 109618 5182
rect 115390 5234 115442 5246
rect 115390 5170 115442 5182
rect 134654 5234 134706 5246
rect 134654 5170 134706 5182
rect 75854 5122 75906 5134
rect 75854 5058 75906 5070
rect 78542 5122 78594 5134
rect 78542 5058 78594 5070
rect 79438 5122 79490 5134
rect 83246 5122 83298 5134
rect 82114 5070 82126 5122
rect 82178 5070 82190 5122
rect 79438 5058 79490 5070
rect 83246 5058 83298 5070
rect 84254 5122 84306 5134
rect 84254 5058 84306 5070
rect 87614 5122 87666 5134
rect 87614 5058 87666 5070
rect 98366 5122 98418 5134
rect 98366 5058 98418 5070
rect 99038 5122 99090 5134
rect 99038 5058 99090 5070
rect 102622 5122 102674 5134
rect 102622 5058 102674 5070
rect 104526 5122 104578 5134
rect 104526 5058 104578 5070
rect 111806 5122 111858 5134
rect 111806 5058 111858 5070
rect 117630 5122 117682 5134
rect 117630 5058 117682 5070
rect 122782 5122 122834 5134
rect 122782 5058 122834 5070
rect 127374 5122 127426 5134
rect 127374 5058 127426 5070
rect 136110 5122 136162 5134
rect 136110 5058 136162 5070
rect 140254 5122 140306 5134
rect 140254 5058 140306 5070
rect 141822 5122 141874 5134
rect 141822 5058 141874 5070
rect 146414 5122 146466 5134
rect 146414 5058 146466 5070
rect 147310 5122 147362 5134
rect 147310 5058 147362 5070
rect 80558 5010 80610 5022
rect 80558 4946 80610 4958
rect 80894 5010 80946 5022
rect 80894 4946 80946 4958
rect 82910 5010 82962 5022
rect 82910 4946 82962 4958
rect 83918 5010 83970 5022
rect 83918 4946 83970 4958
rect 85598 5010 85650 5022
rect 85598 4946 85650 4958
rect 85934 5010 85986 5022
rect 85934 4946 85986 4958
rect 87278 5010 87330 5022
rect 87278 4946 87330 4958
rect 88958 5010 89010 5022
rect 88958 4946 89010 4958
rect 89294 5010 89346 5022
rect 89294 4946 89346 4958
rect 99486 5010 99538 5022
rect 99486 4946 99538 4958
rect 100382 5010 100434 5022
rect 100382 4946 100434 4958
rect 102062 5010 102114 5022
rect 105534 5010 105586 5022
rect 103730 4958 103742 5010
rect 103794 4958 103806 5010
rect 104178 4958 104190 5010
rect 104242 4958 104254 5010
rect 102062 4946 102114 4958
rect 105534 4946 105586 4958
rect 105870 5010 105922 5022
rect 105870 4946 105922 4958
rect 106430 5010 106482 5022
rect 106430 4946 106482 4958
rect 106766 5010 106818 5022
rect 106766 4946 106818 4958
rect 110014 5010 110066 5022
rect 110014 4946 110066 4958
rect 110350 5010 110402 5022
rect 112142 5010 112194 5022
rect 111010 4958 111022 5010
rect 111074 4958 111086 5010
rect 111458 4958 111470 5010
rect 111522 4958 111534 5010
rect 110350 4946 110402 4958
rect 112142 4946 112194 4958
rect 112814 5010 112866 5022
rect 112814 4946 112866 4958
rect 113150 5010 113202 5022
rect 113150 4946 113202 4958
rect 114606 5010 114658 5022
rect 114606 4946 114658 4958
rect 115950 5010 116002 5022
rect 115950 4946 116002 4958
rect 116286 5010 116338 5022
rect 116286 4946 116338 4958
rect 117070 5010 117122 5022
rect 117070 4946 117122 4958
rect 118190 5010 118242 5022
rect 118190 4946 118242 4958
rect 118526 5010 118578 5022
rect 118526 4946 118578 4958
rect 119086 5010 119138 5022
rect 119086 4946 119138 4958
rect 119422 5010 119474 5022
rect 119422 4946 119474 4958
rect 119982 5010 120034 5022
rect 119982 4946 120034 4958
rect 120318 5010 120370 5022
rect 120318 4946 120370 4958
rect 123566 5010 123618 5022
rect 123566 4946 123618 4958
rect 123902 5010 123954 5022
rect 123902 4946 123954 4958
rect 125022 5010 125074 5022
rect 125022 4946 125074 4958
rect 125358 5010 125410 5022
rect 125358 4946 125410 4958
rect 125918 5010 125970 5022
rect 125918 4946 125970 4958
rect 126254 5010 126306 5022
rect 126254 4946 126306 4958
rect 127038 5010 127090 5022
rect 127038 4946 127090 4958
rect 127934 5010 127986 5022
rect 127934 4946 127986 4958
rect 128270 5010 128322 5022
rect 128270 4946 128322 4958
rect 129054 5010 129106 5022
rect 129054 4946 129106 4958
rect 130174 5010 130226 5022
rect 130174 4946 130226 4958
rect 131070 5010 131122 5022
rect 131070 4946 131122 4958
rect 132974 5010 133026 5022
rect 132974 4946 133026 4958
rect 133310 5010 133362 5022
rect 133310 4946 133362 4958
rect 133870 5010 133922 5022
rect 133870 4946 133922 4958
rect 134206 5010 134258 5022
rect 134206 4946 134258 4958
rect 135550 5010 135602 5022
rect 135550 4946 135602 4958
rect 137454 5010 137506 5022
rect 137454 4946 137506 4958
rect 137790 5010 137842 5022
rect 137790 4946 137842 4958
rect 139134 5010 139186 5022
rect 139134 4946 139186 4958
rect 139470 5010 139522 5022
rect 142830 5010 142882 5022
rect 141138 4958 141150 5010
rect 141202 4958 141214 5010
rect 141586 4958 141598 5010
rect 141650 4958 141662 5010
rect 139470 4946 139522 4958
rect 142830 4946 142882 4958
rect 143166 5010 143218 5022
rect 143166 4946 143218 4958
rect 143726 5010 143778 5022
rect 143726 4946 143778 4958
rect 144062 5010 144114 5022
rect 144062 4946 144114 4958
rect 148094 5010 148146 5022
rect 148094 4946 148146 4958
rect 81342 4898 81394 4910
rect 81342 4834 81394 4846
rect 82350 4898 82402 4910
rect 82350 4834 82402 4846
rect 86382 4898 86434 4910
rect 86382 4834 86434 4846
rect 89742 4898 89794 4910
rect 89742 4834 89794 4846
rect 98030 4898 98082 4910
rect 98030 4834 98082 4846
rect 99822 4898 99874 4910
rect 99822 4834 99874 4846
rect 101166 4898 101218 4910
rect 101166 4834 101218 4846
rect 101614 4898 101666 4910
rect 101614 4834 101666 4846
rect 113598 4898 113650 4910
rect 113598 4834 113650 4846
rect 114158 4898 114210 4910
rect 114158 4834 114210 4846
rect 114942 4898 114994 4910
rect 114942 4834 114994 4846
rect 121102 4898 121154 4910
rect 121102 4834 121154 4846
rect 129614 4898 129666 4910
rect 129614 4834 129666 4846
rect 130510 4898 130562 4910
rect 130510 4834 130562 4846
rect 131630 4898 131682 4910
rect 131630 4834 131682 4846
rect 132078 4898 132130 4910
rect 132078 4834 132130 4846
rect 135102 4898 135154 4910
rect 135102 4834 135154 4846
rect 136782 4898 136834 4910
rect 136782 4834 136834 4846
rect 138686 4898 138738 4910
rect 138686 4834 138738 4846
rect 146862 4898 146914 4910
rect 146862 4834 146914 4846
rect 147758 4898 147810 4910
rect 147758 4834 147810 4846
rect 1344 4730 148784 4764
rect 1344 4678 38034 4730
rect 38086 4678 38138 4730
rect 38190 4678 38242 4730
rect 38294 4678 74854 4730
rect 74906 4678 74958 4730
rect 75010 4678 75062 4730
rect 75114 4678 111674 4730
rect 111726 4678 111778 4730
rect 111830 4678 111882 4730
rect 111934 4678 148494 4730
rect 148546 4678 148598 4730
rect 148650 4678 148702 4730
rect 148754 4678 148784 4730
rect 1344 4644 148784 4678
rect 9774 4562 9826 4574
rect 9774 4498 9826 4510
rect 11342 4562 11394 4574
rect 11342 4498 11394 4510
rect 13022 4562 13074 4574
rect 13022 4498 13074 4510
rect 15150 4562 15202 4574
rect 15150 4498 15202 4510
rect 22542 4562 22594 4574
rect 22542 4498 22594 4510
rect 76078 4562 76130 4574
rect 76078 4498 76130 4510
rect 77870 4562 77922 4574
rect 77870 4498 77922 4510
rect 79662 4562 79714 4574
rect 79662 4498 79714 4510
rect 82126 4562 82178 4574
rect 82126 4498 82178 4510
rect 85374 4562 85426 4574
rect 85374 4498 85426 4510
rect 99486 4562 99538 4574
rect 99486 4498 99538 4510
rect 101390 4562 101442 4574
rect 101390 4498 101442 4510
rect 104302 4562 104354 4574
rect 104302 4498 104354 4510
rect 106430 4562 106482 4574
rect 106430 4498 106482 4510
rect 106990 4562 107042 4574
rect 106990 4498 107042 4510
rect 109006 4562 109058 4574
rect 109006 4498 109058 4510
rect 111582 4562 111634 4574
rect 111582 4498 111634 4510
rect 112142 4562 112194 4574
rect 112142 4498 112194 4510
rect 113262 4562 113314 4574
rect 113262 4498 113314 4510
rect 114942 4562 114994 4574
rect 114942 4498 114994 4510
rect 117070 4562 117122 4574
rect 117070 4498 117122 4510
rect 118974 4562 119026 4574
rect 118974 4498 119026 4510
rect 121438 4562 121490 4574
rect 121438 4498 121490 4510
rect 123230 4562 123282 4574
rect 123230 4498 123282 4510
rect 125358 4562 125410 4574
rect 125358 4498 125410 4510
rect 127262 4562 127314 4574
rect 127262 4498 127314 4510
rect 130734 4562 130786 4574
rect 130734 4498 130786 4510
rect 132862 4562 132914 4574
rect 132862 4498 132914 4510
rect 134094 4562 134146 4574
rect 134094 4498 134146 4510
rect 135662 4562 135714 4574
rect 135662 4498 135714 4510
rect 138238 4562 138290 4574
rect 138238 4498 138290 4510
rect 140254 4562 140306 4574
rect 140254 4498 140306 4510
rect 142158 4562 142210 4574
rect 142158 4498 142210 4510
rect 143726 4562 143778 4574
rect 143726 4498 143778 4510
rect 147758 4562 147810 4574
rect 147758 4498 147810 4510
rect 19406 4450 19458 4462
rect 19406 4386 19458 4398
rect 73950 4450 74002 4462
rect 73950 4386 74002 4398
rect 75294 4450 75346 4462
rect 75294 4386 75346 4398
rect 75630 4450 75682 4462
rect 75630 4386 75682 4398
rect 76974 4450 77026 4462
rect 76974 4386 77026 4398
rect 77310 4450 77362 4462
rect 77310 4386 77362 4398
rect 78206 4450 78258 4462
rect 78206 4386 78258 4398
rect 79102 4450 79154 4462
rect 79102 4386 79154 4398
rect 79998 4450 80050 4462
rect 79998 4386 80050 4398
rect 80446 4450 80498 4462
rect 80446 4386 80498 4398
rect 81342 4450 81394 4462
rect 81342 4386 81394 4398
rect 81678 4450 81730 4462
rect 81678 4386 81730 4398
rect 84814 4450 84866 4462
rect 84814 4386 84866 4398
rect 88174 4450 88226 4462
rect 88174 4386 88226 4398
rect 89630 4450 89682 4462
rect 89630 4386 89682 4398
rect 90750 4450 90802 4462
rect 90750 4386 90802 4398
rect 91310 4450 91362 4462
rect 91310 4386 91362 4398
rect 97694 4450 97746 4462
rect 109790 4450 109842 4462
rect 119982 4450 120034 4462
rect 128270 4450 128322 4462
rect 133534 4450 133586 4462
rect 98466 4398 98478 4450
rect 98530 4398 98542 4450
rect 100370 4398 100382 4450
rect 100434 4398 100446 4450
rect 102162 4398 102174 4450
rect 102226 4398 102238 4450
rect 102722 4398 102734 4450
rect 102786 4398 102798 4450
rect 105522 4398 105534 4450
rect 105586 4398 105598 4450
rect 110562 4398 110574 4450
rect 110626 4398 110638 4450
rect 114258 4398 114270 4450
rect 114322 4398 114334 4450
rect 115938 4398 115950 4450
rect 116002 4398 116014 4450
rect 116498 4398 116510 4450
rect 116562 4398 116574 4450
rect 117842 4398 117854 4450
rect 117906 4398 117918 4450
rect 118402 4398 118414 4450
rect 118466 4398 118478 4450
rect 122098 4398 122110 4450
rect 122162 4398 122174 4450
rect 122658 4398 122670 4450
rect 122722 4398 122734 4450
rect 124338 4398 124350 4450
rect 124402 4398 124414 4450
rect 124786 4398 124798 4450
rect 124850 4398 124862 4450
rect 126354 4398 126366 4450
rect 126418 4398 126430 4450
rect 126690 4398 126702 4450
rect 126754 4398 126766 4450
rect 129826 4398 129838 4450
rect 129890 4398 129902 4450
rect 131842 4398 131854 4450
rect 131906 4398 131918 4450
rect 97694 4386 97746 4398
rect 109790 4386 109842 4398
rect 119982 4386 120034 4398
rect 128270 4386 128322 4398
rect 133534 4386 133586 4398
rect 135102 4450 135154 4462
rect 143166 4450 143218 4462
rect 137218 4398 137230 4450
rect 137282 4398 137294 4450
rect 139122 4398 139134 4450
rect 139186 4398 139198 4450
rect 139570 4398 139582 4450
rect 139634 4398 139646 4450
rect 141138 4398 141150 4450
rect 141202 4398 141214 4450
rect 141586 4398 141598 4450
rect 141650 4398 141662 4450
rect 135102 4386 135154 4398
rect 143166 4386 143218 4398
rect 146862 4450 146914 4462
rect 146862 4386 146914 4398
rect 8878 4338 8930 4350
rect 22206 4338 22258 4350
rect 97358 4338 97410 4350
rect 101054 4338 101106 4350
rect 8306 4286 8318 4338
rect 8370 4286 8382 4338
rect 18946 4286 18958 4338
rect 19010 4286 19022 4338
rect 78866 4286 78878 4338
rect 78930 4286 78942 4338
rect 82674 4286 82686 4338
rect 82738 4286 82750 4338
rect 84578 4286 84590 4338
rect 84642 4286 84654 4338
rect 86146 4286 86158 4338
rect 86210 4286 86222 4338
rect 87938 4286 87950 4338
rect 88002 4286 88014 4338
rect 89394 4286 89406 4338
rect 89458 4286 89470 4338
rect 90514 4286 90526 4338
rect 90578 4286 90590 4338
rect 98690 4286 98702 4338
rect 98754 4286 98766 4338
rect 100594 4286 100606 4338
rect 100658 4286 100670 4338
rect 8878 4274 8930 4286
rect 22206 4274 22258 4286
rect 97358 4274 97410 4286
rect 101054 4274 101106 4286
rect 103294 4338 103346 4350
rect 103294 4274 103346 4286
rect 103966 4338 104018 4350
rect 109454 4338 109506 4350
rect 119646 4338 119698 4350
rect 105298 4286 105310 4338
rect 105362 4286 105374 4338
rect 110450 4286 110462 4338
rect 110514 4286 110526 4338
rect 114034 4286 114046 4338
rect 114098 4286 114110 4338
rect 103966 4274 104018 4286
rect 109454 4274 109506 4286
rect 119646 4274 119698 4286
rect 120990 4338 121042 4350
rect 120990 4274 121042 4286
rect 127934 4338 127986 4350
rect 130398 4338 130450 4350
rect 134766 4338 134818 4350
rect 142830 4338 142882 4350
rect 129602 4286 129614 4338
rect 129666 4286 129678 4338
rect 131730 4286 131742 4338
rect 131794 4286 131806 4338
rect 137106 4286 137118 4338
rect 137170 4286 137182 4338
rect 127934 4274 127986 4286
rect 130398 4274 130450 4286
rect 134766 4274 134818 4286
rect 142830 4274 142882 4286
rect 144062 4338 144114 4350
rect 144062 4274 144114 4286
rect 145294 4338 145346 4350
rect 148094 4338 148146 4350
rect 147074 4286 147086 4338
rect 147138 4286 147150 4338
rect 145294 4274 145346 4286
rect 148094 4274 148146 4286
rect 6638 4226 6690 4238
rect 21758 4226 21810 4238
rect 7298 4174 7310 4226
rect 7362 4174 7374 4226
rect 17938 4174 17950 4226
rect 18002 4174 18014 4226
rect 6638 4162 6690 4174
rect 21758 4162 21810 4174
rect 22990 4226 23042 4238
rect 22990 4162 23042 4174
rect 25566 4226 25618 4238
rect 25566 4162 25618 4174
rect 32622 4226 32674 4238
rect 32622 4162 32674 4174
rect 37102 4226 37154 4238
rect 37102 4162 37154 4174
rect 44382 4226 44434 4238
rect 44382 4162 44434 4174
rect 48862 4226 48914 4238
rect 48862 4162 48914 4174
rect 56142 4226 56194 4238
rect 56142 4162 56194 4174
rect 60622 4226 60674 4238
rect 60622 4162 60674 4174
rect 67902 4226 67954 4238
rect 67902 4162 67954 4174
rect 73278 4226 73330 4238
rect 73278 4162 73330 4174
rect 74398 4226 74450 4238
rect 93550 4226 93602 4238
rect 83346 4174 83358 4226
rect 83410 4174 83422 4226
rect 86706 4174 86718 4226
rect 86770 4174 86782 4226
rect 74398 4162 74450 4174
rect 93550 4162 93602 4174
rect 94446 4226 94498 4238
rect 94446 4162 94498 4174
rect 95902 4226 95954 4238
rect 95902 4162 95954 4174
rect 107438 4226 107490 4238
rect 107438 4162 107490 4174
rect 107886 4226 107938 4238
rect 107886 4162 107938 4174
rect 108558 4226 108610 4238
rect 108558 4162 108610 4174
rect 128942 4226 128994 4238
rect 144846 4226 144898 4238
rect 136098 4174 136110 4226
rect 136162 4174 136174 4226
rect 128942 4162 128994 4174
rect 144846 4162 144898 4174
rect 145966 4226 146018 4238
rect 145966 4162 146018 4174
rect 146414 4226 146466 4238
rect 146414 4162 146466 4174
rect 99150 4114 99202 4126
rect 99150 4050 99202 4062
rect 102958 4114 103010 4126
rect 102958 4050 103010 4062
rect 106094 4114 106146 4126
rect 106094 4050 106146 4062
rect 111246 4114 111298 4126
rect 111246 4050 111298 4062
rect 113598 4114 113650 4126
rect 113598 4050 113650 4062
rect 116734 4114 116786 4126
rect 116734 4050 116786 4062
rect 118638 4114 118690 4126
rect 118638 4050 118690 4062
rect 122894 4114 122946 4126
rect 122894 4050 122946 4062
rect 125022 4114 125074 4126
rect 125022 4050 125074 4062
rect 126926 4114 126978 4126
rect 126926 4050 126978 4062
rect 132526 4114 132578 4126
rect 132526 4050 132578 4062
rect 137902 4114 137954 4126
rect 137902 4050 137954 4062
rect 139918 4114 139970 4126
rect 139918 4050 139970 4062
rect 141822 4114 141874 4126
rect 141822 4050 141874 4062
rect 1344 3946 148624 3980
rect 1344 3894 19624 3946
rect 19676 3894 19728 3946
rect 19780 3894 19832 3946
rect 19884 3894 56444 3946
rect 56496 3894 56548 3946
rect 56600 3894 56652 3946
rect 56704 3894 93264 3946
rect 93316 3894 93368 3946
rect 93420 3894 93472 3946
rect 93524 3894 130084 3946
rect 130136 3894 130188 3946
rect 130240 3894 130292 3946
rect 130344 3894 148624 3946
rect 1344 3860 148624 3894
rect 98926 3778 98978 3790
rect 98926 3714 98978 3726
rect 100718 3778 100770 3790
rect 100718 3714 100770 3726
rect 101054 3778 101106 3790
rect 101054 3714 101106 3726
rect 104974 3778 105026 3790
rect 104974 3714 105026 3726
rect 110574 3778 110626 3790
rect 110574 3714 110626 3726
rect 112478 3778 112530 3790
rect 112478 3714 112530 3726
rect 112814 3778 112866 3790
rect 112814 3714 112866 3726
rect 115614 3778 115666 3790
rect 115614 3714 115666 3726
rect 115950 3778 116002 3790
rect 115950 3714 116002 3726
rect 120318 3778 120370 3790
rect 120318 3714 120370 3726
rect 120654 3778 120706 3790
rect 120654 3714 120706 3726
rect 124574 3778 124626 3790
rect 124574 3714 124626 3726
rect 129726 3778 129778 3790
rect 129726 3714 129778 3726
rect 130062 3778 130114 3790
rect 130062 3714 130114 3726
rect 132414 3778 132466 3790
rect 132414 3714 132466 3726
rect 136334 3778 136386 3790
rect 136334 3714 136386 3726
rect 136670 3778 136722 3790
rect 136670 3714 136722 3726
rect 140254 3778 140306 3790
rect 140254 3714 140306 3726
rect 143838 3778 143890 3790
rect 143838 3714 143890 3726
rect 144174 3778 144226 3790
rect 144174 3714 144226 3726
rect 17502 3666 17554 3678
rect 86942 3666 86994 3678
rect 97134 3666 97186 3678
rect 8194 3614 8206 3666
rect 8258 3614 8270 3666
rect 10210 3614 10222 3666
rect 10274 3614 10286 3666
rect 13906 3614 13918 3666
rect 13970 3614 13982 3666
rect 78754 3614 78766 3666
rect 78818 3614 78830 3666
rect 82674 3614 82686 3666
rect 82738 3614 82750 3666
rect 90514 3614 90526 3666
rect 90578 3614 90590 3666
rect 17502 3602 17554 3614
rect 86942 3602 86994 3614
rect 97134 3602 97186 3614
rect 126030 3666 126082 3678
rect 126030 3602 126082 3614
rect 126590 3666 126642 3678
rect 126590 3602 126642 3614
rect 20638 3554 20690 3566
rect 73726 3554 73778 3566
rect 6738 3502 6750 3554
rect 6802 3502 6814 3554
rect 8866 3502 8878 3554
rect 8930 3502 8942 3554
rect 10994 3502 11006 3554
rect 11058 3502 11070 3554
rect 12786 3502 12798 3554
rect 12850 3502 12862 3554
rect 14914 3502 14926 3554
rect 14978 3502 14990 3554
rect 16706 3502 16718 3554
rect 16770 3502 16782 3554
rect 20066 3502 20078 3554
rect 20130 3502 20142 3554
rect 22642 3502 22654 3554
rect 22706 3502 22718 3554
rect 20638 3490 20690 3502
rect 73726 3490 73778 3502
rect 75518 3554 75570 3566
rect 86494 3554 86546 3566
rect 93774 3554 93826 3566
rect 76290 3502 76302 3554
rect 76354 3502 76366 3554
rect 78082 3502 78094 3554
rect 78146 3502 78158 3554
rect 80210 3502 80222 3554
rect 80274 3502 80286 3554
rect 82002 3502 82014 3554
rect 82066 3502 82078 3554
rect 85362 3502 85374 3554
rect 85426 3502 85438 3554
rect 88162 3502 88174 3554
rect 88226 3502 88238 3554
rect 89842 3502 89854 3554
rect 89906 3502 89918 3554
rect 91970 3502 91982 3554
rect 92034 3502 92046 3554
rect 75518 3490 75570 3502
rect 86494 3490 86546 3502
rect 93774 3490 93826 3502
rect 98590 3554 98642 3566
rect 104638 3554 104690 3566
rect 110238 3554 110290 3566
rect 124238 3554 124290 3566
rect 132078 3554 132130 3566
rect 139918 3554 139970 3566
rect 145630 3554 145682 3566
rect 104178 3502 104190 3554
rect 104242 3502 104254 3554
rect 106754 3502 106766 3554
rect 106818 3502 106830 3554
rect 111794 3502 111806 3554
rect 111858 3502 111870 3554
rect 114594 3502 114606 3554
rect 114658 3502 114670 3554
rect 116722 3502 116734 3554
rect 116786 3502 116798 3554
rect 119634 3502 119646 3554
rect 119698 3502 119710 3554
rect 127474 3502 127486 3554
rect 127538 3502 127550 3554
rect 131394 3502 131406 3554
rect 131458 3502 131470 3554
rect 134194 3502 134206 3554
rect 134258 3502 134270 3554
rect 141138 3502 141150 3554
rect 141202 3502 141214 3554
rect 145058 3502 145070 3554
rect 145122 3502 145134 3554
rect 98590 3490 98642 3502
rect 104638 3490 104690 3502
rect 110238 3490 110290 3502
rect 124238 3490 124290 3502
rect 132078 3490 132130 3502
rect 139918 3490 139970 3502
rect 145630 3490 145682 3502
rect 23438 3442 23490 3454
rect 6066 3390 6078 3442
rect 6130 3390 6142 3442
rect 11890 3390 11902 3442
rect 11954 3390 11966 3442
rect 15810 3390 15822 3442
rect 15874 3390 15886 3442
rect 19170 3390 19182 3442
rect 19234 3390 19246 3442
rect 21746 3390 21758 3442
rect 21810 3390 21822 3442
rect 23438 3378 23490 3390
rect 23886 3442 23938 3454
rect 23886 3378 23938 3390
rect 25566 3442 25618 3454
rect 25566 3378 25618 3390
rect 26798 3442 26850 3454
rect 26798 3378 26850 3390
rect 27246 3442 27298 3454
rect 27246 3378 27298 3390
rect 28590 3442 28642 3454
rect 28590 3378 28642 3390
rect 29262 3442 29314 3454
rect 29262 3378 29314 3390
rect 30158 3442 30210 3454
rect 30158 3378 30210 3390
rect 30606 3442 30658 3454
rect 30606 3378 30658 3390
rect 32062 3442 32114 3454
rect 32062 3378 32114 3390
rect 33518 3442 33570 3454
rect 33518 3378 33570 3390
rect 33966 3442 34018 3454
rect 33966 3378 34018 3390
rect 35198 3442 35250 3454
rect 35198 3378 35250 3390
rect 35646 3442 35698 3454
rect 35646 3378 35698 3390
rect 37326 3442 37378 3454
rect 37326 3378 37378 3390
rect 38558 3442 38610 3454
rect 38558 3378 38610 3390
rect 39006 3442 39058 3454
rect 39006 3378 39058 3390
rect 40350 3442 40402 3454
rect 40350 3378 40402 3390
rect 41022 3442 41074 3454
rect 41022 3378 41074 3390
rect 41918 3442 41970 3454
rect 41918 3378 41970 3390
rect 42366 3442 42418 3454
rect 42366 3378 42418 3390
rect 43822 3442 43874 3454
rect 43822 3378 43874 3390
rect 45278 3442 45330 3454
rect 45278 3378 45330 3390
rect 45726 3442 45778 3454
rect 45726 3378 45778 3390
rect 46958 3442 47010 3454
rect 46958 3378 47010 3390
rect 47406 3442 47458 3454
rect 47406 3378 47458 3390
rect 49086 3442 49138 3454
rect 49086 3378 49138 3390
rect 50318 3442 50370 3454
rect 50318 3378 50370 3390
rect 50766 3442 50818 3454
rect 50766 3378 50818 3390
rect 52110 3442 52162 3454
rect 52110 3378 52162 3390
rect 52782 3442 52834 3454
rect 52782 3378 52834 3390
rect 53678 3442 53730 3454
rect 53678 3378 53730 3390
rect 54126 3442 54178 3454
rect 54126 3378 54178 3390
rect 55582 3442 55634 3454
rect 55582 3378 55634 3390
rect 57038 3442 57090 3454
rect 57038 3378 57090 3390
rect 57486 3442 57538 3454
rect 57486 3378 57538 3390
rect 58718 3442 58770 3454
rect 58718 3378 58770 3390
rect 59166 3442 59218 3454
rect 59166 3378 59218 3390
rect 60846 3442 60898 3454
rect 60846 3378 60898 3390
rect 62078 3442 62130 3454
rect 62078 3378 62130 3390
rect 62526 3442 62578 3454
rect 62526 3378 62578 3390
rect 63870 3442 63922 3454
rect 63870 3378 63922 3390
rect 64542 3442 64594 3454
rect 64542 3378 64594 3390
rect 65438 3442 65490 3454
rect 65438 3378 65490 3390
rect 65886 3442 65938 3454
rect 65886 3378 65938 3390
rect 67342 3442 67394 3454
rect 67342 3378 67394 3390
rect 68798 3442 68850 3454
rect 68798 3378 68850 3390
rect 69246 3442 69298 3454
rect 69246 3378 69298 3390
rect 70478 3442 70530 3454
rect 70478 3378 70530 3390
rect 70926 3442 70978 3454
rect 70926 3378 70978 3390
rect 72494 3442 72546 3454
rect 72494 3378 72546 3390
rect 74286 3442 74338 3454
rect 86158 3442 86210 3454
rect 94670 3442 94722 3454
rect 77186 3390 77198 3442
rect 77250 3390 77262 3442
rect 81106 3390 81118 3442
rect 81170 3390 81182 3442
rect 84690 3390 84702 3442
rect 84754 3390 84766 3442
rect 88946 3390 88958 3442
rect 89010 3390 89022 3442
rect 92866 3390 92878 3442
rect 92930 3390 92942 3442
rect 74286 3378 74338 3390
rect 86158 3378 86210 3390
rect 94670 3378 94722 3390
rect 96126 3442 96178 3454
rect 101726 3442 101778 3454
rect 97794 3390 97806 3442
rect 97858 3390 97870 3442
rect 98354 3390 98366 3442
rect 98418 3390 98430 3442
rect 99922 3390 99934 3442
rect 99986 3390 99998 3442
rect 100482 3390 100494 3442
rect 100546 3390 100558 3442
rect 96126 3378 96178 3390
rect 101726 3378 101778 3390
rect 102622 3442 102674 3454
rect 105982 3442 106034 3454
rect 104066 3390 104078 3442
rect 104130 3390 104142 3442
rect 102622 3378 102674 3390
rect 105982 3378 106034 3390
rect 106542 3442 106594 3454
rect 106542 3378 106594 3390
rect 107886 3442 107938 3454
rect 107886 3378 107938 3390
rect 108670 3442 108722 3454
rect 113822 3442 113874 3454
rect 117742 3442 117794 3454
rect 109442 3390 109454 3442
rect 109506 3390 109518 3442
rect 110002 3390 110014 3442
rect 110066 3390 110078 3442
rect 111682 3390 111694 3442
rect 111746 3390 111758 3442
rect 116498 3390 116510 3442
rect 116562 3390 116574 3442
rect 108670 3378 108722 3390
rect 113822 3378 113874 3390
rect 117742 3378 117794 3390
rect 118302 3442 118354 3454
rect 118302 3378 118354 3390
rect 118638 3442 118690 3454
rect 121326 3442 121378 3454
rect 119522 3390 119534 3442
rect 119586 3390 119598 3442
rect 118638 3378 118690 3390
rect 121326 3378 121378 3390
rect 122222 3442 122274 3454
rect 125246 3442 125298 3454
rect 123666 3390 123678 3442
rect 123730 3390 123742 3442
rect 124002 3390 124014 3442
rect 124066 3390 124078 3442
rect 122222 3378 122274 3390
rect 125246 3378 125298 3390
rect 125582 3442 125634 3454
rect 125582 3378 125634 3390
rect 127262 3442 127314 3454
rect 127262 3378 127314 3390
rect 128046 3442 128098 3454
rect 133422 3442 133474 3454
rect 137342 3442 137394 3454
rect 128930 3390 128942 3442
rect 128994 3390 129006 3442
rect 129378 3390 129390 3442
rect 129442 3390 129454 3442
rect 131282 3390 131294 3442
rect 131346 3390 131358 3442
rect 135538 3390 135550 3442
rect 135602 3390 135614 3442
rect 136098 3390 136110 3442
rect 136162 3390 136174 3442
rect 128046 3378 128098 3390
rect 133422 3378 133474 3390
rect 137342 3378 137394 3390
rect 138126 3442 138178 3454
rect 142158 3442 142210 3454
rect 146078 3442 146130 3454
rect 139346 3390 139358 3442
rect 139410 3390 139422 3442
rect 139570 3390 139582 3442
rect 139634 3390 139646 3442
rect 143266 3390 143278 3442
rect 143330 3390 143342 3442
rect 143490 3390 143502 3442
rect 143554 3390 143566 3442
rect 138126 3378 138178 3390
rect 142158 3378 142210 3390
rect 146078 3378 146130 3390
rect 147198 3442 147250 3454
rect 147198 3378 147250 3390
rect 148094 3442 148146 3454
rect 148094 3378 148146 3390
rect 24222 3330 24274 3342
rect 24222 3266 24274 3278
rect 25902 3330 25954 3342
rect 25902 3266 25954 3278
rect 27582 3330 27634 3342
rect 27582 3266 27634 3278
rect 29598 3330 29650 3342
rect 29598 3266 29650 3278
rect 30942 3330 30994 3342
rect 30942 3266 30994 3278
rect 32398 3330 32450 3342
rect 32398 3266 32450 3278
rect 34302 3330 34354 3342
rect 34302 3266 34354 3278
rect 35982 3330 36034 3342
rect 35982 3266 36034 3278
rect 37662 3330 37714 3342
rect 37662 3266 37714 3278
rect 39342 3330 39394 3342
rect 39342 3266 39394 3278
rect 41358 3330 41410 3342
rect 41358 3266 41410 3278
rect 42702 3330 42754 3342
rect 42702 3266 42754 3278
rect 44158 3330 44210 3342
rect 44158 3266 44210 3278
rect 46062 3330 46114 3342
rect 46062 3266 46114 3278
rect 47742 3330 47794 3342
rect 47742 3266 47794 3278
rect 49422 3330 49474 3342
rect 49422 3266 49474 3278
rect 51102 3330 51154 3342
rect 51102 3266 51154 3278
rect 53118 3330 53170 3342
rect 53118 3266 53170 3278
rect 54462 3330 54514 3342
rect 54462 3266 54514 3278
rect 55918 3330 55970 3342
rect 55918 3266 55970 3278
rect 57822 3330 57874 3342
rect 57822 3266 57874 3278
rect 59502 3330 59554 3342
rect 59502 3266 59554 3278
rect 61182 3330 61234 3342
rect 61182 3266 61234 3278
rect 62862 3330 62914 3342
rect 62862 3266 62914 3278
rect 64878 3330 64930 3342
rect 64878 3266 64930 3278
rect 66222 3330 66274 3342
rect 66222 3266 66274 3278
rect 67678 3330 67730 3342
rect 67678 3266 67730 3278
rect 69582 3330 69634 3342
rect 69582 3266 69634 3278
rect 71262 3330 71314 3342
rect 71262 3266 71314 3278
rect 72830 3330 72882 3342
rect 72830 3266 72882 3278
rect 73390 3330 73442 3342
rect 73390 3266 73442 3278
rect 74622 3330 74674 3342
rect 74622 3266 74674 3278
rect 75182 3330 75234 3342
rect 75182 3266 75234 3278
rect 94110 3330 94162 3342
rect 94110 3266 94162 3278
rect 95006 3330 95058 3342
rect 95006 3266 95058 3278
rect 96462 3330 96514 3342
rect 96462 3266 96514 3278
rect 102062 3330 102114 3342
rect 102062 3266 102114 3278
rect 102958 3330 103010 3342
rect 102958 3266 103010 3278
rect 105646 3330 105698 3342
rect 105646 3266 105698 3278
rect 108222 3330 108274 3342
rect 108222 3266 108274 3278
rect 113486 3330 113538 3342
rect 113486 3266 113538 3278
rect 114382 3330 114434 3342
rect 114382 3266 114434 3278
rect 117406 3330 117458 3342
rect 117406 3266 117458 3278
rect 121662 3330 121714 3342
rect 121662 3266 121714 3278
rect 122558 3330 122610 3342
rect 122558 3266 122610 3278
rect 133086 3330 133138 3342
rect 133086 3266 133138 3278
rect 133982 3330 134034 3342
rect 133982 3266 134034 3278
rect 137678 3330 137730 3342
rect 137678 3266 137730 3278
rect 140926 3330 140978 3342
rect 140926 3266 140978 3278
rect 141822 3330 141874 3342
rect 141822 3266 141874 3278
rect 144846 3330 144898 3342
rect 144846 3266 144898 3278
rect 146862 3330 146914 3342
rect 146862 3266 146914 3278
rect 147758 3330 147810 3342
rect 147758 3266 147810 3278
rect 1344 3162 148784 3196
rect 1344 3110 38034 3162
rect 38086 3110 38138 3162
rect 38190 3110 38242 3162
rect 38294 3110 74854 3162
rect 74906 3110 74958 3162
rect 75010 3110 75062 3162
rect 75114 3110 111674 3162
rect 111726 3110 111778 3162
rect 111830 3110 111882 3162
rect 111934 3110 148494 3162
rect 148546 3110 148598 3162
rect 148650 3110 148702 3162
rect 148754 3110 148784 3162
rect 1344 3076 148784 3110
rect 104514 2942 104526 2994
rect 104578 2991 104590 2994
rect 105634 2991 105646 2994
rect 104578 2945 105646 2991
rect 104578 2942 104590 2945
rect 105634 2942 105646 2945
rect 105698 2942 105710 2994
rect 139906 2942 139918 2994
rect 139970 2991 139982 2994
rect 140914 2991 140926 2994
rect 139970 2945 140926 2991
rect 139970 2942 139982 2945
rect 140914 2942 140926 2945
rect 140978 2942 140990 2994
<< via1 >>
rect 19624 36822 19676 36874
rect 19728 36822 19780 36874
rect 19832 36822 19884 36874
rect 56444 36822 56496 36874
rect 56548 36822 56600 36874
rect 56652 36822 56704 36874
rect 93264 36822 93316 36874
rect 93368 36822 93420 36874
rect 93472 36822 93524 36874
rect 130084 36822 130136 36874
rect 130188 36822 130240 36874
rect 130292 36822 130344 36874
rect 145854 36542 145906 36594
rect 144846 36430 144898 36482
rect 146862 36430 146914 36482
rect 147758 36318 147810 36370
rect 143838 36206 143890 36258
rect 144286 36206 144338 36258
rect 38034 36038 38086 36090
rect 38138 36038 38190 36090
rect 38242 36038 38294 36090
rect 74854 36038 74906 36090
rect 74958 36038 75010 36090
rect 75062 36038 75114 36090
rect 111674 36038 111726 36090
rect 111778 36038 111830 36090
rect 111882 36038 111934 36090
rect 148494 36038 148546 36090
rect 148598 36038 148650 36090
rect 148702 36038 148754 36090
rect 145966 35758 146018 35810
rect 145070 35646 145122 35698
rect 146974 35646 147026 35698
rect 144286 35534 144338 35586
rect 147758 35534 147810 35586
rect 19624 35254 19676 35306
rect 19728 35254 19780 35306
rect 19832 35254 19884 35306
rect 56444 35254 56496 35306
rect 56548 35254 56600 35306
rect 56652 35254 56704 35306
rect 93264 35254 93316 35306
rect 93368 35254 93420 35306
rect 93472 35254 93524 35306
rect 130084 35254 130136 35306
rect 130188 35254 130240 35306
rect 130292 35254 130344 35306
rect 146078 34974 146130 35026
rect 145070 34862 145122 34914
rect 146862 34862 146914 34914
rect 147758 34750 147810 34802
rect 144510 34638 144562 34690
rect 38034 34470 38086 34522
rect 38138 34470 38190 34522
rect 38242 34470 38294 34522
rect 74854 34470 74906 34522
rect 74958 34470 75010 34522
rect 75062 34470 75114 34522
rect 111674 34470 111726 34522
rect 111778 34470 111830 34522
rect 111882 34470 111934 34522
rect 148494 34470 148546 34522
rect 148598 34470 148650 34522
rect 148702 34470 148754 34522
rect 146414 34078 146466 34130
rect 147086 34078 147138 34130
rect 145406 33966 145458 34018
rect 145854 33966 145906 34018
rect 147758 33966 147810 34018
rect 19624 33686 19676 33738
rect 19728 33686 19780 33738
rect 19832 33686 19884 33738
rect 56444 33686 56496 33738
rect 56548 33686 56600 33738
rect 56652 33686 56704 33738
rect 93264 33686 93316 33738
rect 93368 33686 93420 33738
rect 93472 33686 93524 33738
rect 130084 33686 130136 33738
rect 130188 33686 130240 33738
rect 130292 33686 130344 33738
rect 146302 33294 146354 33346
rect 146862 33294 146914 33346
rect 147758 33182 147810 33234
rect 38034 32902 38086 32954
rect 38138 32902 38190 32954
rect 38242 32902 38294 32954
rect 74854 32902 74906 32954
rect 74958 32902 75010 32954
rect 75062 32902 75114 32954
rect 111674 32902 111726 32954
rect 111778 32902 111830 32954
rect 111882 32902 111934 32954
rect 148494 32902 148546 32954
rect 148598 32902 148650 32954
rect 148702 32902 148754 32954
rect 19624 32118 19676 32170
rect 19728 32118 19780 32170
rect 19832 32118 19884 32170
rect 56444 32118 56496 32170
rect 56548 32118 56600 32170
rect 56652 32118 56704 32170
rect 93264 32118 93316 32170
rect 93368 32118 93420 32170
rect 93472 32118 93524 32170
rect 130084 32118 130136 32170
rect 130188 32118 130240 32170
rect 130292 32118 130344 32170
rect 146862 31726 146914 31778
rect 147758 31614 147810 31666
rect 146302 31502 146354 31554
rect 38034 31334 38086 31386
rect 38138 31334 38190 31386
rect 38242 31334 38294 31386
rect 74854 31334 74906 31386
rect 74958 31334 75010 31386
rect 75062 31334 75114 31386
rect 111674 31334 111726 31386
rect 111778 31334 111830 31386
rect 111882 31334 111934 31386
rect 148494 31334 148546 31386
rect 148598 31334 148650 31386
rect 148702 31334 148754 31386
rect 146414 30942 146466 30994
rect 146862 30942 146914 30994
rect 147758 30830 147810 30882
rect 19624 30550 19676 30602
rect 19728 30550 19780 30602
rect 19832 30550 19884 30602
rect 56444 30550 56496 30602
rect 56548 30550 56600 30602
rect 56652 30550 56704 30602
rect 93264 30550 93316 30602
rect 93368 30550 93420 30602
rect 93472 30550 93524 30602
rect 130084 30550 130136 30602
rect 130188 30550 130240 30602
rect 130292 30550 130344 30602
rect 146302 30158 146354 30210
rect 147086 30158 147138 30210
rect 147758 30046 147810 30098
rect 38034 29766 38086 29818
rect 38138 29766 38190 29818
rect 38242 29766 38294 29818
rect 74854 29766 74906 29818
rect 74958 29766 75010 29818
rect 75062 29766 75114 29818
rect 111674 29766 111726 29818
rect 111778 29766 111830 29818
rect 111882 29766 111934 29818
rect 148494 29766 148546 29818
rect 148598 29766 148650 29818
rect 148702 29766 148754 29818
rect 146414 29374 146466 29426
rect 146862 29374 146914 29426
rect 147758 29262 147810 29314
rect 19624 28982 19676 29034
rect 19728 28982 19780 29034
rect 19832 28982 19884 29034
rect 56444 28982 56496 29034
rect 56548 28982 56600 29034
rect 56652 28982 56704 29034
rect 93264 28982 93316 29034
rect 93368 28982 93420 29034
rect 93472 28982 93524 29034
rect 130084 28982 130136 29034
rect 130188 28982 130240 29034
rect 130292 28982 130344 29034
rect 146302 28590 146354 28642
rect 146862 28590 146914 28642
rect 147758 28590 147810 28642
rect 38034 28198 38086 28250
rect 38138 28198 38190 28250
rect 38242 28198 38294 28250
rect 74854 28198 74906 28250
rect 74958 28198 75010 28250
rect 75062 28198 75114 28250
rect 111674 28198 111726 28250
rect 111778 28198 111830 28250
rect 111882 28198 111934 28250
rect 148494 28198 148546 28250
rect 148598 28198 148650 28250
rect 148702 28198 148754 28250
rect 146414 27806 146466 27858
rect 147086 27806 147138 27858
rect 147758 27694 147810 27746
rect 19624 27414 19676 27466
rect 19728 27414 19780 27466
rect 19832 27414 19884 27466
rect 56444 27414 56496 27466
rect 56548 27414 56600 27466
rect 56652 27414 56704 27466
rect 93264 27414 93316 27466
rect 93368 27414 93420 27466
rect 93472 27414 93524 27466
rect 130084 27414 130136 27466
rect 130188 27414 130240 27466
rect 130292 27414 130344 27466
rect 146302 27134 146354 27186
rect 146862 27022 146914 27074
rect 147758 26910 147810 26962
rect 38034 26630 38086 26682
rect 38138 26630 38190 26682
rect 38242 26630 38294 26682
rect 74854 26630 74906 26682
rect 74958 26630 75010 26682
rect 75062 26630 75114 26682
rect 111674 26630 111726 26682
rect 111778 26630 111830 26682
rect 111882 26630 111934 26682
rect 148494 26630 148546 26682
rect 148598 26630 148650 26682
rect 148702 26630 148754 26682
rect 19624 25846 19676 25898
rect 19728 25846 19780 25898
rect 19832 25846 19884 25898
rect 56444 25846 56496 25898
rect 56548 25846 56600 25898
rect 56652 25846 56704 25898
rect 93264 25846 93316 25898
rect 93368 25846 93420 25898
rect 93472 25846 93524 25898
rect 130084 25846 130136 25898
rect 130188 25846 130240 25898
rect 130292 25846 130344 25898
rect 146862 25454 146914 25506
rect 147758 25342 147810 25394
rect 146302 25230 146354 25282
rect 38034 25062 38086 25114
rect 38138 25062 38190 25114
rect 38242 25062 38294 25114
rect 74854 25062 74906 25114
rect 74958 25062 75010 25114
rect 75062 25062 75114 25114
rect 111674 25062 111726 25114
rect 111778 25062 111830 25114
rect 111882 25062 111934 25114
rect 148494 25062 148546 25114
rect 148598 25062 148650 25114
rect 148702 25062 148754 25114
rect 146862 24670 146914 24722
rect 146414 24558 146466 24610
rect 147758 24558 147810 24610
rect 19624 24278 19676 24330
rect 19728 24278 19780 24330
rect 19832 24278 19884 24330
rect 56444 24278 56496 24330
rect 56548 24278 56600 24330
rect 56652 24278 56704 24330
rect 93264 24278 93316 24330
rect 93368 24278 93420 24330
rect 93472 24278 93524 24330
rect 130084 24278 130136 24330
rect 130188 24278 130240 24330
rect 130292 24278 130344 24330
rect 146862 23886 146914 23938
rect 147758 23774 147810 23826
rect 146302 23662 146354 23714
rect 38034 23494 38086 23546
rect 38138 23494 38190 23546
rect 38242 23494 38294 23546
rect 74854 23494 74906 23546
rect 74958 23494 75010 23546
rect 75062 23494 75114 23546
rect 111674 23494 111726 23546
rect 111778 23494 111830 23546
rect 111882 23494 111934 23546
rect 148494 23494 148546 23546
rect 148598 23494 148650 23546
rect 148702 23494 148754 23546
rect 146414 23102 146466 23154
rect 146862 23102 146914 23154
rect 147758 22990 147810 23042
rect 19624 22710 19676 22762
rect 19728 22710 19780 22762
rect 19832 22710 19884 22762
rect 56444 22710 56496 22762
rect 56548 22710 56600 22762
rect 56652 22710 56704 22762
rect 93264 22710 93316 22762
rect 93368 22710 93420 22762
rect 93472 22710 93524 22762
rect 130084 22710 130136 22762
rect 130188 22710 130240 22762
rect 130292 22710 130344 22762
rect 146302 22318 146354 22370
rect 146862 22318 146914 22370
rect 147758 22206 147810 22258
rect 38034 21926 38086 21978
rect 38138 21926 38190 21978
rect 38242 21926 38294 21978
rect 74854 21926 74906 21978
rect 74958 21926 75010 21978
rect 75062 21926 75114 21978
rect 111674 21926 111726 21978
rect 111778 21926 111830 21978
rect 111882 21926 111934 21978
rect 148494 21926 148546 21978
rect 148598 21926 148650 21978
rect 148702 21926 148754 21978
rect 146862 21534 146914 21586
rect 146414 21422 146466 21474
rect 147758 21422 147810 21474
rect 19624 21142 19676 21194
rect 19728 21142 19780 21194
rect 19832 21142 19884 21194
rect 56444 21142 56496 21194
rect 56548 21142 56600 21194
rect 56652 21142 56704 21194
rect 93264 21142 93316 21194
rect 93368 21142 93420 21194
rect 93472 21142 93524 21194
rect 130084 21142 130136 21194
rect 130188 21142 130240 21194
rect 130292 21142 130344 21194
rect 146302 20750 146354 20802
rect 146862 20750 146914 20802
rect 147758 20638 147810 20690
rect 38034 20358 38086 20410
rect 38138 20358 38190 20410
rect 38242 20358 38294 20410
rect 74854 20358 74906 20410
rect 74958 20358 75010 20410
rect 75062 20358 75114 20410
rect 111674 20358 111726 20410
rect 111778 20358 111830 20410
rect 111882 20358 111934 20410
rect 148494 20358 148546 20410
rect 148598 20358 148650 20410
rect 148702 20358 148754 20410
rect 19624 19574 19676 19626
rect 19728 19574 19780 19626
rect 19832 19574 19884 19626
rect 56444 19574 56496 19626
rect 56548 19574 56600 19626
rect 56652 19574 56704 19626
rect 93264 19574 93316 19626
rect 93368 19574 93420 19626
rect 93472 19574 93524 19626
rect 130084 19574 130136 19626
rect 130188 19574 130240 19626
rect 130292 19574 130344 19626
rect 146302 19182 146354 19234
rect 146862 19182 146914 19234
rect 147758 19070 147810 19122
rect 38034 18790 38086 18842
rect 38138 18790 38190 18842
rect 38242 18790 38294 18842
rect 74854 18790 74906 18842
rect 74958 18790 75010 18842
rect 75062 18790 75114 18842
rect 111674 18790 111726 18842
rect 111778 18790 111830 18842
rect 111882 18790 111934 18842
rect 148494 18790 148546 18842
rect 148598 18790 148650 18842
rect 148702 18790 148754 18842
rect 114046 18622 114098 18674
rect 113710 18398 113762 18450
rect 146862 18398 146914 18450
rect 113150 18286 113202 18338
rect 146414 18286 146466 18338
rect 147758 18286 147810 18338
rect 19624 18006 19676 18058
rect 19728 18006 19780 18058
rect 19832 18006 19884 18058
rect 56444 18006 56496 18058
rect 56548 18006 56600 18058
rect 56652 18006 56704 18058
rect 93264 18006 93316 18058
rect 93368 18006 93420 18058
rect 93472 18006 93524 18058
rect 130084 18006 130136 18058
rect 130188 18006 130240 18058
rect 130292 18006 130344 18058
rect 146862 17614 146914 17666
rect 147758 17502 147810 17554
rect 146302 17390 146354 17442
rect 38034 17222 38086 17274
rect 38138 17222 38190 17274
rect 38242 17222 38294 17274
rect 74854 17222 74906 17274
rect 74958 17222 75010 17274
rect 75062 17222 75114 17274
rect 111674 17222 111726 17274
rect 111778 17222 111830 17274
rect 111882 17222 111934 17274
rect 148494 17222 148546 17274
rect 148598 17222 148650 17274
rect 148702 17222 148754 17274
rect 146414 16942 146466 16994
rect 146862 16830 146914 16882
rect 147758 16830 147810 16882
rect 19624 16438 19676 16490
rect 19728 16438 19780 16490
rect 19832 16438 19884 16490
rect 56444 16438 56496 16490
rect 56548 16438 56600 16490
rect 56652 16438 56704 16490
rect 93264 16438 93316 16490
rect 93368 16438 93420 16490
rect 93472 16438 93524 16490
rect 130084 16438 130136 16490
rect 130188 16438 130240 16490
rect 130292 16438 130344 16490
rect 146862 16046 146914 16098
rect 147758 15934 147810 15986
rect 146302 15822 146354 15874
rect 38034 15654 38086 15706
rect 38138 15654 38190 15706
rect 38242 15654 38294 15706
rect 74854 15654 74906 15706
rect 74958 15654 75010 15706
rect 75062 15654 75114 15706
rect 111674 15654 111726 15706
rect 111778 15654 111830 15706
rect 111882 15654 111934 15706
rect 148494 15654 148546 15706
rect 148598 15654 148650 15706
rect 148702 15654 148754 15706
rect 146414 15374 146466 15426
rect 146862 15262 146914 15314
rect 147758 15150 147810 15202
rect 19624 14870 19676 14922
rect 19728 14870 19780 14922
rect 19832 14870 19884 14922
rect 56444 14870 56496 14922
rect 56548 14870 56600 14922
rect 56652 14870 56704 14922
rect 93264 14870 93316 14922
rect 93368 14870 93420 14922
rect 93472 14870 93524 14922
rect 130084 14870 130136 14922
rect 130188 14870 130240 14922
rect 130292 14870 130344 14922
rect 146302 14478 146354 14530
rect 146862 14478 146914 14530
rect 147758 14366 147810 14418
rect 38034 14086 38086 14138
rect 38138 14086 38190 14138
rect 38242 14086 38294 14138
rect 74854 14086 74906 14138
rect 74958 14086 75010 14138
rect 75062 14086 75114 14138
rect 111674 14086 111726 14138
rect 111778 14086 111830 14138
rect 111882 14086 111934 14138
rect 148494 14086 148546 14138
rect 148598 14086 148650 14138
rect 148702 14086 148754 14138
rect 19624 13302 19676 13354
rect 19728 13302 19780 13354
rect 19832 13302 19884 13354
rect 56444 13302 56496 13354
rect 56548 13302 56600 13354
rect 56652 13302 56704 13354
rect 93264 13302 93316 13354
rect 93368 13302 93420 13354
rect 93472 13302 93524 13354
rect 130084 13302 130136 13354
rect 130188 13302 130240 13354
rect 130292 13302 130344 13354
rect 146302 12910 146354 12962
rect 146862 12910 146914 12962
rect 101502 12798 101554 12850
rect 101838 12798 101890 12850
rect 147758 12798 147810 12850
rect 38034 12518 38086 12570
rect 38138 12518 38190 12570
rect 38242 12518 38294 12570
rect 74854 12518 74906 12570
rect 74958 12518 75010 12570
rect 75062 12518 75114 12570
rect 111674 12518 111726 12570
rect 111778 12518 111830 12570
rect 111882 12518 111934 12570
rect 148494 12518 148546 12570
rect 148598 12518 148650 12570
rect 148702 12518 148754 12570
rect 100718 12350 100770 12402
rect 100494 12126 100546 12178
rect 146862 12126 146914 12178
rect 101166 12014 101218 12066
rect 146414 12014 146466 12066
rect 147758 12014 147810 12066
rect 19624 11734 19676 11786
rect 19728 11734 19780 11786
rect 19832 11734 19884 11786
rect 56444 11734 56496 11786
rect 56548 11734 56600 11786
rect 56652 11734 56704 11786
rect 93264 11734 93316 11786
rect 93368 11734 93420 11786
rect 93472 11734 93524 11786
rect 130084 11734 130136 11786
rect 130188 11734 130240 11786
rect 130292 11734 130344 11786
rect 146302 11342 146354 11394
rect 146862 11342 146914 11394
rect 99486 11230 99538 11282
rect 99822 11230 99874 11282
rect 147758 11230 147810 11282
rect 38034 10950 38086 11002
rect 38138 10950 38190 11002
rect 38242 10950 38294 11002
rect 74854 10950 74906 11002
rect 74958 10950 75010 11002
rect 75062 10950 75114 11002
rect 111674 10950 111726 11002
rect 111778 10950 111830 11002
rect 111882 10950 111934 11002
rect 148494 10950 148546 11002
rect 148598 10950 148650 11002
rect 148702 10950 148754 11002
rect 147758 10670 147810 10722
rect 148094 10558 148146 10610
rect 147310 10446 147362 10498
rect 19624 10166 19676 10218
rect 19728 10166 19780 10218
rect 19832 10166 19884 10218
rect 56444 10166 56496 10218
rect 56548 10166 56600 10218
rect 56652 10166 56704 10218
rect 93264 10166 93316 10218
rect 93368 10166 93420 10218
rect 93472 10166 93524 10218
rect 130084 10166 130136 10218
rect 130188 10166 130240 10218
rect 130292 10166 130344 10218
rect 148094 9662 148146 9714
rect 147310 9550 147362 9602
rect 147758 9550 147810 9602
rect 38034 9382 38086 9434
rect 38138 9382 38190 9434
rect 38242 9382 38294 9434
rect 74854 9382 74906 9434
rect 74958 9382 75010 9434
rect 75062 9382 75114 9434
rect 111674 9382 111726 9434
rect 111778 9382 111830 9434
rect 111882 9382 111934 9434
rect 148494 9382 148546 9434
rect 148598 9382 148650 9434
rect 148702 9382 148754 9434
rect 147758 9102 147810 9154
rect 147310 8990 147362 9042
rect 148094 8990 148146 9042
rect 19624 8598 19676 8650
rect 19728 8598 19780 8650
rect 19832 8598 19884 8650
rect 56444 8598 56496 8650
rect 56548 8598 56600 8650
rect 56652 8598 56704 8650
rect 93264 8598 93316 8650
rect 93368 8598 93420 8650
rect 93472 8598 93524 8650
rect 130084 8598 130136 8650
rect 130188 8598 130240 8650
rect 130292 8598 130344 8650
rect 134878 8094 134930 8146
rect 135326 8094 135378 8146
rect 148094 8094 148146 8146
rect 134542 7982 134594 8034
rect 147310 7982 147362 8034
rect 147758 7982 147810 8034
rect 38034 7814 38086 7866
rect 38138 7814 38190 7866
rect 38242 7814 38294 7866
rect 74854 7814 74906 7866
rect 74958 7814 75010 7866
rect 75062 7814 75114 7866
rect 111674 7814 111726 7866
rect 111778 7814 111830 7866
rect 111882 7814 111934 7866
rect 148494 7814 148546 7866
rect 148598 7814 148650 7866
rect 148702 7814 148754 7866
rect 99598 7646 99650 7698
rect 113486 7646 113538 7698
rect 99374 7422 99426 7474
rect 113150 7422 113202 7474
rect 19624 7030 19676 7082
rect 19728 7030 19780 7082
rect 19832 7030 19884 7082
rect 56444 7030 56496 7082
rect 56548 7030 56600 7082
rect 56652 7030 56704 7082
rect 93264 7030 93316 7082
rect 93368 7030 93420 7082
rect 93472 7030 93524 7082
rect 130084 7030 130136 7082
rect 130188 7030 130240 7082
rect 130292 7030 130344 7082
rect 129278 6526 129330 6578
rect 147310 6526 147362 6578
rect 148094 6526 148146 6578
rect 103518 6414 103570 6466
rect 111582 6414 111634 6466
rect 128606 6414 128658 6466
rect 130958 6414 131010 6466
rect 140926 6414 140978 6466
rect 141262 6414 141314 6466
rect 147758 6414 147810 6466
rect 38034 6246 38086 6298
rect 38138 6246 38190 6298
rect 38242 6246 38294 6298
rect 74854 6246 74906 6298
rect 74958 6246 75010 6298
rect 75062 6246 75114 6298
rect 111674 6246 111726 6298
rect 111778 6246 111830 6298
rect 111882 6246 111934 6298
rect 148494 6246 148546 6298
rect 148598 6246 148650 6298
rect 148702 6246 148754 6298
rect 84478 6078 84530 6130
rect 88398 6078 88450 6130
rect 105534 6078 105586 6130
rect 112142 6078 112194 6130
rect 131406 6078 131458 6130
rect 140814 6078 140866 6130
rect 141710 6078 141762 6130
rect 142606 6078 142658 6130
rect 130062 5966 130114 6018
rect 147758 5966 147810 6018
rect 103966 5854 104018 5906
rect 104414 5854 104466 5906
rect 105198 5854 105250 5906
rect 111246 5854 111298 5906
rect 111918 5854 111970 5906
rect 129726 5854 129778 5906
rect 131070 5854 131122 5906
rect 140478 5854 140530 5906
rect 141374 5854 141426 5906
rect 142270 5854 142322 5906
rect 148094 5854 148146 5906
rect 82686 5742 82738 5794
rect 83582 5742 83634 5794
rect 99598 5742 99650 5794
rect 102510 5742 102562 5794
rect 102958 5742 103010 5794
rect 103518 5742 103570 5794
rect 110238 5742 110290 5794
rect 110798 5742 110850 5794
rect 113262 5742 113314 5794
rect 114158 5742 114210 5794
rect 115614 5742 115666 5794
rect 116062 5742 116114 5794
rect 117070 5742 117122 5794
rect 117518 5742 117570 5794
rect 117854 5742 117906 5794
rect 118302 5742 118354 5794
rect 119198 5742 119250 5794
rect 123902 5742 123954 5794
rect 127598 5742 127650 5794
rect 128270 5742 128322 5794
rect 129278 5742 129330 5794
rect 130510 5742 130562 5794
rect 131966 5742 132018 5794
rect 132862 5742 132914 5794
rect 133758 5742 133810 5794
rect 138798 5742 138850 5794
rect 139582 5742 139634 5794
rect 139918 5742 139970 5794
rect 143054 5742 143106 5794
rect 143502 5742 143554 5794
rect 147310 5742 147362 5794
rect 19624 5462 19676 5514
rect 19728 5462 19780 5514
rect 19832 5462 19884 5514
rect 56444 5462 56496 5514
rect 56548 5462 56600 5514
rect 56652 5462 56704 5514
rect 93264 5462 93316 5514
rect 93368 5462 93420 5514
rect 93472 5462 93524 5514
rect 130084 5462 130136 5514
rect 130188 5462 130240 5514
rect 130292 5462 130344 5514
rect 104862 5294 104914 5346
rect 142158 5294 142210 5346
rect 77646 5182 77698 5234
rect 88062 5182 88114 5234
rect 90190 5182 90242 5234
rect 103070 5182 103122 5234
rect 109566 5182 109618 5234
rect 115390 5182 115442 5234
rect 134654 5182 134706 5234
rect 75854 5070 75906 5122
rect 78542 5070 78594 5122
rect 79438 5070 79490 5122
rect 82126 5070 82178 5122
rect 83246 5070 83298 5122
rect 84254 5070 84306 5122
rect 87614 5070 87666 5122
rect 98366 5070 98418 5122
rect 99038 5070 99090 5122
rect 102622 5070 102674 5122
rect 104526 5070 104578 5122
rect 111806 5070 111858 5122
rect 117630 5070 117682 5122
rect 122782 5070 122834 5122
rect 127374 5070 127426 5122
rect 136110 5070 136162 5122
rect 140254 5070 140306 5122
rect 141822 5070 141874 5122
rect 146414 5070 146466 5122
rect 147310 5070 147362 5122
rect 80558 4958 80610 5010
rect 80894 4958 80946 5010
rect 82910 4958 82962 5010
rect 83918 4958 83970 5010
rect 85598 4958 85650 5010
rect 85934 4958 85986 5010
rect 87278 4958 87330 5010
rect 88958 4958 89010 5010
rect 89294 4958 89346 5010
rect 99486 4958 99538 5010
rect 100382 4958 100434 5010
rect 102062 4958 102114 5010
rect 103742 4958 103794 5010
rect 104190 4958 104242 5010
rect 105534 4958 105586 5010
rect 105870 4958 105922 5010
rect 106430 4958 106482 5010
rect 106766 4958 106818 5010
rect 110014 4958 110066 5010
rect 110350 4958 110402 5010
rect 111022 4958 111074 5010
rect 111470 4958 111522 5010
rect 112142 4958 112194 5010
rect 112814 4958 112866 5010
rect 113150 4958 113202 5010
rect 114606 4958 114658 5010
rect 115950 4958 116002 5010
rect 116286 4958 116338 5010
rect 117070 4958 117122 5010
rect 118190 4958 118242 5010
rect 118526 4958 118578 5010
rect 119086 4958 119138 5010
rect 119422 4958 119474 5010
rect 119982 4958 120034 5010
rect 120318 4958 120370 5010
rect 123566 4958 123618 5010
rect 123902 4958 123954 5010
rect 125022 4958 125074 5010
rect 125358 4958 125410 5010
rect 125918 4958 125970 5010
rect 126254 4958 126306 5010
rect 127038 4958 127090 5010
rect 127934 4958 127986 5010
rect 128270 4958 128322 5010
rect 129054 4958 129106 5010
rect 130174 4958 130226 5010
rect 131070 4958 131122 5010
rect 132974 4958 133026 5010
rect 133310 4958 133362 5010
rect 133870 4958 133922 5010
rect 134206 4958 134258 5010
rect 135550 4958 135602 5010
rect 137454 4958 137506 5010
rect 137790 4958 137842 5010
rect 139134 4958 139186 5010
rect 139470 4958 139522 5010
rect 141150 4958 141202 5010
rect 141598 4958 141650 5010
rect 142830 4958 142882 5010
rect 143166 4958 143218 5010
rect 143726 4958 143778 5010
rect 144062 4958 144114 5010
rect 148094 4958 148146 5010
rect 81342 4846 81394 4898
rect 82350 4846 82402 4898
rect 86382 4846 86434 4898
rect 89742 4846 89794 4898
rect 98030 4846 98082 4898
rect 99822 4846 99874 4898
rect 101166 4846 101218 4898
rect 101614 4846 101666 4898
rect 113598 4846 113650 4898
rect 114158 4846 114210 4898
rect 114942 4846 114994 4898
rect 121102 4846 121154 4898
rect 129614 4846 129666 4898
rect 130510 4846 130562 4898
rect 131630 4846 131682 4898
rect 132078 4846 132130 4898
rect 135102 4846 135154 4898
rect 136782 4846 136834 4898
rect 138686 4846 138738 4898
rect 146862 4846 146914 4898
rect 147758 4846 147810 4898
rect 38034 4678 38086 4730
rect 38138 4678 38190 4730
rect 38242 4678 38294 4730
rect 74854 4678 74906 4730
rect 74958 4678 75010 4730
rect 75062 4678 75114 4730
rect 111674 4678 111726 4730
rect 111778 4678 111830 4730
rect 111882 4678 111934 4730
rect 148494 4678 148546 4730
rect 148598 4678 148650 4730
rect 148702 4678 148754 4730
rect 9774 4510 9826 4562
rect 11342 4510 11394 4562
rect 13022 4510 13074 4562
rect 15150 4510 15202 4562
rect 22542 4510 22594 4562
rect 76078 4510 76130 4562
rect 77870 4510 77922 4562
rect 79662 4510 79714 4562
rect 82126 4510 82178 4562
rect 85374 4510 85426 4562
rect 99486 4510 99538 4562
rect 101390 4510 101442 4562
rect 104302 4510 104354 4562
rect 106430 4510 106482 4562
rect 106990 4510 107042 4562
rect 109006 4510 109058 4562
rect 111582 4510 111634 4562
rect 112142 4510 112194 4562
rect 113262 4510 113314 4562
rect 114942 4510 114994 4562
rect 117070 4510 117122 4562
rect 118974 4510 119026 4562
rect 121438 4510 121490 4562
rect 123230 4510 123282 4562
rect 125358 4510 125410 4562
rect 127262 4510 127314 4562
rect 130734 4510 130786 4562
rect 132862 4510 132914 4562
rect 134094 4510 134146 4562
rect 135662 4510 135714 4562
rect 138238 4510 138290 4562
rect 140254 4510 140306 4562
rect 142158 4510 142210 4562
rect 143726 4510 143778 4562
rect 147758 4510 147810 4562
rect 19406 4398 19458 4450
rect 73950 4398 74002 4450
rect 75294 4398 75346 4450
rect 75630 4398 75682 4450
rect 76974 4398 77026 4450
rect 77310 4398 77362 4450
rect 78206 4398 78258 4450
rect 79102 4398 79154 4450
rect 79998 4398 80050 4450
rect 80446 4398 80498 4450
rect 81342 4398 81394 4450
rect 81678 4398 81730 4450
rect 84814 4398 84866 4450
rect 88174 4398 88226 4450
rect 89630 4398 89682 4450
rect 90750 4398 90802 4450
rect 91310 4398 91362 4450
rect 97694 4398 97746 4450
rect 98478 4398 98530 4450
rect 100382 4398 100434 4450
rect 102174 4398 102226 4450
rect 102734 4398 102786 4450
rect 105534 4398 105586 4450
rect 109790 4398 109842 4450
rect 110574 4398 110626 4450
rect 114270 4398 114322 4450
rect 115950 4398 116002 4450
rect 116510 4398 116562 4450
rect 117854 4398 117906 4450
rect 118414 4398 118466 4450
rect 119982 4398 120034 4450
rect 122110 4398 122162 4450
rect 122670 4398 122722 4450
rect 124350 4398 124402 4450
rect 124798 4398 124850 4450
rect 126366 4398 126418 4450
rect 126702 4398 126754 4450
rect 128270 4398 128322 4450
rect 129838 4398 129890 4450
rect 131854 4398 131906 4450
rect 133534 4398 133586 4450
rect 135102 4398 135154 4450
rect 137230 4398 137282 4450
rect 139134 4398 139186 4450
rect 139582 4398 139634 4450
rect 141150 4398 141202 4450
rect 141598 4398 141650 4450
rect 143166 4398 143218 4450
rect 146862 4398 146914 4450
rect 8318 4286 8370 4338
rect 8878 4286 8930 4338
rect 18958 4286 19010 4338
rect 22206 4286 22258 4338
rect 78878 4286 78930 4338
rect 82686 4286 82738 4338
rect 84590 4286 84642 4338
rect 86158 4286 86210 4338
rect 87950 4286 88002 4338
rect 89406 4286 89458 4338
rect 90526 4286 90578 4338
rect 97358 4286 97410 4338
rect 98702 4286 98754 4338
rect 100606 4286 100658 4338
rect 101054 4286 101106 4338
rect 103294 4286 103346 4338
rect 103966 4286 104018 4338
rect 105310 4286 105362 4338
rect 109454 4286 109506 4338
rect 110462 4286 110514 4338
rect 114046 4286 114098 4338
rect 119646 4286 119698 4338
rect 120990 4286 121042 4338
rect 127934 4286 127986 4338
rect 129614 4286 129666 4338
rect 130398 4286 130450 4338
rect 131742 4286 131794 4338
rect 134766 4286 134818 4338
rect 137118 4286 137170 4338
rect 142830 4286 142882 4338
rect 144062 4286 144114 4338
rect 145294 4286 145346 4338
rect 147086 4286 147138 4338
rect 148094 4286 148146 4338
rect 6638 4174 6690 4226
rect 7310 4174 7362 4226
rect 17950 4174 18002 4226
rect 21758 4174 21810 4226
rect 22990 4174 23042 4226
rect 25566 4174 25618 4226
rect 32622 4174 32674 4226
rect 37102 4174 37154 4226
rect 44382 4174 44434 4226
rect 48862 4174 48914 4226
rect 56142 4174 56194 4226
rect 60622 4174 60674 4226
rect 67902 4174 67954 4226
rect 73278 4174 73330 4226
rect 74398 4174 74450 4226
rect 83358 4174 83410 4226
rect 86718 4174 86770 4226
rect 93550 4174 93602 4226
rect 94446 4174 94498 4226
rect 95902 4174 95954 4226
rect 107438 4174 107490 4226
rect 107886 4174 107938 4226
rect 108558 4174 108610 4226
rect 128942 4174 128994 4226
rect 136110 4174 136162 4226
rect 144846 4174 144898 4226
rect 145966 4174 146018 4226
rect 146414 4174 146466 4226
rect 99150 4062 99202 4114
rect 102958 4062 103010 4114
rect 106094 4062 106146 4114
rect 111246 4062 111298 4114
rect 113598 4062 113650 4114
rect 116734 4062 116786 4114
rect 118638 4062 118690 4114
rect 122894 4062 122946 4114
rect 125022 4062 125074 4114
rect 126926 4062 126978 4114
rect 132526 4062 132578 4114
rect 137902 4062 137954 4114
rect 139918 4062 139970 4114
rect 141822 4062 141874 4114
rect 19624 3894 19676 3946
rect 19728 3894 19780 3946
rect 19832 3894 19884 3946
rect 56444 3894 56496 3946
rect 56548 3894 56600 3946
rect 56652 3894 56704 3946
rect 93264 3894 93316 3946
rect 93368 3894 93420 3946
rect 93472 3894 93524 3946
rect 130084 3894 130136 3946
rect 130188 3894 130240 3946
rect 130292 3894 130344 3946
rect 98926 3726 98978 3778
rect 100718 3726 100770 3778
rect 101054 3726 101106 3778
rect 104974 3726 105026 3778
rect 110574 3726 110626 3778
rect 112478 3726 112530 3778
rect 112814 3726 112866 3778
rect 115614 3726 115666 3778
rect 115950 3726 116002 3778
rect 120318 3726 120370 3778
rect 120654 3726 120706 3778
rect 124574 3726 124626 3778
rect 129726 3726 129778 3778
rect 130062 3726 130114 3778
rect 132414 3726 132466 3778
rect 136334 3726 136386 3778
rect 136670 3726 136722 3778
rect 140254 3726 140306 3778
rect 143838 3726 143890 3778
rect 144174 3726 144226 3778
rect 8206 3614 8258 3666
rect 10222 3614 10274 3666
rect 13918 3614 13970 3666
rect 17502 3614 17554 3666
rect 78766 3614 78818 3666
rect 82686 3614 82738 3666
rect 86942 3614 86994 3666
rect 90526 3614 90578 3666
rect 97134 3614 97186 3666
rect 126030 3614 126082 3666
rect 126590 3614 126642 3666
rect 6750 3502 6802 3554
rect 8878 3502 8930 3554
rect 11006 3502 11058 3554
rect 12798 3502 12850 3554
rect 14926 3502 14978 3554
rect 16718 3502 16770 3554
rect 20078 3502 20130 3554
rect 20638 3502 20690 3554
rect 22654 3502 22706 3554
rect 73726 3502 73778 3554
rect 75518 3502 75570 3554
rect 76302 3502 76354 3554
rect 78094 3502 78146 3554
rect 80222 3502 80274 3554
rect 82014 3502 82066 3554
rect 85374 3502 85426 3554
rect 86494 3502 86546 3554
rect 88174 3502 88226 3554
rect 89854 3502 89906 3554
rect 91982 3502 92034 3554
rect 93774 3502 93826 3554
rect 98590 3502 98642 3554
rect 104190 3502 104242 3554
rect 104638 3502 104690 3554
rect 106766 3502 106818 3554
rect 110238 3502 110290 3554
rect 111806 3502 111858 3554
rect 114606 3502 114658 3554
rect 116734 3502 116786 3554
rect 119646 3502 119698 3554
rect 124238 3502 124290 3554
rect 127486 3502 127538 3554
rect 131406 3502 131458 3554
rect 132078 3502 132130 3554
rect 134206 3502 134258 3554
rect 139918 3502 139970 3554
rect 141150 3502 141202 3554
rect 145070 3502 145122 3554
rect 145630 3502 145682 3554
rect 6078 3390 6130 3442
rect 11902 3390 11954 3442
rect 15822 3390 15874 3442
rect 19182 3390 19234 3442
rect 21758 3390 21810 3442
rect 23438 3390 23490 3442
rect 23886 3390 23938 3442
rect 25566 3390 25618 3442
rect 26798 3390 26850 3442
rect 27246 3390 27298 3442
rect 28590 3390 28642 3442
rect 29262 3390 29314 3442
rect 30158 3390 30210 3442
rect 30606 3390 30658 3442
rect 32062 3390 32114 3442
rect 33518 3390 33570 3442
rect 33966 3390 34018 3442
rect 35198 3390 35250 3442
rect 35646 3390 35698 3442
rect 37326 3390 37378 3442
rect 38558 3390 38610 3442
rect 39006 3390 39058 3442
rect 40350 3390 40402 3442
rect 41022 3390 41074 3442
rect 41918 3390 41970 3442
rect 42366 3390 42418 3442
rect 43822 3390 43874 3442
rect 45278 3390 45330 3442
rect 45726 3390 45778 3442
rect 46958 3390 47010 3442
rect 47406 3390 47458 3442
rect 49086 3390 49138 3442
rect 50318 3390 50370 3442
rect 50766 3390 50818 3442
rect 52110 3390 52162 3442
rect 52782 3390 52834 3442
rect 53678 3390 53730 3442
rect 54126 3390 54178 3442
rect 55582 3390 55634 3442
rect 57038 3390 57090 3442
rect 57486 3390 57538 3442
rect 58718 3390 58770 3442
rect 59166 3390 59218 3442
rect 60846 3390 60898 3442
rect 62078 3390 62130 3442
rect 62526 3390 62578 3442
rect 63870 3390 63922 3442
rect 64542 3390 64594 3442
rect 65438 3390 65490 3442
rect 65886 3390 65938 3442
rect 67342 3390 67394 3442
rect 68798 3390 68850 3442
rect 69246 3390 69298 3442
rect 70478 3390 70530 3442
rect 70926 3390 70978 3442
rect 72494 3390 72546 3442
rect 74286 3390 74338 3442
rect 77198 3390 77250 3442
rect 81118 3390 81170 3442
rect 84702 3390 84754 3442
rect 86158 3390 86210 3442
rect 88958 3390 89010 3442
rect 92878 3390 92930 3442
rect 94670 3390 94722 3442
rect 96126 3390 96178 3442
rect 97806 3390 97858 3442
rect 98366 3390 98418 3442
rect 99934 3390 99986 3442
rect 100494 3390 100546 3442
rect 101726 3390 101778 3442
rect 102622 3390 102674 3442
rect 104078 3390 104130 3442
rect 105982 3390 106034 3442
rect 106542 3390 106594 3442
rect 107886 3390 107938 3442
rect 108670 3390 108722 3442
rect 109454 3390 109506 3442
rect 110014 3390 110066 3442
rect 111694 3390 111746 3442
rect 113822 3390 113874 3442
rect 116510 3390 116562 3442
rect 117742 3390 117794 3442
rect 118302 3390 118354 3442
rect 118638 3390 118690 3442
rect 119534 3390 119586 3442
rect 121326 3390 121378 3442
rect 122222 3390 122274 3442
rect 123678 3390 123730 3442
rect 124014 3390 124066 3442
rect 125246 3390 125298 3442
rect 125582 3390 125634 3442
rect 127262 3390 127314 3442
rect 128046 3390 128098 3442
rect 128942 3390 128994 3442
rect 129390 3390 129442 3442
rect 131294 3390 131346 3442
rect 133422 3390 133474 3442
rect 135550 3390 135602 3442
rect 136110 3390 136162 3442
rect 137342 3390 137394 3442
rect 138126 3390 138178 3442
rect 139358 3390 139410 3442
rect 139582 3390 139634 3442
rect 142158 3390 142210 3442
rect 143278 3390 143330 3442
rect 143502 3390 143554 3442
rect 146078 3390 146130 3442
rect 147198 3390 147250 3442
rect 148094 3390 148146 3442
rect 24222 3278 24274 3330
rect 25902 3278 25954 3330
rect 27582 3278 27634 3330
rect 29598 3278 29650 3330
rect 30942 3278 30994 3330
rect 32398 3278 32450 3330
rect 34302 3278 34354 3330
rect 35982 3278 36034 3330
rect 37662 3278 37714 3330
rect 39342 3278 39394 3330
rect 41358 3278 41410 3330
rect 42702 3278 42754 3330
rect 44158 3278 44210 3330
rect 46062 3278 46114 3330
rect 47742 3278 47794 3330
rect 49422 3278 49474 3330
rect 51102 3278 51154 3330
rect 53118 3278 53170 3330
rect 54462 3278 54514 3330
rect 55918 3278 55970 3330
rect 57822 3278 57874 3330
rect 59502 3278 59554 3330
rect 61182 3278 61234 3330
rect 62862 3278 62914 3330
rect 64878 3278 64930 3330
rect 66222 3278 66274 3330
rect 67678 3278 67730 3330
rect 69582 3278 69634 3330
rect 71262 3278 71314 3330
rect 72830 3278 72882 3330
rect 73390 3278 73442 3330
rect 74622 3278 74674 3330
rect 75182 3278 75234 3330
rect 94110 3278 94162 3330
rect 95006 3278 95058 3330
rect 96462 3278 96514 3330
rect 102062 3278 102114 3330
rect 102958 3278 103010 3330
rect 105646 3278 105698 3330
rect 108222 3278 108274 3330
rect 113486 3278 113538 3330
rect 114382 3278 114434 3330
rect 117406 3278 117458 3330
rect 121662 3278 121714 3330
rect 122558 3278 122610 3330
rect 133086 3278 133138 3330
rect 133982 3278 134034 3330
rect 137678 3278 137730 3330
rect 140926 3278 140978 3330
rect 141822 3278 141874 3330
rect 144846 3278 144898 3330
rect 146862 3278 146914 3330
rect 147758 3278 147810 3330
rect 38034 3110 38086 3162
rect 38138 3110 38190 3162
rect 38242 3110 38294 3162
rect 74854 3110 74906 3162
rect 74958 3110 75010 3162
rect 75062 3110 75114 3162
rect 111674 3110 111726 3162
rect 111778 3110 111830 3162
rect 111882 3110 111934 3162
rect 148494 3110 148546 3162
rect 148598 3110 148650 3162
rect 148702 3110 148754 3162
rect 104526 2942 104578 2994
rect 105646 2942 105698 2994
rect 139918 2942 139970 2994
rect 140926 2942 140978 2994
<< metal2 >>
rect 146076 38836 146132 38846
rect 145964 37940 146020 37950
rect 145852 37044 145908 37054
rect 19622 36876 19886 36886
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19622 36810 19886 36820
rect 56442 36876 56706 36886
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56442 36810 56706 36820
rect 93262 36876 93526 36886
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93262 36810 93526 36820
rect 130082 36876 130346 36886
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130082 36810 130346 36820
rect 145852 36594 145908 36988
rect 145852 36542 145854 36594
rect 145906 36542 145908 36594
rect 145852 36530 145908 36542
rect 144284 36484 144340 36494
rect 141708 36260 141764 36270
rect 38032 36092 38296 36102
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38032 36026 38296 36036
rect 74852 36092 75116 36102
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 74852 36026 75116 36036
rect 111672 36092 111936 36102
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111672 36026 111936 36036
rect 19622 35308 19886 35318
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19622 35242 19886 35252
rect 56442 35308 56706 35318
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56442 35242 56706 35252
rect 93262 35308 93526 35318
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93262 35242 93526 35252
rect 130082 35308 130346 35318
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130082 35242 130346 35252
rect 38032 34524 38296 34534
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38032 34458 38296 34468
rect 74852 34524 75116 34534
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 74852 34458 75116 34468
rect 111672 34524 111936 34534
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111672 34458 111936 34468
rect 139356 34020 139412 34030
rect 19622 33740 19886 33750
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19622 33674 19886 33684
rect 56442 33740 56706 33750
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56442 33674 56706 33684
rect 93262 33740 93526 33750
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93262 33674 93526 33684
rect 130082 33740 130346 33750
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130082 33674 130346 33684
rect 134204 33348 134260 33358
rect 38032 32956 38296 32966
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38032 32890 38296 32900
rect 74852 32956 75116 32966
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 74852 32890 75116 32900
rect 111672 32956 111936 32966
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111672 32890 111936 32900
rect 19622 32172 19886 32182
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19622 32106 19886 32116
rect 56442 32172 56706 32182
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56442 32106 56706 32116
rect 93262 32172 93526 32182
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93262 32106 93526 32116
rect 130082 32172 130346 32182
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130082 32106 130346 32116
rect 38032 31388 38296 31398
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38032 31322 38296 31332
rect 74852 31388 75116 31398
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 74852 31322 75116 31332
rect 111672 31388 111936 31398
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111672 31322 111936 31332
rect 131404 30996 131460 31006
rect 19622 30604 19886 30614
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19622 30538 19886 30548
rect 56442 30604 56706 30614
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56442 30538 56706 30548
rect 93262 30604 93526 30614
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93262 30538 93526 30548
rect 130082 30604 130346 30614
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130082 30538 130346 30548
rect 38032 29820 38296 29830
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38032 29754 38296 29764
rect 74852 29820 75116 29830
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 74852 29754 75116 29764
rect 111672 29820 111936 29830
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111672 29754 111936 29764
rect 128268 29428 128324 29438
rect 19622 29036 19886 29046
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19622 28970 19886 28980
rect 56442 29036 56706 29046
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56442 28970 56706 28980
rect 93262 29036 93526 29046
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93262 28970 93526 28980
rect 38032 28252 38296 28262
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38032 28186 38296 28196
rect 74852 28252 75116 28262
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 74852 28186 75116 28196
rect 111672 28252 111936 28262
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111672 28186 111936 28196
rect 126252 27748 126308 27758
rect 19622 27468 19886 27478
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19622 27402 19886 27412
rect 56442 27468 56706 27478
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56442 27402 56706 27412
rect 93262 27468 93526 27478
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93262 27402 93526 27412
rect 38032 26684 38296 26694
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38032 26618 38296 26628
rect 74852 26684 75116 26694
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 74852 26618 75116 26628
rect 111672 26684 111936 26694
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111672 26618 111936 26628
rect 19622 25900 19886 25910
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19622 25834 19886 25844
rect 56442 25900 56706 25910
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56442 25834 56706 25844
rect 93262 25900 93526 25910
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93262 25834 93526 25844
rect 123452 25284 123508 25294
rect 38032 25116 38296 25126
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38032 25050 38296 25060
rect 74852 25116 75116 25126
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 74852 25050 75116 25060
rect 111672 25116 111936 25126
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111672 25050 111936 25060
rect 19622 24332 19886 24342
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19622 24266 19886 24276
rect 56442 24332 56706 24342
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56442 24266 56706 24276
rect 93262 24332 93526 24342
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93262 24266 93526 24276
rect 38032 23548 38296 23558
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38032 23482 38296 23492
rect 74852 23548 75116 23558
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 74852 23482 75116 23492
rect 111672 23548 111936 23558
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111672 23482 111936 23492
rect 121884 23156 121940 23166
rect 19622 22764 19886 22774
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19622 22698 19886 22708
rect 56442 22764 56706 22774
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56442 22698 56706 22708
rect 93262 22764 93526 22774
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93262 22698 93526 22708
rect 115164 22372 115220 22382
rect 38032 21980 38296 21990
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38032 21914 38296 21924
rect 74852 21980 75116 21990
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 74852 21914 75116 21924
rect 111672 21980 111936 21990
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111672 21914 111936 21924
rect 19622 21196 19886 21206
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19622 21130 19886 21140
rect 56442 21196 56706 21206
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56442 21130 56706 21140
rect 93262 21196 93526 21206
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93262 21130 93526 21140
rect 114044 20804 114100 20814
rect 38032 20412 38296 20422
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38032 20346 38296 20356
rect 74852 20412 75116 20422
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 74852 20346 75116 20356
rect 111672 20412 111936 20422
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111672 20346 111936 20356
rect 19622 19628 19886 19638
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19622 19562 19886 19572
rect 56442 19628 56706 19638
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56442 19562 56706 19572
rect 93262 19628 93526 19638
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93262 19562 93526 19572
rect 110348 19236 110404 19246
rect 38032 18844 38296 18854
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38032 18778 38296 18788
rect 74852 18844 75116 18854
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 74852 18778 75116 18788
rect 106764 18340 106820 18350
rect 19622 18060 19886 18070
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19622 17994 19886 18004
rect 56442 18060 56706 18070
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56442 17994 56706 18004
rect 93262 18060 93526 18070
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93262 17994 93526 18004
rect 38032 17276 38296 17286
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38032 17210 38296 17220
rect 74852 17276 75116 17286
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 74852 17210 75116 17220
rect 19622 16492 19886 16502
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19622 16426 19886 16436
rect 56442 16492 56706 16502
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56442 16426 56706 16436
rect 93262 16492 93526 16502
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93262 16426 93526 16436
rect 38032 15708 38296 15718
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38032 15642 38296 15652
rect 74852 15708 75116 15718
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 74852 15642 75116 15652
rect 101836 15428 101892 15438
rect 19622 14924 19886 14934
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19622 14858 19886 14868
rect 56442 14924 56706 14934
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56442 14858 56706 14868
rect 93262 14924 93526 14934
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93262 14858 93526 14868
rect 100716 14532 100772 14542
rect 38032 14140 38296 14150
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38032 14074 38296 14084
rect 74852 14140 75116 14150
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 74852 14074 75116 14084
rect 19622 13356 19886 13366
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19622 13290 19886 13300
rect 56442 13356 56706 13366
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56442 13290 56706 13300
rect 93262 13356 93526 13366
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93262 13290 93526 13300
rect 99820 12964 99876 12974
rect 38032 12572 38296 12582
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38032 12506 38296 12516
rect 74852 12572 75116 12582
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 74852 12506 75116 12516
rect 19622 11788 19886 11798
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19622 11722 19886 11732
rect 56442 11788 56706 11798
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56442 11722 56706 11732
rect 93262 11788 93526 11798
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93262 11722 93526 11732
rect 98924 11284 98980 11294
rect 38032 11004 38296 11014
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38032 10938 38296 10948
rect 74852 11004 75116 11014
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 74852 10938 75116 10948
rect 59500 10500 59556 10510
rect 42700 10388 42756 10398
rect 19622 10220 19886 10230
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19622 10154 19886 10164
rect 38032 9436 38296 9446
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38032 9370 38296 9380
rect 41356 9044 41412 9054
rect 15148 8932 15204 8942
rect 13468 7364 13524 7374
rect 11788 5908 11844 5918
rect 10108 5796 10164 5806
rect 9660 5124 9716 5134
rect 8316 4340 8372 4350
rect 8316 4246 8372 4284
rect 8876 4340 8932 4350
rect 8876 4246 8932 4284
rect 9660 4340 9716 5068
rect 9660 4274 9716 4284
rect 9772 4564 9828 4574
rect 10108 4564 10164 5740
rect 9772 4562 10164 4564
rect 9772 4510 9774 4562
rect 9826 4510 10164 4562
rect 9772 4508 10164 4510
rect 11004 4564 11060 4574
rect 6636 4228 6692 4238
rect 7308 4228 7364 4238
rect 6636 3556 6692 4172
rect 6972 4226 7364 4228
rect 6972 4174 7310 4226
rect 7362 4174 7364 4226
rect 6972 4172 7364 4174
rect 6748 3556 6804 3566
rect 6636 3554 6804 3556
rect 6636 3502 6750 3554
rect 6802 3502 6804 3554
rect 6636 3500 6804 3502
rect 6748 3490 6804 3500
rect 5180 3444 5236 3454
rect 5180 800 5236 3388
rect 6076 3444 6132 3454
rect 6076 3350 6132 3388
rect 6972 980 7028 4172
rect 7308 4162 7364 4172
rect 8204 3668 8260 3678
rect 8204 3666 8596 3668
rect 8204 3614 8206 3666
rect 8258 3614 8596 3666
rect 8204 3612 8596 3614
rect 8204 3602 8260 3612
rect 6860 924 7028 980
rect 6860 800 6916 924
rect 8540 800 8596 3612
rect 8876 3556 8932 3566
rect 8876 3462 8932 3500
rect 9772 3556 9828 4508
rect 9772 3490 9828 3500
rect 10220 3666 10276 3678
rect 10220 3614 10222 3666
rect 10274 3614 10276 3666
rect 10220 800 10276 3614
rect 11004 3554 11060 4508
rect 11340 4564 11396 4574
rect 11340 4470 11396 4508
rect 11788 4564 11844 5852
rect 11788 4498 11844 4508
rect 13020 4564 13076 4574
rect 11004 3502 11006 3554
rect 11058 3502 11060 3554
rect 11004 3490 11060 3502
rect 12796 3556 12852 3566
rect 13020 3556 13076 4508
rect 13468 4564 13524 7308
rect 13468 4498 13524 4508
rect 15148 4562 15204 8876
rect 15148 4510 15150 4562
rect 15202 4510 15204 4562
rect 13916 3668 13972 3678
rect 12796 3554 13076 3556
rect 12796 3502 12798 3554
rect 12850 3502 13076 3554
rect 12796 3500 13076 3502
rect 13580 3666 13972 3668
rect 13580 3614 13918 3666
rect 13970 3614 13972 3666
rect 13580 3612 13972 3614
rect 12796 3490 12852 3500
rect 11900 3442 11956 3454
rect 11900 3390 11902 3442
rect 11954 3390 11956 3442
rect 11900 800 11956 3390
rect 13580 800 13636 3612
rect 13916 3602 13972 3612
rect 14924 3556 14980 3566
rect 15148 3556 15204 4510
rect 17500 8820 17556 8830
rect 16940 4228 16996 4238
rect 14924 3554 15204 3556
rect 14924 3502 14926 3554
rect 14978 3502 15204 3554
rect 14924 3500 15204 3502
rect 16716 3556 16772 3566
rect 14924 3490 14980 3500
rect 16716 3462 16772 3500
rect 15260 3444 15316 3454
rect 15260 800 15316 3388
rect 15820 3444 15876 3454
rect 15820 3350 15876 3388
rect 16940 800 16996 4172
rect 17500 3666 17556 8764
rect 19622 8652 19886 8662
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19622 8586 19886 8596
rect 38032 7868 38296 7878
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38032 7802 38296 7812
rect 39116 7588 39172 7598
rect 21644 7252 21700 7262
rect 19622 7084 19886 7094
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19622 7018 19886 7028
rect 19622 5516 19886 5526
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19622 5450 19886 5460
rect 18956 4452 19012 4462
rect 18956 4338 19012 4396
rect 19404 4452 19460 4462
rect 19404 4358 19460 4396
rect 18956 4286 18958 4338
rect 19010 4286 19012 4338
rect 18956 4274 19012 4286
rect 17948 4228 18004 4238
rect 17948 4134 18004 4172
rect 19622 3948 19886 3958
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19622 3882 19886 3892
rect 17500 3614 17502 3666
rect 17554 3614 17556 3666
rect 17500 3556 17556 3614
rect 17500 3490 17556 3500
rect 20076 3556 20132 3566
rect 20076 3462 20132 3500
rect 20636 3556 20692 3566
rect 20636 3462 20692 3500
rect 21644 3556 21700 7196
rect 22540 6804 22596 6814
rect 22540 4562 22596 6748
rect 35980 6580 36036 6590
rect 22540 4510 22542 4562
rect 22594 4510 22596 4562
rect 22540 4498 22596 4510
rect 30716 5684 30772 5694
rect 22204 4338 22260 4350
rect 22204 4286 22206 4338
rect 22258 4286 22260 4338
rect 21756 4228 21812 4238
rect 22204 4228 22260 4286
rect 21756 4226 22260 4228
rect 21756 4174 21758 4226
rect 21810 4174 22260 4226
rect 21756 4172 22260 4174
rect 22988 4226 23044 4238
rect 22988 4174 22990 4226
rect 23042 4174 23044 4226
rect 21756 4162 21812 4172
rect 21644 3490 21700 3500
rect 18620 3444 18676 3454
rect 18620 800 18676 3388
rect 19180 3444 19236 3454
rect 19180 3350 19236 3388
rect 20300 3444 20356 3454
rect 20300 800 20356 3388
rect 21756 3444 21812 3454
rect 21756 3350 21812 3388
rect 21980 800 22036 4172
rect 22652 3668 22708 3678
rect 22652 3554 22708 3612
rect 22988 3668 23044 4174
rect 22988 3602 23044 3612
rect 25564 4226 25620 4238
rect 25564 4174 25566 4226
rect 25618 4174 25620 4226
rect 22652 3502 22654 3554
rect 22706 3502 22708 3554
rect 22652 3490 22708 3502
rect 23436 3444 23492 3454
rect 23884 3444 23940 3454
rect 25564 3444 25620 4174
rect 23436 3442 23940 3444
rect 23436 3390 23438 3442
rect 23490 3390 23886 3442
rect 23938 3390 23940 3442
rect 23436 3388 23940 3390
rect 23436 3378 23492 3388
rect 23660 800 23716 3388
rect 23884 3378 23940 3388
rect 25340 3442 25620 3444
rect 25340 3390 25566 3442
rect 25618 3390 25620 3442
rect 25340 3388 25620 3390
rect 24220 3330 24276 3342
rect 24220 3278 24222 3330
rect 24274 3278 24276 3330
rect 24220 1540 24276 3278
rect 24220 1474 24276 1484
rect 25340 800 25396 3388
rect 25564 3378 25620 3388
rect 26796 3444 26852 3454
rect 27244 3444 27300 3454
rect 26796 3442 27300 3444
rect 26796 3390 26798 3442
rect 26850 3390 27246 3442
rect 27298 3390 27300 3442
rect 26796 3388 27300 3390
rect 26796 3378 26852 3388
rect 25900 3332 25956 3342
rect 25900 3238 25956 3276
rect 27020 800 27076 3388
rect 27244 3378 27300 3388
rect 28588 3444 28644 3454
rect 28700 3444 28756 3454
rect 28588 3442 28700 3444
rect 28588 3390 28590 3442
rect 28642 3390 28700 3442
rect 28588 3388 28700 3390
rect 28588 3378 28644 3388
rect 27580 3330 27636 3342
rect 27580 3278 27582 3330
rect 27634 3278 27636 3330
rect 27580 2996 27636 3278
rect 27580 2930 27636 2940
rect 28700 800 28756 3388
rect 29260 3444 29316 3454
rect 29260 3350 29316 3388
rect 30156 3444 30212 3454
rect 30604 3444 30660 3454
rect 30156 3442 30660 3444
rect 30156 3390 30158 3442
rect 30210 3390 30606 3442
rect 30658 3390 30660 3442
rect 30156 3388 30660 3390
rect 30156 3378 30212 3388
rect 29596 3330 29652 3342
rect 29596 3278 29598 3330
rect 29650 3278 29652 3330
rect 29596 2884 29652 3278
rect 29596 2818 29652 2828
rect 30380 800 30436 3388
rect 30604 3378 30660 3388
rect 30716 3332 30772 5628
rect 32060 4228 32116 4238
rect 32060 3442 32116 4172
rect 32620 4228 32676 4238
rect 32620 4134 32676 4172
rect 32060 3390 32062 3442
rect 32114 3390 32116 3442
rect 30716 3266 30772 3276
rect 30940 3330 30996 3342
rect 30940 3278 30942 3330
rect 30994 3278 30996 3330
rect 30940 2772 30996 3278
rect 30940 2706 30996 2716
rect 32060 800 32116 3390
rect 33516 3444 33572 3454
rect 33964 3444 34020 3454
rect 33516 3442 34020 3444
rect 33516 3390 33518 3442
rect 33570 3390 33966 3442
rect 34018 3390 34020 3442
rect 33516 3388 34020 3390
rect 33516 3378 33572 3388
rect 32396 3330 32452 3342
rect 32396 3278 32398 3330
rect 32450 3278 32452 3330
rect 32396 2548 32452 3278
rect 32396 2482 32452 2492
rect 33740 800 33796 3388
rect 33964 3378 34020 3388
rect 35196 3444 35252 3454
rect 35644 3444 35700 3454
rect 35196 3442 35700 3444
rect 35196 3390 35198 3442
rect 35250 3390 35646 3442
rect 35698 3390 35700 3442
rect 35196 3388 35700 3390
rect 35196 3378 35252 3388
rect 34300 3330 34356 3342
rect 34300 3278 34302 3330
rect 34354 3278 34356 3330
rect 34300 2436 34356 3278
rect 34300 2370 34356 2380
rect 35420 800 35476 3388
rect 35644 3378 35700 3388
rect 35980 3330 36036 6524
rect 38032 6300 38296 6310
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38032 6234 38296 6244
rect 38032 4732 38296 4742
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38032 4666 38296 4676
rect 35980 3278 35982 3330
rect 36034 3278 36036 3330
rect 35980 3266 36036 3278
rect 37100 4226 37156 4238
rect 37100 4174 37102 4226
rect 37154 4174 37156 4226
rect 37100 3444 37156 4174
rect 37324 3444 37380 3454
rect 37100 3442 37380 3444
rect 37100 3390 37326 3442
rect 37378 3390 37380 3442
rect 37100 3388 37380 3390
rect 37100 800 37156 3388
rect 37324 3378 37380 3388
rect 38556 3444 38612 3454
rect 39004 3444 39060 3454
rect 38556 3442 39060 3444
rect 38556 3390 38558 3442
rect 38610 3390 39006 3442
rect 39058 3390 39060 3442
rect 38556 3388 39060 3390
rect 38556 3378 38612 3388
rect 37660 3332 37716 3342
rect 37660 3238 37716 3276
rect 38032 3164 38296 3174
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38032 3098 38296 3108
rect 38780 800 38836 3388
rect 39004 3378 39060 3388
rect 39116 3332 39172 7532
rect 40348 3444 40404 3454
rect 40460 3444 40516 3454
rect 40348 3442 40460 3444
rect 40348 3390 40350 3442
rect 40402 3390 40460 3442
rect 40348 3388 40460 3390
rect 40348 3378 40404 3388
rect 39116 3266 39172 3276
rect 39340 3332 39396 3342
rect 39340 3238 39396 3276
rect 40460 800 40516 3388
rect 41020 3444 41076 3454
rect 41020 3350 41076 3388
rect 41356 3330 41412 8988
rect 42476 4564 42532 4574
rect 41916 3444 41972 3454
rect 42364 3444 42420 3454
rect 41916 3442 42420 3444
rect 41916 3390 41918 3442
rect 41970 3390 42366 3442
rect 42418 3390 42420 3442
rect 41916 3388 42420 3390
rect 41916 3378 41972 3388
rect 41356 3278 41358 3330
rect 41410 3278 41412 3330
rect 41356 3266 41412 3278
rect 42140 800 42196 3388
rect 42364 3378 42420 3388
rect 42476 3332 42532 4508
rect 42476 3266 42532 3276
rect 42700 3330 42756 10332
rect 56442 10220 56706 10230
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56442 10154 56706 10164
rect 56442 8652 56706 8662
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56442 8586 56706 8596
rect 53116 8484 53172 8494
rect 51100 7700 51156 7710
rect 42700 3278 42702 3330
rect 42754 3278 42756 3330
rect 42700 3266 42756 3278
rect 43820 4228 43876 4238
rect 43820 3442 43876 4172
rect 44380 4228 44436 4238
rect 44380 4134 44436 4172
rect 48860 4226 48916 4238
rect 48860 4174 48862 4226
rect 48914 4174 48916 4226
rect 43820 3390 43822 3442
rect 43874 3390 43876 3442
rect 43820 800 43876 3390
rect 45276 3444 45332 3454
rect 45724 3444 45780 3454
rect 45276 3442 45780 3444
rect 45276 3390 45278 3442
rect 45330 3390 45726 3442
rect 45778 3390 45780 3442
rect 45276 3388 45780 3390
rect 45276 3378 45332 3388
rect 44156 3330 44212 3342
rect 44156 3278 44158 3330
rect 44210 3278 44212 3330
rect 44156 1204 44212 3278
rect 44156 1138 44212 1148
rect 45500 800 45556 3388
rect 45724 3378 45780 3388
rect 46956 3444 47012 3454
rect 47404 3444 47460 3454
rect 46956 3442 47460 3444
rect 46956 3390 46958 3442
rect 47010 3390 47406 3442
rect 47458 3390 47460 3442
rect 46956 3388 47460 3390
rect 46956 3378 47012 3388
rect 46060 3330 46116 3342
rect 46060 3278 46062 3330
rect 46114 3278 46116 3330
rect 46060 1316 46116 3278
rect 46060 1250 46116 1260
rect 47180 800 47236 3388
rect 47404 3378 47460 3388
rect 48860 3444 48916 4174
rect 49084 3444 49140 3454
rect 48860 3442 49140 3444
rect 48860 3390 49086 3442
rect 49138 3390 49140 3442
rect 48860 3388 49140 3390
rect 47740 3330 47796 3342
rect 47740 3278 47742 3330
rect 47794 3278 47796 3330
rect 47740 868 47796 3278
rect 47740 802 47796 812
rect 48860 800 48916 3388
rect 49084 3378 49140 3388
rect 50316 3444 50372 3454
rect 50764 3444 50820 3454
rect 50316 3442 50820 3444
rect 50316 3390 50318 3442
rect 50370 3390 50766 3442
rect 50818 3390 50820 3442
rect 50316 3388 50820 3390
rect 50316 3378 50372 3388
rect 49420 3330 49476 3342
rect 49420 3278 49422 3330
rect 49474 3278 49476 3330
rect 49420 1428 49476 3278
rect 49420 1362 49476 1372
rect 50540 800 50596 3388
rect 50764 3378 50820 3388
rect 51100 3330 51156 7644
rect 52108 3444 52164 3454
rect 52220 3444 52276 3454
rect 52108 3442 52220 3444
rect 52108 3390 52110 3442
rect 52162 3390 52220 3442
rect 52108 3388 52220 3390
rect 52108 3378 52164 3388
rect 51100 3278 51102 3330
rect 51154 3278 51156 3330
rect 51100 3266 51156 3278
rect 52220 800 52276 3388
rect 52780 3444 52836 3454
rect 52780 3350 52836 3388
rect 53116 3330 53172 8428
rect 57260 7476 57316 7486
rect 56442 7084 56706 7094
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56442 7018 56706 7028
rect 56442 5516 56706 5526
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56442 5450 56706 5460
rect 55916 5348 55972 5358
rect 55580 4228 55636 4238
rect 54236 4116 54292 4126
rect 53676 3444 53732 3454
rect 54124 3444 54180 3454
rect 53676 3442 54180 3444
rect 53676 3390 53678 3442
rect 53730 3390 54126 3442
rect 54178 3390 54180 3442
rect 53676 3388 54180 3390
rect 53676 3378 53732 3388
rect 53116 3278 53118 3330
rect 53170 3278 53172 3330
rect 53116 3266 53172 3278
rect 53900 800 53956 3388
rect 54124 3378 54180 3388
rect 54236 2996 54292 4060
rect 55580 3442 55636 4172
rect 55580 3390 55582 3442
rect 55634 3390 55636 3442
rect 54460 3332 54516 3342
rect 54460 3238 54516 3276
rect 54236 2930 54292 2940
rect 55580 800 55636 3390
rect 55916 3330 55972 5292
rect 56140 4228 56196 4238
rect 56140 4134 56196 4172
rect 56442 3948 56706 3958
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56442 3882 56706 3892
rect 57260 3668 57316 7420
rect 57260 3602 57316 3612
rect 57036 3444 57092 3454
rect 57484 3444 57540 3454
rect 57036 3442 57540 3444
rect 57036 3390 57038 3442
rect 57090 3390 57486 3442
rect 57538 3390 57540 3442
rect 57036 3388 57540 3390
rect 57036 3378 57092 3388
rect 55916 3278 55918 3330
rect 55970 3278 55972 3330
rect 55916 3266 55972 3278
rect 56924 3332 56980 3342
rect 56924 1092 56980 3276
rect 56924 1026 56980 1036
rect 57260 800 57316 3388
rect 57484 3378 57540 3388
rect 58716 3444 58772 3454
rect 59164 3444 59220 3454
rect 58716 3442 59220 3444
rect 58716 3390 58718 3442
rect 58770 3390 59166 3442
rect 59218 3390 59220 3442
rect 58716 3388 59220 3390
rect 58716 3378 58772 3388
rect 57820 3332 57876 3342
rect 57820 3238 57876 3276
rect 58940 800 58996 3388
rect 59164 3378 59220 3388
rect 59500 3330 59556 10444
rect 93262 10220 93526 10230
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93262 10154 93526 10164
rect 74852 9436 75116 9446
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 74852 9370 75116 9380
rect 90748 9156 90804 9166
rect 82908 8932 82964 8942
rect 74852 7868 75116 7878
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 74852 7802 75116 7812
rect 80556 7364 80612 7374
rect 71260 6916 71316 6926
rect 61292 5236 61348 5246
rect 59500 3278 59502 3330
rect 59554 3278 59556 3330
rect 59500 3266 59556 3278
rect 60396 4900 60452 4910
rect 60396 2884 60452 4844
rect 61292 4452 61348 5180
rect 61292 4386 61348 4396
rect 60396 2818 60452 2828
rect 60620 4226 60676 4238
rect 60620 4174 60622 4226
rect 60674 4174 60676 4226
rect 60620 3444 60676 4174
rect 67340 4228 67396 4238
rect 66220 4004 66276 4014
rect 62636 3668 62692 3678
rect 60844 3444 60900 3454
rect 60620 3442 60900 3444
rect 60620 3390 60846 3442
rect 60898 3390 60900 3442
rect 60620 3388 60900 3390
rect 60620 800 60676 3388
rect 60844 3378 60900 3388
rect 62076 3444 62132 3454
rect 62524 3444 62580 3454
rect 62076 3442 62580 3444
rect 62076 3390 62078 3442
rect 62130 3390 62526 3442
rect 62578 3390 62580 3442
rect 62076 3388 62580 3390
rect 62076 3378 62132 3388
rect 61180 3330 61236 3342
rect 61180 3278 61182 3330
rect 61234 3278 61236 3330
rect 61180 2660 61236 3278
rect 61180 2594 61236 2604
rect 62300 800 62356 3388
rect 62524 3378 62580 3388
rect 62636 2548 62692 3612
rect 63868 3444 63924 3454
rect 63980 3444 64036 3454
rect 63868 3442 63980 3444
rect 63868 3390 63870 3442
rect 63922 3390 63980 3442
rect 63868 3388 63980 3390
rect 63868 3378 63924 3388
rect 62860 3330 62916 3342
rect 62860 3278 62862 3330
rect 62914 3278 62916 3330
rect 62860 2996 62916 3278
rect 62860 2930 62916 2940
rect 62636 2482 62692 2492
rect 63980 800 64036 3388
rect 64540 3444 64596 3454
rect 64540 3350 64596 3388
rect 65436 3444 65492 3454
rect 65884 3444 65940 3454
rect 65436 3442 65940 3444
rect 65436 3390 65438 3442
rect 65490 3390 65886 3442
rect 65938 3390 65940 3442
rect 65436 3388 65940 3390
rect 65436 3378 65492 3388
rect 64092 3332 64148 3342
rect 64092 980 64148 3276
rect 64876 3330 64932 3342
rect 64876 3278 64878 3330
rect 64930 3278 64932 3330
rect 64876 2548 64932 3278
rect 64876 2482 64932 2492
rect 64092 914 64148 924
rect 65660 800 65716 3388
rect 65884 3378 65940 3388
rect 66220 3330 66276 3948
rect 66220 3278 66222 3330
rect 66274 3278 66276 3330
rect 66220 3266 66276 3278
rect 67340 3442 67396 4172
rect 67900 4228 67956 4238
rect 67900 4134 67956 4172
rect 67340 3390 67342 3442
rect 67394 3390 67396 3442
rect 67340 800 67396 3390
rect 68796 3444 68852 3454
rect 69244 3444 69300 3454
rect 68796 3442 69300 3444
rect 68796 3390 68798 3442
rect 68850 3390 69246 3442
rect 69298 3390 69300 3442
rect 68796 3388 69300 3390
rect 68796 3378 68852 3388
rect 67676 3330 67732 3342
rect 67676 3278 67678 3330
rect 67730 3278 67732 3330
rect 67676 2100 67732 3278
rect 67676 2034 67732 2044
rect 69020 800 69076 3388
rect 69244 3378 69300 3388
rect 70476 3444 70532 3454
rect 70924 3444 70980 3454
rect 70476 3442 70980 3444
rect 70476 3390 70478 3442
rect 70530 3390 70926 3442
rect 70978 3390 70980 3442
rect 70476 3388 70980 3390
rect 70476 3378 70532 3388
rect 69580 3330 69636 3342
rect 69580 3278 69582 3330
rect 69634 3278 69636 3330
rect 69580 2212 69636 3278
rect 69580 2146 69636 2156
rect 70700 800 70756 3388
rect 70924 3378 70980 3388
rect 71260 3330 71316 6860
rect 77644 6692 77700 6702
rect 74852 6300 75116 6310
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 74852 6234 75116 6244
rect 76076 6244 76132 6254
rect 75180 5124 75236 5134
rect 74852 4732 75116 4742
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 74852 4666 75116 4676
rect 73948 4452 74004 4462
rect 73724 4396 73948 4452
rect 73388 4340 73444 4350
rect 72492 4228 72548 4238
rect 72492 3444 72548 4172
rect 73276 4228 73332 4238
rect 73276 4134 73332 4172
rect 71260 3278 71262 3330
rect 71314 3278 71316 3330
rect 71260 3266 71316 3278
rect 72380 3442 72548 3444
rect 72380 3390 72494 3442
rect 72546 3390 72548 3442
rect 72380 3388 72548 3390
rect 72380 800 72436 3388
rect 72492 3378 72548 3388
rect 72828 3780 72884 3790
rect 72828 3330 72884 3724
rect 72828 3278 72830 3330
rect 72882 3278 72884 3330
rect 72828 3266 72884 3278
rect 73388 3330 73444 4284
rect 73724 3554 73780 4396
rect 73948 4358 74004 4396
rect 74396 4228 74452 4238
rect 73724 3502 73726 3554
rect 73778 3502 73780 3554
rect 73724 3490 73780 3502
rect 74284 4226 74452 4228
rect 74284 4174 74398 4226
rect 74450 4174 74452 4226
rect 74284 4172 74452 4174
rect 74284 3444 74340 4172
rect 74396 4162 74452 4172
rect 73388 3278 73390 3330
rect 73442 3278 73444 3330
rect 73388 3266 73444 3278
rect 74060 3442 74340 3444
rect 74060 3390 74286 3442
rect 74338 3390 74340 3442
rect 74060 3388 74340 3390
rect 74060 800 74116 3388
rect 74284 3378 74340 3388
rect 74620 3330 74676 3342
rect 74620 3278 74622 3330
rect 74674 3278 74676 3330
rect 74620 2884 74676 3278
rect 75180 3330 75236 5068
rect 75852 5124 75908 5134
rect 75852 5030 75908 5068
rect 75516 5012 75572 5022
rect 75292 4452 75348 4462
rect 75292 4358 75348 4396
rect 75516 3554 75572 4956
rect 76076 4562 76132 6188
rect 77644 5234 77700 6636
rect 79660 5908 79716 5918
rect 77644 5182 77646 5234
rect 77698 5182 77700 5234
rect 76076 4510 76078 4562
rect 76130 4510 76132 4562
rect 75628 4452 75684 4462
rect 76076 4452 76132 4510
rect 75628 4450 75908 4452
rect 75628 4398 75630 4450
rect 75682 4398 75908 4450
rect 75628 4396 75908 4398
rect 75628 4386 75684 4396
rect 75516 3502 75518 3554
rect 75570 3502 75572 3554
rect 75516 3490 75572 3502
rect 75852 3556 75908 4396
rect 76076 4386 76132 4396
rect 76972 5124 77028 5134
rect 76972 4450 77028 5068
rect 77644 5124 77700 5182
rect 77644 5058 77700 5068
rect 77868 5796 77924 5806
rect 77868 4562 77924 5740
rect 77868 4510 77870 4562
rect 77922 4510 77924 4562
rect 77868 4498 77924 4510
rect 78204 5124 78260 5134
rect 76972 4398 76974 4450
rect 77026 4398 77028 4450
rect 76972 4386 77028 4398
rect 77308 4450 77364 4462
rect 77308 4398 77310 4450
rect 77362 4398 77364 4450
rect 76300 3556 76356 3566
rect 75852 3554 76356 3556
rect 75852 3502 76302 3554
rect 76354 3502 76356 3554
rect 75852 3500 76356 3502
rect 77308 3556 77364 4398
rect 78204 4450 78260 5068
rect 78540 5124 78596 5134
rect 78540 5030 78596 5068
rect 78876 5124 78932 5134
rect 78204 4398 78206 4450
rect 78258 4398 78260 4450
rect 78204 4386 78260 4398
rect 78876 4338 78932 5068
rect 79436 5124 79492 5134
rect 79436 5030 79492 5068
rect 79660 4562 79716 5852
rect 80556 5010 80612 7308
rect 82236 7364 82292 7374
rect 82124 5122 82180 5134
rect 82124 5070 82126 5122
rect 82178 5070 82180 5122
rect 80556 4958 80558 5010
rect 80610 4958 80612 5010
rect 80556 4946 80612 4958
rect 80892 5010 80948 5022
rect 80892 4958 80894 5010
rect 80946 4958 80948 5010
rect 80892 4788 80948 4958
rect 80892 4722 80948 4732
rect 81340 4898 81396 4910
rect 81340 4846 81342 4898
rect 81394 4846 81396 4898
rect 81340 4788 81396 4846
rect 81340 4722 81396 4732
rect 82124 4788 82180 5070
rect 82124 4722 82180 4732
rect 79660 4510 79662 4562
rect 79714 4510 79716 4562
rect 79660 4498 79716 4510
rect 82124 4564 82180 4574
rect 82236 4564 82292 7308
rect 82684 5794 82740 5806
rect 82684 5742 82686 5794
rect 82738 5742 82740 5794
rect 82124 4562 82292 4564
rect 82124 4510 82126 4562
rect 82178 4510 82292 4562
rect 82124 4508 82292 4510
rect 82348 4898 82404 4910
rect 82348 4846 82350 4898
rect 82402 4846 82404 4898
rect 79100 4452 79156 4462
rect 79996 4452 80052 4462
rect 79100 4450 79268 4452
rect 79100 4398 79102 4450
rect 79154 4398 79268 4450
rect 79100 4396 79268 4398
rect 79100 4386 79156 4396
rect 78876 4286 78878 4338
rect 78930 4286 78932 4338
rect 78764 3666 78820 3678
rect 78764 3614 78766 3666
rect 78818 3614 78820 3666
rect 78092 3556 78148 3566
rect 77308 3554 78148 3556
rect 77308 3502 78094 3554
rect 78146 3502 78148 3554
rect 77308 3500 78148 3502
rect 76300 3490 76356 3500
rect 78092 3490 78148 3500
rect 75180 3278 75182 3330
rect 75234 3278 75236 3330
rect 75180 3266 75236 3278
rect 75740 3444 75796 3454
rect 74852 3164 75116 3174
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 74852 3098 75116 3108
rect 74620 2818 74676 2828
rect 75740 800 75796 3388
rect 77196 3444 77252 3454
rect 77196 3350 77252 3388
rect 78764 3444 78820 3614
rect 78764 3378 78820 3388
rect 77420 3332 77476 3342
rect 77420 800 77476 3276
rect 78876 868 78932 4286
rect 79212 3556 79268 4396
rect 79996 4358 80052 4396
rect 80444 4452 80500 4462
rect 80444 4358 80500 4396
rect 81340 4452 81396 4462
rect 81340 4358 81396 4396
rect 81676 4450 81732 4462
rect 81676 4398 81678 4450
rect 81730 4398 81732 4450
rect 80220 3556 80276 3566
rect 79212 3554 80276 3556
rect 79212 3502 80222 3554
rect 80274 3502 80276 3554
rect 79212 3500 80276 3502
rect 80220 3490 80276 3500
rect 80780 3556 80836 3566
rect 81676 3556 81732 4398
rect 82124 4452 82180 4508
rect 82124 4386 82180 4396
rect 82348 4340 82404 4846
rect 82684 4788 82740 5742
rect 82908 5010 82964 8876
rect 83916 8820 83972 8830
rect 83580 5794 83636 5806
rect 83580 5742 83582 5794
rect 83634 5742 83636 5794
rect 83244 5124 83300 5134
rect 83244 5030 83300 5068
rect 83580 5124 83636 5742
rect 83580 5058 83636 5068
rect 82908 4958 82910 5010
rect 82962 4958 82964 5010
rect 82908 4946 82964 4958
rect 83916 5010 83972 8764
rect 90524 8820 90580 8830
rect 88956 7476 89012 7486
rect 87276 7252 87332 7262
rect 84476 6356 84532 6366
rect 84476 6132 84532 6300
rect 84252 6130 84532 6132
rect 84252 6078 84478 6130
rect 84530 6078 84532 6130
rect 84252 6076 84532 6078
rect 84252 5122 84308 6076
rect 84476 6066 84532 6076
rect 86940 6356 86996 6366
rect 85372 6020 85428 6030
rect 84252 5070 84254 5122
rect 84306 5070 84308 5122
rect 84252 5058 84308 5070
rect 84588 5124 84644 5134
rect 83916 4958 83918 5010
rect 83970 4958 83972 5010
rect 83916 4946 83972 4958
rect 82684 4722 82740 4732
rect 82684 4340 82740 4350
rect 82348 4338 82740 4340
rect 82348 4286 82686 4338
rect 82738 4286 82740 4338
rect 82348 4284 82740 4286
rect 82684 4274 82740 4284
rect 84588 4338 84644 5068
rect 85372 5124 85428 5964
rect 85372 4562 85428 5068
rect 85596 5236 85652 5246
rect 85596 5010 85652 5180
rect 85596 4958 85598 5010
rect 85650 4958 85652 5010
rect 85596 4946 85652 4958
rect 85932 5010 85988 5022
rect 85932 4958 85934 5010
rect 85986 4958 85988 5010
rect 85932 4900 85988 4958
rect 85932 4834 85988 4844
rect 86380 4900 86436 4910
rect 86380 4806 86436 4844
rect 85372 4510 85374 4562
rect 85426 4510 85428 4562
rect 85372 4498 85428 4510
rect 84588 4286 84590 4338
rect 84642 4286 84644 4338
rect 84588 4274 84644 4286
rect 84812 4450 84868 4462
rect 84812 4398 84814 4450
rect 84866 4398 84868 4450
rect 83356 4226 83412 4238
rect 83356 4174 83358 4226
rect 83410 4174 83412 4226
rect 82684 3666 82740 3678
rect 82684 3614 82686 3666
rect 82738 3614 82740 3666
rect 82012 3556 82068 3566
rect 81676 3554 82068 3556
rect 81676 3502 82014 3554
rect 82066 3502 82068 3554
rect 81676 3500 82068 3502
rect 78876 802 78932 812
rect 79100 3444 79156 3454
rect 79100 800 79156 3388
rect 80780 800 80836 3500
rect 82012 3490 82068 3500
rect 82684 3556 82740 3614
rect 82684 3490 82740 3500
rect 81116 3444 81172 3454
rect 81116 3350 81172 3388
rect 82460 3444 82516 3454
rect 82460 800 82516 3388
rect 83356 3444 83412 4174
rect 84812 3556 84868 4398
rect 86156 4338 86212 4350
rect 86156 4286 86158 4338
rect 86210 4286 86212 4338
rect 85820 4228 85876 4238
rect 85372 3556 85428 3566
rect 84812 3554 85428 3556
rect 84812 3502 85374 3554
rect 85426 3502 85428 3554
rect 84812 3500 85428 3502
rect 85372 3490 85428 3500
rect 83356 3378 83412 3388
rect 84140 3444 84196 3454
rect 84140 800 84196 3388
rect 84700 3444 84756 3454
rect 84700 3350 84756 3388
rect 85820 800 85876 4172
rect 86156 3442 86212 4286
rect 86716 4228 86772 4238
rect 86716 4134 86772 4172
rect 86940 3668 86996 6300
rect 87276 5010 87332 7196
rect 88396 7252 88452 7262
rect 88396 6132 88452 7196
rect 87948 6130 88452 6132
rect 87948 6078 88398 6130
rect 88450 6078 88452 6130
rect 87948 6076 88452 6078
rect 87612 5236 87668 5246
rect 87612 5122 87668 5180
rect 87612 5070 87614 5122
rect 87666 5070 87668 5122
rect 87612 5058 87668 5070
rect 87276 4958 87278 5010
rect 87330 4958 87332 5010
rect 87276 4946 87332 4958
rect 87948 4900 88004 6076
rect 88396 6066 88452 6076
rect 88060 5236 88116 5246
rect 88060 5142 88116 5180
rect 88956 5010 89012 7420
rect 89404 5236 89460 5246
rect 88956 4958 88958 5010
rect 89010 4958 89012 5010
rect 88956 4946 89012 4958
rect 89292 5010 89348 5022
rect 89292 4958 89294 5010
rect 89346 4958 89348 5010
rect 87948 4338 88004 4844
rect 89292 4900 89348 4958
rect 89292 4834 89348 4844
rect 87948 4286 87950 4338
rect 88002 4286 88004 4338
rect 87948 4274 88004 4286
rect 88172 4450 88228 4462
rect 88172 4398 88174 4450
rect 88226 4398 88228 4450
rect 86492 3666 86996 3668
rect 86492 3614 86942 3666
rect 86994 3614 86996 3666
rect 86492 3612 86996 3614
rect 86492 3554 86548 3612
rect 86940 3602 86996 3612
rect 86492 3502 86494 3554
rect 86546 3502 86548 3554
rect 86492 3490 86548 3502
rect 88172 3554 88228 4398
rect 89404 4338 89460 5180
rect 90188 5236 90244 5246
rect 90188 5142 90244 5180
rect 89740 4900 89796 4910
rect 89740 4806 89796 4844
rect 90524 4900 90580 8764
rect 90748 5236 90804 9100
rect 93262 8652 93526 8662
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93262 8586 93526 8596
rect 93262 7084 93526 7094
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93262 7018 93526 7028
rect 97132 5684 97188 5694
rect 93262 5516 93526 5526
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93262 5450 93526 5460
rect 90748 5170 90804 5180
rect 89404 4286 89406 4338
rect 89458 4286 89460 4338
rect 89404 4274 89460 4286
rect 89628 4450 89684 4462
rect 89628 4398 89630 4450
rect 89682 4398 89684 4450
rect 88172 3502 88174 3554
rect 88226 3502 88228 3554
rect 88172 3490 88228 3502
rect 89628 3556 89684 4398
rect 90524 4452 90580 4844
rect 90524 4338 90580 4396
rect 90524 4286 90526 4338
rect 90578 4286 90580 4338
rect 90524 4274 90580 4286
rect 90748 4450 90804 4462
rect 90748 4398 90750 4450
rect 90802 4398 90804 4450
rect 90524 3666 90580 3678
rect 90524 3614 90526 3666
rect 90578 3614 90580 3666
rect 89852 3556 89908 3566
rect 89628 3554 89908 3556
rect 89628 3502 89854 3554
rect 89906 3502 89908 3554
rect 89628 3500 89908 3502
rect 89852 3490 89908 3500
rect 86156 3390 86158 3442
rect 86210 3390 86212 3442
rect 86156 3378 86212 3390
rect 87500 3444 87556 3454
rect 87500 800 87556 3388
rect 88956 3444 89012 3454
rect 88956 3350 89012 3388
rect 89180 3444 89236 3454
rect 89180 800 89236 3388
rect 90524 3444 90580 3614
rect 90748 3556 90804 4398
rect 91308 4452 91364 4462
rect 91308 4358 91364 4396
rect 93548 4228 93604 4238
rect 93548 4226 93716 4228
rect 93548 4174 93550 4226
rect 93602 4174 93716 4226
rect 93548 4172 93716 4174
rect 93548 4162 93604 4172
rect 93262 3948 93526 3958
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93262 3882 93526 3892
rect 91980 3556 92036 3566
rect 90748 3554 92036 3556
rect 90748 3502 91982 3554
rect 92034 3502 92036 3554
rect 90748 3500 92036 3502
rect 91980 3490 92036 3500
rect 92540 3556 92596 3566
rect 93660 3556 93716 4172
rect 94444 4226 94500 4238
rect 94444 4174 94446 4226
rect 94498 4174 94500 4226
rect 93772 3556 93828 3566
rect 93660 3500 93772 3556
rect 90524 3378 90580 3388
rect 90860 3332 90916 3342
rect 90860 800 90916 3276
rect 92540 800 92596 3500
rect 93772 3462 93828 3500
rect 92876 3444 92932 3454
rect 94444 3444 94500 4174
rect 95900 4226 95956 4238
rect 95900 4174 95902 4226
rect 95954 4174 95956 4226
rect 94668 3444 94724 3454
rect 92876 3350 92932 3388
rect 94220 3442 94724 3444
rect 94220 3390 94670 3442
rect 94722 3390 94724 3442
rect 94220 3388 94724 3390
rect 94108 3330 94164 3342
rect 94108 3278 94110 3330
rect 94162 3278 94164 3330
rect 94108 2324 94164 3278
rect 94108 2258 94164 2268
rect 94220 800 94276 3388
rect 94668 3378 94724 3388
rect 95900 3444 95956 4174
rect 97132 3666 97188 5628
rect 98364 5122 98420 5134
rect 98364 5070 98366 5122
rect 98418 5070 98420 5122
rect 97580 4900 97636 4910
rect 97356 4340 97412 4350
rect 97580 4340 97636 4844
rect 98028 4898 98084 4910
rect 98028 4846 98030 4898
rect 98082 4846 98084 4898
rect 97692 4452 97748 4462
rect 98028 4452 98084 4846
rect 98364 4900 98420 5070
rect 98364 4834 98420 4844
rect 98476 4452 98532 4462
rect 98028 4450 98532 4452
rect 98028 4398 98478 4450
rect 98530 4398 98532 4450
rect 98028 4396 98532 4398
rect 97692 4358 97748 4396
rect 97356 4338 97636 4340
rect 97356 4286 97358 4338
rect 97410 4286 97636 4338
rect 97356 4284 97636 4286
rect 97356 4274 97412 4284
rect 97132 3614 97134 3666
rect 97186 3614 97188 3666
rect 96460 3556 96516 3566
rect 96124 3444 96180 3454
rect 95900 3442 96180 3444
rect 95900 3390 96126 3442
rect 96178 3390 96180 3442
rect 95900 3388 96180 3390
rect 95004 3332 95060 3342
rect 95004 3238 95060 3276
rect 95676 2772 95732 2782
rect 95676 1652 95732 2716
rect 95676 1586 95732 1596
rect 95900 800 95956 3388
rect 96124 3378 96180 3388
rect 96460 3330 96516 3500
rect 97132 3444 97188 3614
rect 97132 3378 97188 3388
rect 96460 3278 96462 3330
rect 96514 3278 96516 3330
rect 96460 3266 96516 3278
rect 97580 800 97636 4284
rect 98364 4228 98420 4238
rect 97804 3444 97860 3454
rect 97804 3350 97860 3388
rect 98364 3442 98420 4172
rect 98364 3390 98366 3442
rect 98418 3390 98420 3442
rect 98364 3378 98420 3390
rect 98476 1540 98532 4396
rect 98700 4338 98756 4350
rect 98700 4286 98702 4338
rect 98754 4286 98756 4338
rect 98700 4228 98756 4286
rect 98700 4162 98756 4172
rect 98924 3778 98980 11228
rect 99484 11284 99540 11294
rect 99484 11190 99540 11228
rect 99820 11282 99876 12908
rect 100716 12402 100772 14476
rect 100716 12350 100718 12402
rect 100770 12350 100772 12402
rect 100716 12338 100772 12350
rect 101500 12850 101556 12862
rect 101500 12798 101502 12850
rect 101554 12798 101556 12850
rect 100492 12178 100548 12190
rect 100492 12126 100494 12178
rect 100546 12126 100548 12178
rect 100492 12068 100548 12126
rect 101164 12068 101220 12078
rect 100492 12066 101220 12068
rect 100492 12014 101166 12066
rect 101218 12014 101220 12066
rect 100492 12012 101220 12014
rect 99820 11230 99822 11282
rect 99874 11230 99876 11282
rect 99820 11218 99876 11230
rect 99596 10164 99652 10174
rect 99596 7698 99652 10108
rect 99596 7646 99598 7698
rect 99650 7646 99652 7698
rect 99596 7634 99652 7646
rect 99372 7474 99428 7486
rect 99372 7422 99374 7474
rect 99426 7422 99428 7474
rect 99036 5124 99092 5134
rect 99260 5124 99316 5134
rect 99036 5122 99260 5124
rect 99036 5070 99038 5122
rect 99090 5070 99260 5122
rect 99036 5068 99260 5070
rect 99036 5058 99092 5068
rect 98924 3726 98926 3778
rect 98978 3726 98980 3778
rect 98924 3714 98980 3726
rect 99148 4114 99204 4126
rect 99148 4062 99150 4114
rect 99202 4062 99204 4114
rect 98588 3556 98644 3566
rect 98588 3462 98644 3500
rect 99148 3332 99204 4062
rect 99148 3266 99204 3276
rect 98476 1474 98532 1484
rect 99260 800 99316 5068
rect 99372 4564 99428 7422
rect 99596 5794 99652 5806
rect 99596 5742 99598 5794
rect 99650 5742 99652 5794
rect 99484 5124 99540 5134
rect 99484 5010 99540 5068
rect 99484 4958 99486 5010
rect 99538 4958 99540 5010
rect 99484 4946 99540 4958
rect 99484 4564 99540 4574
rect 99372 4562 99540 4564
rect 99372 4510 99486 4562
rect 99538 4510 99540 4562
rect 99372 4508 99540 4510
rect 99484 4498 99540 4508
rect 99596 4116 99652 5742
rect 100380 5012 100436 5022
rect 99820 4898 99876 4910
rect 99820 4846 99822 4898
rect 99874 4846 99876 4898
rect 99820 4340 99876 4846
rect 100380 4450 100436 4956
rect 100380 4398 100382 4450
rect 100434 4398 100436 4450
rect 100380 4386 100436 4398
rect 100604 5012 100660 5022
rect 100604 4340 100660 4956
rect 99820 4274 99876 4284
rect 100492 4338 100660 4340
rect 100492 4286 100606 4338
rect 100658 4286 100660 4338
rect 100492 4284 100660 4286
rect 100492 4228 100548 4284
rect 100604 4274 100660 4284
rect 100716 4452 100772 4462
rect 99596 4050 99652 4060
rect 99932 4116 99988 4126
rect 99932 3442 99988 4060
rect 99932 3390 99934 3442
rect 99986 3390 99988 3442
rect 99932 3378 99988 3390
rect 100492 3442 100548 4172
rect 100716 3778 100772 4396
rect 100716 3726 100718 3778
rect 100770 3726 100772 3778
rect 100716 3714 100772 3726
rect 100940 3780 100996 12012
rect 101164 12002 101220 12012
rect 101500 8428 101556 12798
rect 101836 12850 101892 15372
rect 101836 12798 101838 12850
rect 101890 12798 101892 12850
rect 101836 12786 101892 12798
rect 105532 14308 105588 14318
rect 102844 12068 102900 12078
rect 102844 10164 102900 12012
rect 102844 10098 102900 10108
rect 101388 8372 101556 8428
rect 101164 4898 101220 4910
rect 101164 4846 101166 4898
rect 101218 4846 101220 4898
rect 101052 4340 101108 4350
rect 101052 4246 101108 4284
rect 101052 3780 101108 3790
rect 100940 3778 101108 3780
rect 100940 3726 101054 3778
rect 101106 3726 101108 3778
rect 100940 3724 101108 3726
rect 101052 3714 101108 3724
rect 100492 3390 100494 3442
rect 100546 3390 100548 3442
rect 100492 3378 100548 3390
rect 101164 980 101220 4846
rect 101388 4562 101444 8372
rect 103516 6468 103572 6478
rect 103516 6466 104132 6468
rect 103516 6414 103518 6466
rect 103570 6414 104132 6466
rect 103516 6412 104132 6414
rect 103516 6402 103572 6412
rect 103068 5908 103124 5918
rect 102508 5794 102564 5806
rect 102956 5796 103012 5806
rect 102508 5742 102510 5794
rect 102562 5742 102564 5794
rect 102060 5012 102116 5022
rect 102060 4918 102116 4956
rect 101388 4510 101390 4562
rect 101442 4510 101444 4562
rect 101388 4498 101444 4510
rect 101612 4898 101668 4910
rect 101612 4846 101614 4898
rect 101666 4846 101668 4898
rect 101612 4452 101668 4846
rect 102508 4564 102564 5742
rect 102844 5794 103012 5796
rect 102844 5742 102958 5794
rect 103010 5742 103012 5794
rect 102844 5740 103012 5742
rect 102620 5124 102676 5134
rect 102620 5030 102676 5068
rect 102844 5012 102900 5740
rect 102956 5730 103012 5740
rect 103068 5234 103124 5852
rect 103964 5908 104020 5918
rect 103964 5814 104020 5852
rect 103068 5182 103070 5234
rect 103122 5182 103124 5234
rect 103068 5124 103124 5182
rect 103068 5058 103124 5068
rect 103516 5794 103572 5806
rect 103516 5742 103518 5794
rect 103570 5742 103572 5794
rect 102508 4508 102676 4564
rect 102172 4452 102228 4462
rect 101612 4450 102228 4452
rect 101612 4398 102174 4450
rect 102226 4398 102228 4450
rect 101612 4396 102228 4398
rect 101612 1652 101668 4396
rect 102172 4386 102228 4396
rect 102060 4116 102116 4126
rect 101612 1586 101668 1596
rect 101724 3442 101780 3454
rect 101724 3390 101726 3442
rect 101778 3390 101780 3442
rect 100940 924 101332 980
rect 100940 800 100996 924
rect 5152 0 5264 800
rect 6832 0 6944 800
rect 8512 0 8624 800
rect 10192 0 10304 800
rect 11872 0 11984 800
rect 13552 0 13664 800
rect 15232 0 15344 800
rect 16912 0 17024 800
rect 18592 0 18704 800
rect 20272 0 20384 800
rect 21952 0 22064 800
rect 23632 0 23744 800
rect 25312 0 25424 800
rect 26992 0 27104 800
rect 28672 0 28784 800
rect 30352 0 30464 800
rect 32032 0 32144 800
rect 33712 0 33824 800
rect 35392 0 35504 800
rect 37072 0 37184 800
rect 38752 0 38864 800
rect 40432 0 40544 800
rect 42112 0 42224 800
rect 43792 0 43904 800
rect 45472 0 45584 800
rect 47152 0 47264 800
rect 48832 0 48944 800
rect 50512 0 50624 800
rect 52192 0 52304 800
rect 53872 0 53984 800
rect 55552 0 55664 800
rect 57232 0 57344 800
rect 58912 0 59024 800
rect 60592 0 60704 800
rect 62272 0 62384 800
rect 63952 0 64064 800
rect 65632 0 65744 800
rect 67312 0 67424 800
rect 68992 0 69104 800
rect 70672 0 70784 800
rect 72352 0 72464 800
rect 74032 0 74144 800
rect 75712 0 75824 800
rect 77392 0 77504 800
rect 79072 0 79184 800
rect 80752 0 80864 800
rect 82432 0 82544 800
rect 84112 0 84224 800
rect 85792 0 85904 800
rect 87472 0 87584 800
rect 89152 0 89264 800
rect 90832 0 90944 800
rect 92512 0 92624 800
rect 94192 0 94304 800
rect 95872 0 95984 800
rect 97552 0 97664 800
rect 99232 0 99344 800
rect 100912 0 101024 800
rect 101276 756 101332 924
rect 101724 756 101780 3390
rect 102060 3330 102116 4060
rect 102060 3278 102062 3330
rect 102114 3278 102116 3330
rect 102060 3266 102116 3278
rect 102620 3442 102676 4508
rect 102732 4450 102788 4462
rect 102732 4398 102734 4450
rect 102786 4398 102788 4450
rect 102732 4340 102788 4398
rect 102732 4274 102788 4284
rect 102620 3390 102622 3442
rect 102674 3390 102676 3442
rect 102620 800 102676 3390
rect 102844 2436 102900 4956
rect 103516 4564 103572 5742
rect 103740 5012 103796 5022
rect 103740 4918 103796 4956
rect 103516 4498 103572 4508
rect 103292 4340 103348 4350
rect 103964 4340 104020 4350
rect 103292 4338 104020 4340
rect 103292 4286 103294 4338
rect 103346 4286 103966 4338
rect 104018 4286 104020 4338
rect 103292 4284 104020 4286
rect 103292 4274 103348 4284
rect 103964 4274 104020 4284
rect 102956 4116 103012 4126
rect 102956 4022 103012 4060
rect 104076 3668 104132 6412
rect 105532 6130 105588 14252
rect 105868 10164 105924 10174
rect 105532 6078 105534 6130
rect 105586 6078 105588 6130
rect 105532 6066 105588 6078
rect 105644 6580 105700 6590
rect 104412 5908 104468 5918
rect 105196 5908 105252 5918
rect 104412 5814 104468 5852
rect 104860 5906 105252 5908
rect 104860 5854 105198 5906
rect 105250 5854 105252 5906
rect 104860 5852 105252 5854
rect 104860 5346 104916 5852
rect 105196 5842 105252 5852
rect 104860 5294 104862 5346
rect 104914 5294 104916 5346
rect 104860 5282 104916 5294
rect 104300 5124 104356 5134
rect 102956 3556 103012 3566
rect 102956 3330 103012 3500
rect 104076 3442 104132 3612
rect 104188 5010 104244 5022
rect 104188 4958 104190 5010
rect 104242 4958 104244 5010
rect 104188 4340 104244 4958
rect 104300 4562 104356 5068
rect 104300 4510 104302 4562
rect 104354 4510 104356 4562
rect 104300 4498 104356 4510
rect 104524 5122 104580 5134
rect 104524 5070 104526 5122
rect 104578 5070 104580 5122
rect 104188 3554 104244 4284
rect 104188 3502 104190 3554
rect 104242 3502 104244 3554
rect 104188 3490 104244 3502
rect 104076 3390 104078 3442
rect 104130 3390 104132 3442
rect 104076 3378 104132 3390
rect 104412 3444 104468 3454
rect 102956 3278 102958 3330
rect 103010 3278 103012 3330
rect 102956 3266 103012 3278
rect 104412 2884 104468 3388
rect 104524 2994 104580 5070
rect 105532 5012 105588 5022
rect 104972 5010 105588 5012
rect 104972 4958 105534 5010
rect 105586 4958 105588 5010
rect 104972 4956 105588 4958
rect 104972 3778 105028 4956
rect 105532 4946 105588 4956
rect 105644 4564 105700 6524
rect 105868 5010 105924 10108
rect 105868 4958 105870 5010
rect 105922 4958 105924 5010
rect 105868 4946 105924 4958
rect 106428 5010 106484 5022
rect 106428 4958 106430 5010
rect 106482 4958 106484 5010
rect 105532 4452 105588 4462
rect 105644 4452 105700 4508
rect 106428 4562 106484 4958
rect 106764 5010 106820 18284
rect 108332 15876 108388 15886
rect 108332 5124 108388 15820
rect 109564 10388 109620 10398
rect 108332 5058 108388 5068
rect 109004 7588 109060 7598
rect 106764 4958 106766 5010
rect 106818 4958 106820 5010
rect 106764 4946 106820 4958
rect 106428 4510 106430 4562
rect 106482 4510 106484 4562
rect 106428 4498 106484 4510
rect 106988 4564 107044 4574
rect 106988 4470 107044 4508
rect 109004 4562 109060 7532
rect 109564 5236 109620 10332
rect 110236 5794 110292 5806
rect 110236 5742 110238 5794
rect 110290 5742 110292 5794
rect 110236 5236 110292 5742
rect 109564 5104 109620 5180
rect 109900 5180 110292 5236
rect 109004 4510 109006 4562
rect 109058 4510 109060 4562
rect 105532 4450 105700 4452
rect 105532 4398 105534 4450
rect 105586 4398 105700 4450
rect 105532 4396 105700 4398
rect 105532 4386 105588 4396
rect 105308 4340 105364 4350
rect 105308 4246 105364 4284
rect 107436 4226 107492 4238
rect 107436 4174 107438 4226
rect 107490 4174 107492 4226
rect 106092 4116 106148 4126
rect 106092 4114 106596 4116
rect 106092 4062 106094 4114
rect 106146 4062 106596 4114
rect 106092 4060 106596 4062
rect 106092 4050 106148 4060
rect 104972 3726 104974 3778
rect 105026 3726 105028 3778
rect 104972 3714 105028 3726
rect 104636 3556 104692 3566
rect 104636 3462 104692 3500
rect 106092 3556 106148 3566
rect 105980 3444 106036 3454
rect 105980 3350 106036 3388
rect 104524 2942 104526 2994
rect 104578 2942 104580 2994
rect 104524 2930 104580 2942
rect 105644 3330 105700 3342
rect 105644 3278 105646 3330
rect 105698 3278 105700 3330
rect 105644 2994 105700 3278
rect 105644 2942 105646 2994
rect 105698 2942 105700 2994
rect 105644 2930 105700 2942
rect 102844 2370 102900 2380
rect 104300 2828 104468 2884
rect 104300 800 104356 2828
rect 106092 2660 106148 3500
rect 106540 3442 106596 4060
rect 106764 3556 106820 3566
rect 106764 3462 106820 3500
rect 106540 3390 106542 3442
rect 106594 3390 106596 3442
rect 106540 3378 106596 3390
rect 107436 3444 107492 4174
rect 107884 4226 107940 4238
rect 107884 4174 107886 4226
rect 107938 4174 107940 4226
rect 107884 3668 107940 4174
rect 108556 4228 108612 4238
rect 108556 4134 108612 4172
rect 107884 3602 107940 3612
rect 108220 3556 108276 3566
rect 107884 3444 107940 3454
rect 107436 3378 107492 3388
rect 107660 3388 107884 3444
rect 105980 2604 106148 2660
rect 105980 800 106036 2604
rect 107660 800 107716 3388
rect 107884 3312 107940 3388
rect 108220 3330 108276 3500
rect 108668 3444 108724 3454
rect 108668 3350 108724 3388
rect 109004 3444 109060 4510
rect 109900 4676 109956 5180
rect 110012 5012 110068 5022
rect 110012 5010 110292 5012
rect 110012 4958 110014 5010
rect 110066 4958 110292 5010
rect 110012 4956 110292 4958
rect 110012 4946 110068 4956
rect 109788 4452 109844 4462
rect 109788 4358 109844 4396
rect 109452 4340 109508 4350
rect 109004 3378 109060 3388
rect 109340 4338 109508 4340
rect 109340 4286 109454 4338
rect 109506 4286 109508 4338
rect 109340 4284 109508 4286
rect 109340 4228 109396 4284
rect 109452 4274 109508 4284
rect 108220 3278 108222 3330
rect 108274 3278 108276 3330
rect 108220 3266 108276 3278
rect 109340 800 109396 4172
rect 109900 3668 109956 4620
rect 109900 3602 109956 3612
rect 110012 4340 110068 4350
rect 109452 3444 109508 3454
rect 109452 3350 109508 3388
rect 110012 3442 110068 4284
rect 110236 4116 110292 4956
rect 110348 5010 110404 19180
rect 111672 18844 111936 18854
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111672 18778 111936 18788
rect 114044 18674 114100 20748
rect 114044 18622 114046 18674
rect 114098 18622 114100 18674
rect 114044 18610 114100 18622
rect 113708 18450 113764 18462
rect 113708 18398 113710 18450
rect 113762 18398 113764 18450
rect 113148 18340 113204 18350
rect 113708 18340 113764 18398
rect 113148 18338 113764 18340
rect 113148 18286 113150 18338
rect 113202 18286 113764 18338
rect 113148 18284 113764 18286
rect 111672 17276 111936 17286
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111672 17210 111936 17220
rect 111672 15708 111936 15718
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111672 15642 111936 15652
rect 111672 14140 111936 14150
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111672 14074 111936 14084
rect 111672 12572 111936 12582
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111672 12506 111936 12516
rect 111672 11004 111936 11014
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111672 10938 111936 10948
rect 111672 9436 111936 9446
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111672 9370 111936 9380
rect 112140 9268 112196 9278
rect 110348 4958 110350 5010
rect 110402 4958 110404 5010
rect 110348 4946 110404 4958
rect 110572 9044 110628 9054
rect 110572 4564 110628 8988
rect 111672 7868 111936 7878
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111672 7802 111936 7812
rect 111580 6468 111636 6478
rect 111468 6466 111636 6468
rect 111468 6414 111582 6466
rect 111634 6414 111636 6466
rect 111468 6412 111636 6414
rect 111244 5908 111300 5918
rect 111244 5814 111300 5852
rect 111468 5908 111524 6412
rect 111580 6402 111636 6412
rect 111672 6300 111936 6310
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111672 6234 111936 6244
rect 112140 6130 112196 9212
rect 113148 8428 113204 18284
rect 112140 6078 112142 6130
rect 112194 6078 112196 6130
rect 112140 6066 112196 6078
rect 112700 8372 113204 8428
rect 111468 5842 111524 5852
rect 111916 5908 111972 5918
rect 111916 5906 112084 5908
rect 111916 5854 111918 5906
rect 111970 5854 112084 5906
rect 111916 5852 112084 5854
rect 111916 5842 111972 5852
rect 110572 4450 110628 4508
rect 110572 4398 110574 4450
rect 110626 4398 110628 4450
rect 110572 4386 110628 4398
rect 110796 5794 110852 5806
rect 110796 5742 110798 5794
rect 110850 5742 110852 5794
rect 110460 4340 110516 4350
rect 110460 4246 110516 4284
rect 110796 4340 110852 5742
rect 111020 5236 111076 5246
rect 111020 5010 111076 5180
rect 111804 5124 111860 5134
rect 111804 5030 111860 5068
rect 111020 4958 111022 5010
rect 111074 4958 111076 5010
rect 111020 4946 111076 4958
rect 111468 5010 111524 5022
rect 111468 4958 111470 5010
rect 111522 4958 111524 5010
rect 110796 4274 110852 4284
rect 111468 4340 111524 4958
rect 111672 4732 111936 4742
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111672 4666 111936 4676
rect 111580 4564 111636 4574
rect 112028 4564 112084 5852
rect 112252 5124 112308 5134
rect 112140 5012 112196 5022
rect 112140 4918 112196 4956
rect 111580 4562 112084 4564
rect 111580 4510 111582 4562
rect 111634 4510 112084 4562
rect 111580 4508 112084 4510
rect 112140 4564 112196 4574
rect 111580 4498 111636 4508
rect 112140 4470 112196 4508
rect 111468 4274 111524 4284
rect 111804 4340 111860 4350
rect 110236 4060 110628 4116
rect 110572 3778 110628 4060
rect 110572 3726 110574 3778
rect 110626 3726 110628 3778
rect 110572 3714 110628 3726
rect 111244 4114 111300 4126
rect 111244 4062 111246 4114
rect 111298 4062 111300 4114
rect 110236 3556 110292 3566
rect 110236 3462 110292 3500
rect 110012 3390 110014 3442
rect 110066 3390 110068 3442
rect 110012 3378 110068 3390
rect 111020 3444 111076 3454
rect 111020 800 111076 3388
rect 111244 3332 111300 4062
rect 111692 3668 111748 3678
rect 111692 3442 111748 3612
rect 111804 3554 111860 4284
rect 112252 3892 112308 5068
rect 112252 3826 112308 3836
rect 112476 4452 112532 4462
rect 112476 3778 112532 4396
rect 112476 3726 112478 3778
rect 112530 3726 112532 3778
rect 112476 3714 112532 3726
rect 112700 3780 112756 8372
rect 113484 7812 113540 7822
rect 113484 7698 113540 7756
rect 113484 7646 113486 7698
rect 113538 7646 113540 7698
rect 113484 7634 113540 7646
rect 113148 7474 113204 7486
rect 113148 7422 113150 7474
rect 113202 7422 113204 7474
rect 113148 5572 113204 7422
rect 114268 6804 114324 6814
rect 113260 5796 113316 5806
rect 113260 5794 113428 5796
rect 113260 5742 113262 5794
rect 113314 5742 113428 5794
rect 113260 5740 113428 5742
rect 113260 5730 113316 5740
rect 113148 5516 113316 5572
rect 112812 5012 112868 5022
rect 112812 4918 112868 4956
rect 113148 5012 113204 5022
rect 113148 4918 113204 4956
rect 113260 4562 113316 5516
rect 113260 4510 113262 4562
rect 113314 4510 113316 4562
rect 113260 4498 113316 4510
rect 112812 3780 112868 3790
rect 112700 3778 112868 3780
rect 112700 3726 112814 3778
rect 112866 3726 112868 3778
rect 112700 3724 112868 3726
rect 112812 3714 112868 3724
rect 111804 3502 111806 3554
rect 111858 3502 111860 3554
rect 111804 3490 111860 3502
rect 112812 3556 112868 3566
rect 111692 3390 111694 3442
rect 111746 3390 111748 3442
rect 111692 3378 111748 3390
rect 111244 3266 111300 3276
rect 111672 3164 111936 3174
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111672 3098 111936 3108
rect 112476 2548 112532 2558
rect 112476 1540 112532 2492
rect 112476 1474 112532 1484
rect 112812 1204 112868 3500
rect 113372 3444 113428 5740
rect 114156 5794 114212 5806
rect 114156 5742 114158 5794
rect 114210 5742 114212 5794
rect 114156 5684 114212 5742
rect 113932 5628 114212 5684
rect 113372 3378 113428 3388
rect 113596 4898 113652 4910
rect 113596 4846 113598 4898
rect 113650 4846 113652 4898
rect 113596 4114 113652 4846
rect 113596 4062 113598 4114
rect 113650 4062 113652 4114
rect 113484 3332 113540 3342
rect 113484 3238 113540 3276
rect 113596 2324 113652 4062
rect 113820 3444 113876 3454
rect 113820 3350 113876 3388
rect 113596 2258 113652 2268
rect 113932 3332 113988 5628
rect 114044 5236 114100 5246
rect 114044 4338 114100 5180
rect 114044 4286 114046 4338
rect 114098 4286 114100 4338
rect 114044 4274 114100 4286
rect 114156 4900 114212 4910
rect 114044 3892 114100 3902
rect 114044 3444 114100 3836
rect 114156 3444 114212 4844
rect 114268 4564 114324 6748
rect 114604 5010 114660 5022
rect 114604 4958 114606 5010
rect 114658 4958 114660 5010
rect 114604 4900 114660 4958
rect 115164 5012 115220 22316
rect 118412 21476 118468 21486
rect 116620 16996 116676 17006
rect 115948 11396 116004 11406
rect 115948 7812 116004 11340
rect 116620 10164 116676 16940
rect 116620 10098 116676 10108
rect 118412 9268 118468 21420
rect 119420 19348 119476 19358
rect 119196 17444 119252 17454
rect 119196 14308 119252 17388
rect 119196 14242 119252 14252
rect 118412 9202 118468 9212
rect 115948 7746 116004 7756
rect 118524 6804 118580 6814
rect 117852 5908 117908 5918
rect 115612 5796 115668 5806
rect 116060 5796 116116 5806
rect 117068 5796 117124 5806
rect 115612 5794 115892 5796
rect 115612 5742 115614 5794
rect 115666 5742 115892 5794
rect 115612 5740 115892 5742
rect 115612 5730 115668 5740
rect 115388 5236 115444 5246
rect 115388 5142 115444 5180
rect 115164 4946 115220 4956
rect 115612 5012 115668 5022
rect 114604 4834 114660 4844
rect 114940 4900 114996 4910
rect 114940 4898 115108 4900
rect 114940 4846 114942 4898
rect 114994 4846 115108 4898
rect 114940 4844 115108 4846
rect 114940 4834 114996 4844
rect 114940 4564 114996 4574
rect 114268 4562 114996 4564
rect 114268 4510 114942 4562
rect 114994 4510 114996 4562
rect 114268 4508 114996 4510
rect 114268 4450 114324 4508
rect 114940 4498 114996 4508
rect 114268 4398 114270 4450
rect 114322 4398 114324 4450
rect 114268 4386 114324 4398
rect 115052 3892 115108 4844
rect 115052 3826 115108 3836
rect 115612 3778 115668 4956
rect 115612 3726 115614 3778
rect 115666 3726 115668 3778
rect 115612 3714 115668 3726
rect 115836 4452 115892 5740
rect 116060 5794 116228 5796
rect 116060 5742 116062 5794
rect 116114 5742 116228 5794
rect 116060 5740 116228 5742
rect 116060 5730 116116 5740
rect 115948 5012 116004 5022
rect 115948 4918 116004 4956
rect 115948 4452 116004 4462
rect 115836 4450 116004 4452
rect 115836 4398 115950 4450
rect 116002 4398 116004 4450
rect 115836 4396 116004 4398
rect 114604 3556 114660 3566
rect 115836 3556 115892 4396
rect 115948 4386 116004 4396
rect 115948 3892 116004 3902
rect 115948 3778 116004 3836
rect 115948 3726 115950 3778
rect 116002 3726 116004 3778
rect 115948 3714 116004 3726
rect 116172 3668 116228 5740
rect 117068 5794 117236 5796
rect 117068 5742 117070 5794
rect 117122 5742 117236 5794
rect 117068 5740 117236 5742
rect 117068 5730 117124 5740
rect 116284 5012 116340 5022
rect 117068 5012 117124 5022
rect 116284 4918 116340 4956
rect 116956 5010 117124 5012
rect 116956 4958 117070 5010
rect 117122 4958 117124 5010
rect 116956 4956 117124 4958
rect 116508 4452 116564 4462
rect 116956 4452 117012 4956
rect 117068 4946 117124 4956
rect 117068 4564 117124 4574
rect 117068 4470 117124 4508
rect 116508 4450 117012 4452
rect 116508 4398 116510 4450
rect 116562 4398 117012 4450
rect 116508 4396 117012 4398
rect 116508 4386 116564 4396
rect 116172 3602 116228 3612
rect 116508 3668 116564 3678
rect 115836 3500 116004 3556
rect 114604 3462 114660 3500
rect 114380 3444 114436 3454
rect 114156 3388 114324 3444
rect 114044 3378 114100 3388
rect 112812 1138 112868 1148
rect 112700 924 113092 980
rect 112700 800 112756 924
rect 101276 700 101780 756
rect 102592 0 102704 800
rect 104272 0 104384 800
rect 105952 0 106064 800
rect 107632 0 107744 800
rect 109312 0 109424 800
rect 110992 0 111104 800
rect 112672 0 112784 800
rect 113036 756 113092 924
rect 113932 756 113988 3276
rect 114268 1540 114324 3388
rect 114380 3330 114436 3388
rect 114380 3278 114382 3330
rect 114434 3278 114436 3330
rect 114380 3266 114436 3278
rect 114268 1484 114436 1540
rect 114380 800 114436 1484
rect 115948 1316 116004 3500
rect 115948 1250 116004 1260
rect 116060 3444 116116 3454
rect 116060 800 116116 3388
rect 116508 3442 116564 3612
rect 116620 3556 116676 4396
rect 116732 4116 116788 4126
rect 116732 4114 117124 4116
rect 116732 4062 116734 4114
rect 116786 4062 117124 4114
rect 116732 4060 117124 4062
rect 116732 4050 116788 4060
rect 116732 3556 116788 3566
rect 116620 3500 116732 3556
rect 116732 3462 116788 3500
rect 116508 3390 116510 3442
rect 116562 3390 116564 3442
rect 116508 3378 116564 3390
rect 117068 3220 117124 4060
rect 117180 3444 117236 5740
rect 117516 5794 117572 5806
rect 117516 5742 117518 5794
rect 117570 5742 117572 5794
rect 117516 4452 117572 5742
rect 117852 5794 117908 5852
rect 117852 5742 117854 5794
rect 117906 5742 117908 5794
rect 117628 5124 117684 5134
rect 117628 5030 117684 5068
rect 117852 5124 117908 5742
rect 117852 5058 117908 5068
rect 118300 5794 118356 5806
rect 118300 5742 118302 5794
rect 118354 5742 118356 5794
rect 118188 5010 118244 5022
rect 118188 4958 118190 5010
rect 118242 4958 118244 5010
rect 118188 4564 118244 4958
rect 118188 4498 118244 4508
rect 117852 4452 117908 4462
rect 117516 4450 117908 4452
rect 117516 4398 117854 4450
rect 117906 4398 117908 4450
rect 117516 4396 117908 4398
rect 117180 3378 117236 3388
rect 117740 3444 117796 3454
rect 117740 3350 117796 3388
rect 117404 3330 117460 3342
rect 117404 3278 117406 3330
rect 117458 3278 117460 3330
rect 117404 3220 117460 3278
rect 117068 3164 117460 3220
rect 117852 1204 117908 4396
rect 118300 3442 118356 5742
rect 118524 5010 118580 6748
rect 119196 5794 119252 5806
rect 119196 5742 119198 5794
rect 119250 5742 119252 5794
rect 118524 4958 118526 5010
rect 118578 4958 118580 5010
rect 118524 4946 118580 4958
rect 119084 5010 119140 5022
rect 119084 4958 119086 5010
rect 119138 4958 119140 5010
rect 118972 4564 119028 4574
rect 119084 4564 119140 4958
rect 118972 4562 119140 4564
rect 118972 4510 118974 4562
rect 119026 4510 119140 4562
rect 118972 4508 119140 4510
rect 118972 4498 119028 4508
rect 118412 4450 118468 4462
rect 118412 4398 118414 4450
rect 118466 4398 118468 4450
rect 118412 3556 118468 4398
rect 118412 3490 118468 3500
rect 118636 4114 118692 4126
rect 118636 4062 118638 4114
rect 118690 4062 118692 4114
rect 118300 3390 118302 3442
rect 118354 3390 118356 3442
rect 118300 3388 118356 3390
rect 117852 1138 117908 1148
rect 117964 3332 118356 3388
rect 118636 3442 118692 4062
rect 118636 3390 118638 3442
rect 118690 3390 118692 3442
rect 118636 3378 118692 3390
rect 119196 3444 119252 5742
rect 119420 5010 119476 19292
rect 120316 11732 120372 11742
rect 119420 4958 119422 5010
rect 119474 4958 119476 5010
rect 119420 4946 119476 4958
rect 119980 5012 120036 5022
rect 119980 5010 120260 5012
rect 119980 4958 119982 5010
rect 120034 4958 120260 5010
rect 119980 4956 120260 4958
rect 119980 4946 120036 4956
rect 120204 4564 120260 4956
rect 120316 5010 120372 11676
rect 120316 4958 120318 5010
rect 120370 4958 120372 5010
rect 120316 4946 120372 4958
rect 121436 7700 121492 7710
rect 121100 4898 121156 4910
rect 121100 4846 121102 4898
rect 121154 4846 121156 4898
rect 120204 4508 120708 4564
rect 119980 4452 120036 4462
rect 119980 4450 120372 4452
rect 119980 4398 119982 4450
rect 120034 4398 120372 4450
rect 119980 4396 120372 4398
rect 119980 4386 120036 4396
rect 119644 4340 119700 4350
rect 119196 3378 119252 3388
rect 119420 4284 119644 4340
rect 117964 980 118020 3332
rect 117740 924 118020 980
rect 117740 800 117796 924
rect 119420 800 119476 4284
rect 119644 4208 119700 4284
rect 120316 3778 120372 4396
rect 120316 3726 120318 3778
rect 120370 3726 120372 3778
rect 120316 3714 120372 3726
rect 120652 3778 120708 4508
rect 120988 4340 121044 4350
rect 120988 4246 121044 4284
rect 120652 3726 120654 3778
rect 120706 3726 120708 3778
rect 120652 3714 120708 3726
rect 120988 3668 121044 3678
rect 119644 3556 119700 3566
rect 119644 3462 119700 3500
rect 119532 3444 119588 3454
rect 119532 1428 119588 3388
rect 120988 2660 121044 3612
rect 120988 2594 121044 2604
rect 121100 3444 121156 4846
rect 121436 4562 121492 7644
rect 121884 5012 121940 23100
rect 123452 11732 123508 25228
rect 123452 11666 123508 11676
rect 125132 23716 125188 23726
rect 124012 10948 124068 10958
rect 123676 8484 123732 8494
rect 121884 4946 121940 4956
rect 122780 5122 122836 5134
rect 122780 5070 122782 5122
rect 122834 5070 122836 5122
rect 121436 4510 121438 4562
rect 121490 4510 121492 4562
rect 121436 4452 121492 4510
rect 122108 4452 122164 4462
rect 121436 4450 122164 4452
rect 121436 4398 122110 4450
rect 122162 4398 122164 4450
rect 121436 4396 122164 4398
rect 122108 4386 122164 4396
rect 122668 4452 122724 4462
rect 122668 4358 122724 4396
rect 121660 4116 121716 4126
rect 121324 3444 121380 3454
rect 121100 3442 121380 3444
rect 121100 3390 121326 3442
rect 121378 3390 121380 3442
rect 121100 3388 121380 3390
rect 119532 1362 119588 1372
rect 121100 800 121156 3388
rect 121324 3378 121380 3388
rect 121660 3330 121716 4060
rect 122556 3556 122612 3566
rect 122220 3444 122276 3454
rect 122220 3350 122276 3388
rect 121660 3278 121662 3330
rect 121714 3278 121716 3330
rect 121660 3266 121716 3278
rect 122556 3330 122612 3500
rect 122556 3278 122558 3330
rect 122610 3278 122612 3330
rect 122556 3266 122612 3278
rect 122780 3444 122836 5070
rect 123564 5012 123620 5022
rect 123228 5010 123620 5012
rect 123228 4958 123566 5010
rect 123618 4958 123620 5010
rect 123228 4956 123620 4958
rect 123228 4562 123284 4956
rect 123564 4946 123620 4956
rect 123228 4510 123230 4562
rect 123282 4510 123284 4562
rect 123228 4498 123284 4510
rect 122892 4116 122948 4126
rect 122892 4022 122948 4060
rect 122780 800 122836 3388
rect 123676 3892 123732 8428
rect 123900 5796 123956 5806
rect 123900 5702 123956 5740
rect 123900 5012 123956 5022
rect 124012 5012 124068 10892
rect 125132 6804 125188 23660
rect 125132 6738 125188 6748
rect 125356 7588 125412 7598
rect 123900 5010 124068 5012
rect 123900 4958 123902 5010
rect 123954 4958 124068 5010
rect 123900 4956 124068 4958
rect 124348 5796 124404 5806
rect 123900 4946 123956 4956
rect 123676 3442 123732 3836
rect 123676 3390 123678 3442
rect 123730 3390 123732 3442
rect 123676 3378 123732 3390
rect 124012 4452 124068 4462
rect 124012 3442 124068 4396
rect 124348 4450 124404 5740
rect 125020 5012 125076 5022
rect 124348 4398 124350 4450
rect 124402 4398 124404 4450
rect 124236 3556 124292 3566
rect 124236 3462 124292 3500
rect 124012 3390 124014 3442
rect 124066 3390 124068 3442
rect 124012 3378 124068 3390
rect 124348 1204 124404 4398
rect 124572 5010 125076 5012
rect 124572 4958 125022 5010
rect 125074 4958 125076 5010
rect 124572 4956 125076 4958
rect 124572 3778 124628 4956
rect 125020 4946 125076 4956
rect 125356 5010 125412 7532
rect 125916 5348 125972 5358
rect 125916 5236 125972 5292
rect 125916 5180 126084 5236
rect 125916 5012 125972 5022
rect 125356 4958 125358 5010
rect 125410 4958 125412 5010
rect 125356 4946 125412 4958
rect 125468 5010 125972 5012
rect 125468 4958 125918 5010
rect 125970 4958 125972 5010
rect 125468 4956 125972 4958
rect 125356 4564 125412 4574
rect 125468 4564 125524 4956
rect 125916 4946 125972 4956
rect 125356 4562 125524 4564
rect 125356 4510 125358 4562
rect 125410 4510 125524 4562
rect 125356 4508 125524 4510
rect 125356 4498 125412 4508
rect 124796 4452 124852 4462
rect 126028 4452 126084 5180
rect 126252 5010 126308 27692
rect 127708 10500 127764 10510
rect 127596 8148 127652 8158
rect 127596 5794 127652 8092
rect 127708 6580 127764 10444
rect 128268 8428 128324 29372
rect 130082 29036 130346 29046
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130082 28970 130346 28980
rect 130082 27468 130346 27478
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130082 27402 130346 27412
rect 130082 25900 130346 25910
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130082 25834 130346 25844
rect 130082 24332 130346 24342
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130082 24266 130346 24276
rect 130082 22764 130346 22774
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130082 22698 130346 22708
rect 130082 21196 130346 21206
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130082 21130 130346 21140
rect 130082 19628 130346 19638
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130082 19562 130346 19572
rect 130082 18060 130346 18070
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130082 17994 130346 18004
rect 130082 16492 130346 16502
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130082 16426 130346 16436
rect 130082 14924 130346 14934
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130082 14858 130346 14868
rect 130082 13356 130346 13366
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130082 13290 130346 13300
rect 130082 11788 130346 11798
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130082 11722 130346 11732
rect 130082 10220 130346 10230
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130082 10154 130346 10164
rect 130082 8652 130346 8662
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130082 8586 130346 8596
rect 127708 6514 127764 6524
rect 128156 8372 128324 8428
rect 127596 5742 127598 5794
rect 127650 5742 127652 5794
rect 127036 5124 127092 5134
rect 126252 4958 126254 5010
rect 126306 4958 126308 5010
rect 126252 4946 126308 4958
rect 126700 5012 126756 5022
rect 126364 4452 126420 4462
rect 126028 4450 126420 4452
rect 126028 4398 126366 4450
rect 126418 4398 126420 4450
rect 126028 4396 126420 4398
rect 124796 4358 124852 4396
rect 125020 4116 125076 4126
rect 125020 4114 125300 4116
rect 125020 4062 125022 4114
rect 125074 4062 125300 4114
rect 125020 4060 125300 4062
rect 125020 4050 125076 4060
rect 124572 3726 124574 3778
rect 124626 3726 124628 3778
rect 124572 3714 124628 3726
rect 124348 1138 124404 1148
rect 124460 3444 124516 3454
rect 124460 800 124516 3388
rect 125244 3442 125300 4060
rect 126028 3892 126084 3902
rect 126028 3666 126084 3836
rect 126028 3614 126030 3666
rect 126082 3614 126084 3666
rect 126028 3602 126084 3614
rect 126364 3668 126420 4396
rect 126700 4452 126756 4956
rect 127036 5010 127092 5068
rect 127372 5124 127428 5134
rect 127596 5124 127652 5742
rect 127372 5122 127652 5124
rect 127372 5070 127374 5122
rect 127426 5070 127652 5122
rect 127372 5068 127652 5070
rect 127372 5058 127428 5068
rect 127036 4958 127038 5010
rect 127090 4958 127092 5010
rect 127036 4946 127092 4958
rect 127932 5010 127988 5022
rect 127932 4958 127934 5010
rect 127986 4958 127988 5010
rect 127260 4564 127316 4574
rect 127260 4470 127316 4508
rect 127932 4564 127988 4958
rect 128156 5012 128212 8372
rect 130082 7084 130346 7094
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130082 7018 130346 7028
rect 129276 6580 129332 6590
rect 129276 6486 129332 6524
rect 129836 6580 129892 6590
rect 128604 6466 128660 6478
rect 128604 6414 128606 6466
rect 128658 6414 128660 6466
rect 128268 5796 128324 5806
rect 128268 5794 128436 5796
rect 128268 5742 128270 5794
rect 128322 5742 128436 5794
rect 128268 5740 128436 5742
rect 128268 5730 128324 5740
rect 128268 5012 128324 5022
rect 128156 5010 128324 5012
rect 128156 4958 128270 5010
rect 128322 4958 128324 5010
rect 128156 4956 128324 4958
rect 128268 4946 128324 4956
rect 128380 4788 128436 5740
rect 127932 4498 127988 4508
rect 128156 4732 128436 4788
rect 126700 4320 126756 4396
rect 127932 4340 127988 4350
rect 128156 4340 128212 4732
rect 127820 4338 128212 4340
rect 127820 4286 127934 4338
rect 127986 4286 128212 4338
rect 127820 4284 128212 4286
rect 128268 4450 128324 4462
rect 128268 4398 128270 4450
rect 128322 4398 128324 4450
rect 126924 4116 126980 4126
rect 126924 4114 127204 4116
rect 126924 4062 126926 4114
rect 126978 4062 127204 4114
rect 126924 4060 127204 4062
rect 126924 4050 126980 4060
rect 126588 3668 126644 3678
rect 126364 3666 126644 3668
rect 126364 3614 126590 3666
rect 126642 3614 126644 3666
rect 126364 3612 126644 3614
rect 126588 3602 126644 3612
rect 126140 3556 126196 3566
rect 125244 3390 125246 3442
rect 125298 3390 125300 3442
rect 125244 3378 125300 3390
rect 125580 3444 125636 3454
rect 125580 3350 125636 3388
rect 126140 800 126196 3500
rect 127148 3444 127204 4060
rect 127484 3556 127540 3566
rect 127484 3462 127540 3500
rect 127260 3444 127316 3454
rect 127148 3442 127316 3444
rect 127148 3390 127262 3442
rect 127314 3390 127316 3442
rect 127148 3388 127316 3390
rect 127260 3378 127316 3388
rect 127820 800 127876 4284
rect 127932 4274 127988 4284
rect 128268 3892 128324 4398
rect 128268 3826 128324 3836
rect 128044 3444 128100 3454
rect 128044 3350 128100 3388
rect 128604 3332 128660 6414
rect 129724 5906 129780 5918
rect 129724 5854 129726 5906
rect 129778 5854 129780 5906
rect 129276 5796 129332 5806
rect 129724 5796 129780 5854
rect 129276 5794 129780 5796
rect 129276 5742 129278 5794
rect 129330 5742 129780 5794
rect 129276 5740 129780 5742
rect 129276 5730 129332 5740
rect 129052 5012 129108 5022
rect 129052 4918 129108 4956
rect 129388 4340 129444 4350
rect 128940 4228 128996 4238
rect 128828 4226 128996 4228
rect 128828 4174 128942 4226
rect 128994 4174 128996 4226
rect 128828 4172 128996 4174
rect 128828 3556 128884 4172
rect 128940 4162 128996 4172
rect 128828 3490 128884 3500
rect 129388 3556 129444 4284
rect 128940 3442 128996 3454
rect 128940 3390 128942 3442
rect 128994 3390 128996 3442
rect 128940 3332 128996 3390
rect 129388 3442 129444 3500
rect 129388 3390 129390 3442
rect 129442 3390 129444 3442
rect 129388 3378 129444 3390
rect 128604 3276 128996 3332
rect 128940 980 128996 3276
rect 128940 914 128996 924
rect 129500 800 129556 5740
rect 129612 4900 129668 4910
rect 129612 4806 129668 4844
rect 129836 4450 129892 6524
rect 130956 6466 131012 6478
rect 130956 6414 130958 6466
rect 131010 6414 131012 6466
rect 130956 6132 131012 6414
rect 130956 6076 131236 6132
rect 130060 6020 130116 6030
rect 129948 6018 130116 6020
rect 129948 5966 130062 6018
rect 130114 5966 130116 6018
rect 129948 5964 130116 5966
rect 129948 5236 130004 5964
rect 130060 5954 130116 5964
rect 131068 5908 131124 5918
rect 130732 5906 131124 5908
rect 130732 5854 131070 5906
rect 131122 5854 131124 5906
rect 130732 5852 131124 5854
rect 130508 5796 130564 5806
rect 130508 5794 130676 5796
rect 130508 5742 130510 5794
rect 130562 5742 130676 5794
rect 130508 5740 130676 5742
rect 130508 5730 130564 5740
rect 130082 5516 130346 5526
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130082 5450 130346 5460
rect 129948 5180 130452 5236
rect 130172 5012 130228 5022
rect 129836 4398 129838 4450
rect 129890 4398 129892 4450
rect 129836 4386 129892 4398
rect 129948 5010 130228 5012
rect 129948 4958 130174 5010
rect 130226 4958 130228 5010
rect 129948 4956 130228 4958
rect 129612 4340 129668 4350
rect 129612 4246 129668 4284
rect 129724 3892 129780 3902
rect 129724 3778 129780 3836
rect 129724 3726 129726 3778
rect 129778 3726 129780 3778
rect 129724 3714 129780 3726
rect 129948 3780 130004 4956
rect 130172 4946 130228 4956
rect 130396 4338 130452 5180
rect 130508 4898 130564 4910
rect 130508 4846 130510 4898
rect 130562 4846 130564 4898
rect 130508 4676 130564 4846
rect 130620 4900 130676 5740
rect 130620 4834 130676 4844
rect 130508 4610 130564 4620
rect 130732 4562 130788 5852
rect 131068 5842 131124 5852
rect 130732 4510 130734 4562
rect 130786 4510 130788 4562
rect 130732 4498 130788 4510
rect 131068 5010 131124 5022
rect 131068 4958 131070 5010
rect 131122 4958 131124 5010
rect 130396 4286 130398 4338
rect 130450 4286 130452 4338
rect 130396 4274 130452 4286
rect 130082 3948 130346 3958
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130082 3882 130346 3892
rect 130060 3780 130116 3790
rect 129948 3778 130116 3780
rect 129948 3726 130062 3778
rect 130114 3726 130116 3778
rect 129948 3724 130116 3726
rect 130060 3714 130116 3724
rect 131068 3556 131124 4958
rect 131180 3668 131236 6076
rect 131404 6130 131460 30940
rect 131404 6078 131406 6130
rect 131458 6078 131460 6130
rect 131404 6066 131460 6078
rect 131964 5796 132020 5806
rect 132860 5796 132916 5806
rect 131852 5794 132020 5796
rect 131852 5742 131966 5794
rect 132018 5742 132020 5794
rect 131852 5740 132020 5742
rect 131628 4900 131684 4910
rect 131628 4806 131684 4844
rect 131852 4450 131908 5740
rect 131964 5730 132020 5740
rect 132748 5794 132916 5796
rect 132748 5742 132862 5794
rect 132914 5742 132916 5794
rect 132748 5740 132916 5742
rect 132412 5012 132468 5022
rect 132076 4900 132132 4910
rect 132076 4806 132132 4844
rect 131852 4398 131854 4450
rect 131906 4398 131908 4450
rect 131740 4338 131796 4350
rect 131740 4286 131742 4338
rect 131794 4286 131796 4338
rect 131292 3668 131348 3678
rect 131180 3612 131292 3668
rect 131068 3490 131124 3500
rect 131180 3444 131236 3454
rect 131180 800 131236 3388
rect 131292 3442 131348 3612
rect 131404 3556 131460 3566
rect 131404 3462 131460 3500
rect 131740 3556 131796 4286
rect 131740 3490 131796 3500
rect 131292 3390 131294 3442
rect 131346 3390 131348 3442
rect 131292 3378 131348 3390
rect 131852 2996 131908 4398
rect 132412 3778 132468 4956
rect 132412 3726 132414 3778
rect 132466 3726 132468 3778
rect 132412 3714 132468 3726
rect 132524 4114 132580 4126
rect 132524 4062 132526 4114
rect 132578 4062 132580 4114
rect 132076 3554 132132 3566
rect 132076 3502 132078 3554
rect 132130 3502 132132 3554
rect 132076 3332 132132 3502
rect 132076 3266 132132 3276
rect 132524 3220 132580 4062
rect 132748 3444 132804 5740
rect 132860 5730 132916 5740
rect 133756 5794 133812 5806
rect 133756 5742 133758 5794
rect 133810 5742 133812 5794
rect 133756 5684 133812 5742
rect 133756 5628 134036 5684
rect 133084 5236 133140 5246
rect 132972 5012 133028 5022
rect 132972 4918 133028 4956
rect 133084 4788 133140 5180
rect 133308 5236 133364 5246
rect 133308 5010 133364 5180
rect 133308 4958 133310 5010
rect 133362 4958 133364 5010
rect 133308 4946 133364 4958
rect 133868 5010 133924 5022
rect 133868 4958 133870 5010
rect 133922 4958 133924 5010
rect 133084 4732 133588 4788
rect 132860 4564 132916 4574
rect 132860 4470 132916 4508
rect 133532 4450 133588 4732
rect 133868 4564 133924 4958
rect 133868 4498 133924 4508
rect 133532 4398 133534 4450
rect 133586 4398 133588 4450
rect 133532 4386 133588 4398
rect 133980 3556 134036 5628
rect 134092 5012 134148 5022
rect 134092 4562 134148 4956
rect 134204 5010 134260 33292
rect 136892 31556 136948 31566
rect 135212 27188 135268 27198
rect 135212 10948 135268 27132
rect 135324 24612 135380 24622
rect 135324 19348 135380 24556
rect 135324 19282 135380 19292
rect 135212 10882 135268 10892
rect 134876 8148 134932 8158
rect 134876 8054 134932 8092
rect 135324 8148 135380 8158
rect 135324 8054 135380 8092
rect 134540 8034 134596 8046
rect 134540 7982 134542 8034
rect 134594 7982 134596 8034
rect 134540 5236 134596 7982
rect 136556 6244 136612 6254
rect 134652 5236 134708 5246
rect 134540 5234 134708 5236
rect 134540 5182 134654 5234
rect 134706 5182 134708 5234
rect 134540 5180 134708 5182
rect 134204 4958 134206 5010
rect 134258 4958 134260 5010
rect 134204 4946 134260 4958
rect 134652 5012 134708 5180
rect 136108 5124 136164 5134
rect 135996 5122 136164 5124
rect 135996 5070 136110 5122
rect 136162 5070 136164 5122
rect 135996 5068 136164 5070
rect 134652 4946 134708 4956
rect 135548 5012 135604 5022
rect 135100 4900 135156 4910
rect 134092 4510 134094 4562
rect 134146 4510 134148 4562
rect 134092 4498 134148 4510
rect 134988 4898 135156 4900
rect 134988 4846 135102 4898
rect 135154 4846 135156 4898
rect 134988 4844 135156 4846
rect 134764 4340 134820 4350
rect 134988 4340 135044 4844
rect 135100 4834 135156 4844
rect 135548 4564 135604 4956
rect 135660 4564 135716 4574
rect 135548 4562 135716 4564
rect 135548 4510 135662 4562
rect 135714 4510 135716 4562
rect 135548 4508 135716 4510
rect 135660 4498 135716 4508
rect 135100 4452 135156 4462
rect 135100 4358 135156 4396
rect 134540 4338 135044 4340
rect 134540 4286 134766 4338
rect 134818 4286 135044 4338
rect 134540 4284 135044 4286
rect 134204 3556 134260 3566
rect 133980 3554 134260 3556
rect 133980 3502 134206 3554
rect 134258 3502 134260 3554
rect 133980 3500 134260 3502
rect 132748 3378 132804 3388
rect 133420 3444 133476 3454
rect 133420 3350 133476 3388
rect 133084 3332 133140 3342
rect 133084 3238 133140 3276
rect 133980 3330 134036 3342
rect 133980 3278 133982 3330
rect 134034 3278 134036 3330
rect 132524 3154 132580 3164
rect 133980 3220 134036 3278
rect 133980 3154 134036 3164
rect 131852 2930 131908 2940
rect 132860 924 133252 980
rect 132860 800 132916 924
rect 113036 700 113988 756
rect 114352 0 114464 800
rect 116032 0 116144 800
rect 117712 0 117824 800
rect 119392 0 119504 800
rect 121072 0 121184 800
rect 122752 0 122864 800
rect 124432 0 124544 800
rect 126112 0 126224 800
rect 127792 0 127904 800
rect 129472 0 129584 800
rect 131152 0 131264 800
rect 132832 0 132944 800
rect 133196 756 133252 924
rect 134204 756 134260 3500
rect 134540 800 134596 4284
rect 134764 4274 134820 4284
rect 135548 3444 135604 3454
rect 135996 3444 136052 5068
rect 136108 5058 136164 5068
rect 136332 4452 136388 4462
rect 135548 3442 136052 3444
rect 135548 3390 135550 3442
rect 135602 3390 136052 3442
rect 135548 3388 136052 3390
rect 136108 4340 136164 4350
rect 136108 4226 136164 4284
rect 136108 4174 136110 4226
rect 136162 4174 136164 4226
rect 136108 3442 136164 4174
rect 136332 3778 136388 4396
rect 136332 3726 136334 3778
rect 136386 3726 136388 3778
rect 136332 3714 136388 3726
rect 136444 3668 136500 3678
rect 136108 3390 136110 3442
rect 136162 3390 136164 3442
rect 135548 1540 135604 3388
rect 136108 3378 136164 3390
rect 136220 3444 136276 3454
rect 135548 1474 135604 1484
rect 136220 800 136276 3388
rect 136444 2100 136500 3612
rect 136556 3220 136612 6188
rect 136892 5236 136948 31500
rect 139244 28644 139300 28654
rect 139244 27748 139300 28588
rect 139244 27682 139300 27692
rect 136892 5170 136948 5180
rect 137788 6804 137844 6814
rect 137452 5012 137508 5022
rect 136892 5010 137508 5012
rect 136892 4958 137454 5010
rect 137506 4958 137508 5010
rect 136892 4956 137508 4958
rect 136780 4898 136836 4910
rect 136780 4846 136782 4898
rect 136834 4846 136836 4898
rect 136780 4452 136836 4846
rect 136780 4386 136836 4396
rect 136892 4116 136948 4956
rect 137452 4946 137508 4956
rect 137788 5010 137844 6748
rect 139356 6692 139412 33964
rect 140812 33908 140868 33918
rect 139356 6636 139524 6692
rect 138796 5796 138852 5806
rect 138796 5794 139412 5796
rect 138796 5742 138798 5794
rect 138850 5742 139412 5794
rect 138796 5740 139412 5742
rect 138796 5730 138852 5740
rect 137788 4958 137790 5010
rect 137842 4958 137844 5010
rect 137788 4946 137844 4958
rect 139132 5010 139188 5022
rect 139132 4958 139134 5010
rect 139186 4958 139188 5010
rect 138684 4898 138740 4910
rect 138684 4846 138686 4898
rect 138738 4846 138740 4898
rect 138236 4676 138292 4686
rect 138236 4562 138292 4620
rect 138236 4510 138238 4562
rect 138290 4510 138292 4562
rect 138236 4498 138292 4510
rect 137228 4452 137284 4462
rect 137116 4340 137172 4350
rect 137116 4246 137172 4284
rect 136668 4060 136948 4116
rect 137228 4116 137284 4396
rect 138684 4452 138740 4846
rect 139132 4676 139188 4958
rect 139132 4610 139188 4620
rect 139132 4452 139188 4462
rect 138684 4450 139188 4452
rect 138684 4398 139134 4450
rect 139186 4398 139188 4450
rect 138684 4396 139188 4398
rect 137900 4116 137956 4126
rect 136668 3778 136724 4060
rect 137228 4050 137284 4060
rect 137676 4114 137956 4116
rect 137676 4062 137902 4114
rect 137954 4062 137956 4114
rect 137676 4060 137956 4062
rect 136668 3726 136670 3778
rect 136722 3726 136724 3778
rect 136668 3714 136724 3726
rect 137340 3444 137396 3454
rect 137340 3350 137396 3388
rect 137676 3330 137732 4060
rect 137900 4050 137956 4060
rect 137676 3278 137678 3330
rect 137730 3278 137732 3330
rect 137676 3266 137732 3278
rect 137900 3556 137956 3566
rect 136556 3154 136612 3164
rect 136444 2034 136500 2044
rect 137900 800 137956 3500
rect 138124 3444 138180 3454
rect 138124 3350 138180 3388
rect 138684 2212 138740 4396
rect 139132 4386 139188 4396
rect 139356 3668 139412 5740
rect 139468 5010 139524 6636
rect 140812 6130 140868 33852
rect 140812 6078 140814 6130
rect 140866 6078 140868 6130
rect 140812 6066 140868 6078
rect 140924 6466 140980 6478
rect 140924 6414 140926 6466
rect 140978 6414 140980 6466
rect 140140 5908 140196 5918
rect 140476 5908 140532 5918
rect 139468 4958 139470 5010
rect 139522 4958 139524 5010
rect 139468 4946 139524 4958
rect 139580 5794 139636 5806
rect 139580 5742 139582 5794
rect 139634 5742 139636 5794
rect 139580 4676 139636 5742
rect 139916 5796 139972 5806
rect 139916 5702 139972 5740
rect 139356 3442 139412 3612
rect 139356 3390 139358 3442
rect 139410 3390 139412 3442
rect 139356 3378 139412 3390
rect 139468 4620 139636 4676
rect 139692 4900 139748 4910
rect 139468 3332 139524 4620
rect 139580 4452 139636 4462
rect 139580 3442 139636 4396
rect 139692 3892 139748 4844
rect 140140 4564 140196 5852
rect 140364 5906 140532 5908
rect 140364 5854 140478 5906
rect 140530 5854 140532 5906
rect 140364 5852 140532 5854
rect 140252 5122 140308 5134
rect 140252 5070 140254 5122
rect 140306 5070 140308 5122
rect 140252 4900 140308 5070
rect 140252 4834 140308 4844
rect 140252 4564 140308 4574
rect 140140 4562 140308 4564
rect 140140 4510 140254 4562
rect 140306 4510 140308 4562
rect 140140 4508 140308 4510
rect 140252 4498 140308 4508
rect 139916 4116 139972 4126
rect 139916 4114 140084 4116
rect 139916 4062 139918 4114
rect 139970 4062 140084 4114
rect 139916 4060 140084 4062
rect 139916 4050 139972 4060
rect 139692 3826 139748 3836
rect 139916 3554 139972 3566
rect 139916 3502 139918 3554
rect 139970 3502 139972 3554
rect 139580 3390 139582 3442
rect 139634 3390 139636 3442
rect 139580 3378 139636 3390
rect 139692 3444 139748 3454
rect 139468 3108 139524 3276
rect 139468 3042 139524 3052
rect 139692 2548 139748 3388
rect 139916 2994 139972 3502
rect 140028 3332 140084 4060
rect 140252 3780 140308 3790
rect 140364 3780 140420 5852
rect 140476 5842 140532 5852
rect 140924 5796 140980 6414
rect 140924 5124 140980 5740
rect 140924 5058 140980 5068
rect 141260 6466 141316 6478
rect 141260 6414 141262 6466
rect 141314 6414 141316 6466
rect 141148 5010 141204 5022
rect 141148 4958 141150 5010
rect 141202 4958 141204 5010
rect 141148 4900 141204 4958
rect 141148 4834 141204 4844
rect 141148 4450 141204 4462
rect 141148 4398 141150 4450
rect 141202 4398 141204 4450
rect 141148 4116 141204 4398
rect 140252 3778 140420 3780
rect 140252 3726 140254 3778
rect 140306 3726 140420 3778
rect 140252 3724 140420 3726
rect 141036 4060 141204 4116
rect 140252 3714 140308 3724
rect 140028 3266 140084 3276
rect 140924 3330 140980 3342
rect 140924 3278 140926 3330
rect 140978 3278 140980 3330
rect 139916 2942 139918 2994
rect 139970 2942 139972 2994
rect 139916 2930 139972 2942
rect 140924 2994 140980 3278
rect 141036 3108 141092 4060
rect 141148 3556 141204 3566
rect 141260 3556 141316 6414
rect 141708 6130 141764 36204
rect 143836 36260 143892 36270
rect 144284 36260 144340 36428
rect 144844 36484 144900 36494
rect 144844 36390 144900 36428
rect 143836 36166 143892 36204
rect 144060 36258 144340 36260
rect 144060 36206 144286 36258
rect 144338 36206 144340 36258
rect 144060 36204 144340 36206
rect 141708 6078 141710 6130
rect 141762 6078 141764 6130
rect 141708 6066 141764 6078
rect 142604 35588 142660 35598
rect 142604 6130 142660 35532
rect 142604 6078 142606 6130
rect 142658 6078 142660 6130
rect 142604 6066 142660 6078
rect 143164 33572 143220 33582
rect 141372 5908 141428 5918
rect 141372 5814 141428 5852
rect 142268 5906 142324 5918
rect 142268 5854 142270 5906
rect 142322 5854 142324 5906
rect 142156 5348 142212 5358
rect 142268 5348 142324 5854
rect 142156 5346 142324 5348
rect 142156 5294 142158 5346
rect 142210 5294 142324 5346
rect 142156 5292 142324 5294
rect 143052 5794 143108 5806
rect 143052 5742 143054 5794
rect 143106 5742 143108 5794
rect 142156 5282 142212 5292
rect 141596 5124 141652 5134
rect 141596 5010 141652 5068
rect 141596 4958 141598 5010
rect 141650 4958 141652 5010
rect 141596 4450 141652 4958
rect 141820 5122 141876 5134
rect 141820 5070 141822 5122
rect 141874 5070 141876 5122
rect 141820 4676 141876 5070
rect 141820 4610 141876 4620
rect 142828 5010 142884 5022
rect 142828 4958 142830 5010
rect 142882 4958 142884 5010
rect 142156 4564 142212 4574
rect 142156 4470 142212 4508
rect 142828 4564 142884 4958
rect 142828 4498 142884 4508
rect 141596 4398 141598 4450
rect 141650 4398 141652 4450
rect 141596 4386 141652 4398
rect 142828 4338 142884 4350
rect 142828 4286 142830 4338
rect 142882 4286 142884 4338
rect 141204 3500 141316 3556
rect 141372 4228 141428 4238
rect 141148 3462 141204 3500
rect 141372 3220 141428 4172
rect 142828 4228 142884 4286
rect 142828 4162 142884 4172
rect 142940 4340 142996 4350
rect 141820 4116 141876 4126
rect 141820 4114 142100 4116
rect 141820 4062 141822 4114
rect 141874 4062 142100 4114
rect 141820 4060 142100 4062
rect 141820 4050 141876 4060
rect 141820 3332 141876 3342
rect 141820 3238 141876 3276
rect 142044 3332 142100 4060
rect 142156 3444 142212 3454
rect 142156 3350 142212 3388
rect 142044 3266 142100 3276
rect 141036 3042 141092 3052
rect 141260 3164 141428 3220
rect 140924 2942 140926 2994
rect 140978 2942 140980 2994
rect 140924 2930 140980 2942
rect 138684 2146 138740 2156
rect 139580 2492 139748 2548
rect 139580 800 139636 2492
rect 141260 800 141316 3164
rect 142940 800 142996 4284
rect 143052 4228 143108 5742
rect 143164 5010 143220 33516
rect 143164 4958 143166 5010
rect 143218 4958 143220 5010
rect 143164 4946 143220 4958
rect 143276 6916 143332 6926
rect 143052 4162 143108 4172
rect 143164 4450 143220 4462
rect 143164 4398 143166 4450
rect 143218 4398 143220 4450
rect 143164 3780 143220 4398
rect 143164 3714 143220 3724
rect 143276 4228 143332 6860
rect 143276 3442 143332 4172
rect 143276 3390 143278 3442
rect 143330 3390 143332 3442
rect 143276 3378 143332 3390
rect 143500 5794 143556 5806
rect 143500 5742 143502 5794
rect 143554 5742 143556 5794
rect 143500 5124 143556 5742
rect 143500 3442 143556 5068
rect 143724 5012 143780 5022
rect 143724 5010 144004 5012
rect 143724 4958 143726 5010
rect 143778 4958 144004 5010
rect 143724 4956 144004 4958
rect 143724 4946 143780 4956
rect 143724 4676 143780 4686
rect 143724 4562 143780 4620
rect 143724 4510 143726 4562
rect 143778 4510 143780 4562
rect 143724 4498 143780 4510
rect 143948 4116 144004 4956
rect 144060 5010 144116 36204
rect 144284 36194 144340 36204
rect 145964 35810 146020 37884
rect 145964 35758 145966 35810
rect 146018 35758 146020 35810
rect 145964 35746 146020 35758
rect 145068 35698 145124 35710
rect 145068 35646 145070 35698
rect 145122 35646 145124 35698
rect 144284 35588 144340 35598
rect 144284 35494 144340 35532
rect 145068 35588 145124 35646
rect 145068 35522 145124 35532
rect 146076 35026 146132 38780
rect 146860 36482 146916 36494
rect 146860 36430 146862 36482
rect 146914 36430 146916 36482
rect 146860 36260 146916 36430
rect 146860 36194 146916 36204
rect 147756 36370 147812 36382
rect 147756 36318 147758 36370
rect 147810 36318 147812 36370
rect 147756 36260 147812 36318
rect 147756 36194 147812 36204
rect 148492 36092 148756 36102
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148492 36026 148756 36036
rect 146076 34974 146078 35026
rect 146130 34974 146132 35026
rect 146076 34962 146132 34974
rect 146972 35698 147028 35710
rect 146972 35646 146974 35698
rect 147026 35646 147028 35698
rect 145068 34916 145124 34926
rect 144508 34914 145124 34916
rect 144508 34862 145070 34914
rect 145122 34862 145124 34914
rect 144508 34860 145124 34862
rect 144508 34690 144564 34860
rect 145068 34850 145124 34860
rect 146860 34914 146916 34926
rect 146860 34862 146862 34914
rect 146914 34862 146916 34914
rect 144508 34638 144510 34690
rect 144562 34638 144564 34690
rect 144508 33572 144564 34638
rect 146412 34132 146468 34142
rect 146412 34038 146468 34076
rect 145404 34018 145460 34030
rect 145404 33966 145406 34018
rect 145458 33966 145460 34018
rect 145404 33908 145460 33966
rect 145852 34020 145908 34030
rect 145852 33926 145908 33964
rect 146860 34020 146916 34862
rect 146860 33954 146916 33964
rect 145404 33842 145460 33852
rect 146972 33908 147028 35646
rect 147756 35586 147812 35598
rect 147756 35534 147758 35586
rect 147810 35534 147812 35586
rect 147756 35364 147812 35534
rect 147756 35298 147812 35308
rect 147756 34802 147812 34814
rect 147756 34750 147758 34802
rect 147810 34750 147812 34802
rect 147756 34356 147812 34750
rect 148492 34524 148756 34534
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148492 34458 148756 34468
rect 147756 34290 147812 34300
rect 147084 34132 147140 34142
rect 147084 34038 147140 34076
rect 147868 34132 147924 34142
rect 146972 33842 147028 33852
rect 147756 34018 147812 34030
rect 147756 33966 147758 34018
rect 147810 33966 147812 34018
rect 147756 33684 147812 33966
rect 147756 33618 147812 33628
rect 144508 33506 144564 33516
rect 146300 33348 146356 33358
rect 146300 33254 146356 33292
rect 146860 33348 146916 33358
rect 146860 33254 146916 33292
rect 147756 33234 147812 33246
rect 147756 33182 147758 33234
rect 147810 33182 147812 33234
rect 147756 32564 147812 33182
rect 147756 32498 147812 32508
rect 146860 31778 146916 31790
rect 146860 31726 146862 31778
rect 146914 31726 146916 31778
rect 146300 31556 146356 31566
rect 146300 31462 146356 31500
rect 146860 31556 146916 31726
rect 147756 31668 147812 31678
rect 147756 31574 147812 31612
rect 146860 31490 146916 31500
rect 146412 30996 146468 31006
rect 146412 30902 146468 30940
rect 146860 30996 146916 31006
rect 146860 30902 146916 30940
rect 147756 30882 147812 30894
rect 147756 30830 147758 30882
rect 147810 30830 147812 30882
rect 147756 30772 147812 30830
rect 147756 30706 147812 30716
rect 146300 30212 146356 30222
rect 146300 30118 146356 30156
rect 147084 30212 147140 30222
rect 147084 30118 147140 30156
rect 147756 30098 147812 30110
rect 147756 30046 147758 30098
rect 147810 30046 147812 30098
rect 147756 29988 147812 30046
rect 147756 29922 147812 29932
rect 146412 29428 146468 29438
rect 146412 29334 146468 29372
rect 146860 29428 146916 29438
rect 146860 29334 146916 29372
rect 147756 29314 147812 29326
rect 147756 29262 147758 29314
rect 147810 29262 147812 29314
rect 147756 28980 147812 29262
rect 147756 28914 147812 28924
rect 146300 28644 146356 28654
rect 146300 28550 146356 28588
rect 146860 28644 146916 28654
rect 146860 28550 146916 28588
rect 147756 28642 147812 28654
rect 147756 28590 147758 28642
rect 147810 28590 147812 28642
rect 147756 28084 147812 28590
rect 147756 28018 147812 28028
rect 146412 27860 146468 27870
rect 146412 27766 146468 27804
rect 147084 27860 147140 27870
rect 147084 27766 147140 27804
rect 147756 27746 147812 27758
rect 147756 27694 147758 27746
rect 147810 27694 147812 27746
rect 146300 27188 146356 27198
rect 146300 27094 146356 27132
rect 146860 27188 146916 27198
rect 146860 27074 146916 27132
rect 147756 27188 147812 27694
rect 147756 27122 147812 27132
rect 146860 27022 146862 27074
rect 146914 27022 146916 27074
rect 146860 27010 146916 27022
rect 147756 26962 147812 26974
rect 147756 26910 147758 26962
rect 147810 26910 147812 26962
rect 147756 26292 147812 26910
rect 147756 26226 147812 26236
rect 146860 25506 146916 25518
rect 146860 25454 146862 25506
rect 146914 25454 146916 25506
rect 146300 25284 146356 25294
rect 146300 25190 146356 25228
rect 146860 25284 146916 25454
rect 147756 25396 147812 25406
rect 147756 25302 147812 25340
rect 146860 25218 146916 25228
rect 146860 24722 146916 24734
rect 146860 24670 146862 24722
rect 146914 24670 146916 24722
rect 146412 24612 146468 24622
rect 146412 24518 146468 24556
rect 146860 24612 146916 24670
rect 146860 24546 146916 24556
rect 147756 24610 147812 24622
rect 147756 24558 147758 24610
rect 147810 24558 147812 24610
rect 147756 24500 147812 24558
rect 147756 24434 147812 24444
rect 146860 23938 146916 23950
rect 146860 23886 146862 23938
rect 146914 23886 146916 23938
rect 146300 23716 146356 23726
rect 146300 23622 146356 23660
rect 146860 23716 146916 23886
rect 146860 23650 146916 23660
rect 147756 23826 147812 23838
rect 147756 23774 147758 23826
rect 147810 23774 147812 23826
rect 147756 23716 147812 23774
rect 147756 23650 147812 23660
rect 146412 23156 146468 23166
rect 146412 23062 146468 23100
rect 146860 23156 146916 23166
rect 146860 23062 146916 23100
rect 147756 23042 147812 23054
rect 147756 22990 147758 23042
rect 147810 22990 147812 23042
rect 147756 22708 147812 22990
rect 147756 22642 147812 22652
rect 146300 22372 146356 22382
rect 146300 22278 146356 22316
rect 146860 22372 146916 22382
rect 146860 22278 146916 22316
rect 147756 22258 147812 22270
rect 147756 22206 147758 22258
rect 147810 22206 147812 22258
rect 147756 21924 147812 22206
rect 147756 21858 147812 21868
rect 146860 21586 146916 21598
rect 146860 21534 146862 21586
rect 146914 21534 146916 21586
rect 146412 21476 146468 21486
rect 146412 21382 146468 21420
rect 146860 21476 146916 21534
rect 146860 21410 146916 21420
rect 147756 21474 147812 21486
rect 147756 21422 147758 21474
rect 147810 21422 147812 21474
rect 147756 20916 147812 21422
rect 147756 20850 147812 20860
rect 146300 20804 146356 20814
rect 146300 20710 146356 20748
rect 146860 20804 146916 20814
rect 146860 20710 146916 20748
rect 147756 20690 147812 20702
rect 147756 20638 147758 20690
rect 147810 20638 147812 20690
rect 147756 20244 147812 20638
rect 147756 20178 147812 20188
rect 146300 19236 146356 19246
rect 146300 19142 146356 19180
rect 146860 19236 146916 19246
rect 146860 19142 146916 19180
rect 147756 19124 147812 19134
rect 147756 19030 147812 19068
rect 146860 18450 146916 18462
rect 146860 18398 146862 18450
rect 146914 18398 146916 18450
rect 146412 18340 146468 18350
rect 146412 18246 146468 18284
rect 146860 18340 146916 18398
rect 146860 18274 146916 18284
rect 147756 18338 147812 18350
rect 147756 18286 147758 18338
rect 147810 18286 147812 18338
rect 147756 18228 147812 18286
rect 147756 18162 147812 18172
rect 146860 17666 146916 17678
rect 146860 17614 146862 17666
rect 146914 17614 146916 17666
rect 146300 17444 146356 17454
rect 146300 17350 146356 17388
rect 146860 17444 146916 17614
rect 146860 17378 146916 17388
rect 147756 17554 147812 17566
rect 147756 17502 147758 17554
rect 147810 17502 147812 17554
rect 147756 17444 147812 17502
rect 147756 17378 147812 17388
rect 146412 16996 146468 17006
rect 146412 16902 146468 16940
rect 146860 16996 146916 17006
rect 146860 16882 146916 16940
rect 146860 16830 146862 16882
rect 146914 16830 146916 16882
rect 146860 16818 146916 16830
rect 147756 16882 147812 16894
rect 147756 16830 147758 16882
rect 147810 16830 147812 16882
rect 147756 16436 147812 16830
rect 147756 16370 147812 16380
rect 146860 16098 146916 16110
rect 146860 16046 146862 16098
rect 146914 16046 146916 16098
rect 146300 15876 146356 15886
rect 146300 15782 146356 15820
rect 146860 15876 146916 16046
rect 146860 15810 146916 15820
rect 147756 15986 147812 15998
rect 147756 15934 147758 15986
rect 147810 15934 147812 15986
rect 147756 15540 147812 15934
rect 147756 15474 147812 15484
rect 146412 15428 146468 15438
rect 146412 15334 146468 15372
rect 146860 15428 146916 15438
rect 146860 15314 146916 15372
rect 146860 15262 146862 15314
rect 146914 15262 146916 15314
rect 146860 15250 146916 15262
rect 147756 15202 147812 15214
rect 147756 15150 147758 15202
rect 147810 15150 147812 15202
rect 147756 14644 147812 15150
rect 147756 14578 147812 14588
rect 146300 14532 146356 14542
rect 146300 14438 146356 14476
rect 146860 14532 146916 14542
rect 146860 14438 146916 14476
rect 147756 14418 147812 14430
rect 147756 14366 147758 14418
rect 147810 14366 147812 14418
rect 147756 13748 147812 14366
rect 147756 13682 147812 13692
rect 146300 12964 146356 12974
rect 146300 12870 146356 12908
rect 146860 12964 146916 12974
rect 146860 12870 146916 12908
rect 147756 12852 147812 12862
rect 147756 12758 147812 12796
rect 146860 12178 146916 12190
rect 146860 12126 146862 12178
rect 146914 12126 146916 12178
rect 146412 12068 146468 12078
rect 146412 11974 146468 12012
rect 146860 12068 146916 12126
rect 146860 12002 146916 12012
rect 147756 12066 147812 12078
rect 147756 12014 147758 12066
rect 147810 12014 147812 12066
rect 147756 11956 147812 12014
rect 147756 11890 147812 11900
rect 146300 11396 146356 11406
rect 146300 11302 146356 11340
rect 146860 11396 146916 11406
rect 146860 11302 146916 11340
rect 147756 11282 147812 11294
rect 147756 11230 147758 11282
rect 147810 11230 147812 11282
rect 147756 11172 147812 11230
rect 147756 11106 147812 11116
rect 147756 10724 147812 10734
rect 147532 10722 147812 10724
rect 147532 10670 147758 10722
rect 147810 10670 147812 10722
rect 147532 10668 147812 10670
rect 147308 10498 147364 10510
rect 147308 10446 147310 10498
rect 147362 10446 147364 10498
rect 147308 10164 147364 10446
rect 147308 10098 147364 10108
rect 147308 9602 147364 9614
rect 147308 9550 147310 9602
rect 147362 9550 147364 9602
rect 147308 9268 147364 9550
rect 147308 9202 147364 9212
rect 147308 9044 147364 9054
rect 147308 8950 147364 8988
rect 147532 8148 147588 10668
rect 147756 10658 147812 10668
rect 147756 9604 147812 9614
rect 147644 9602 147812 9604
rect 147644 9550 147758 9602
rect 147810 9550 147812 9602
rect 147644 9548 147812 9550
rect 147644 8820 147700 9548
rect 147756 9538 147812 9548
rect 147756 9156 147812 9166
rect 147756 9062 147812 9100
rect 147644 8754 147700 8764
rect 147532 8082 147588 8092
rect 147308 8036 147364 8046
rect 147308 7942 147364 7980
rect 147756 8034 147812 8046
rect 147756 7982 147758 8034
rect 147810 7982 147812 8034
rect 144060 4958 144062 5010
rect 144114 4958 144116 5010
rect 144060 4946 144116 4958
rect 146076 7364 146132 7374
rect 146076 4564 146132 7308
rect 147756 7252 147812 7982
rect 147756 7186 147812 7196
rect 147868 6804 147924 34076
rect 148492 32956 148756 32966
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148492 32890 148756 32900
rect 148492 31388 148756 31398
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148492 31322 148756 31332
rect 147868 6738 147924 6748
rect 147980 30212 148036 30222
rect 147644 6692 147700 6702
rect 147308 6580 147364 6590
rect 147308 6486 147364 6524
rect 147308 5794 147364 5806
rect 147308 5742 147310 5794
rect 147362 5742 147364 5794
rect 147308 5684 147364 5742
rect 147308 5618 147364 5628
rect 146412 5124 146468 5134
rect 146412 5122 146580 5124
rect 146412 5070 146414 5122
rect 146466 5070 146580 5122
rect 146412 5068 146580 5070
rect 146412 5058 146468 5068
rect 146076 4498 146132 4508
rect 145180 4452 145236 4462
rect 144060 4340 144116 4350
rect 144060 4246 144116 4284
rect 144844 4228 144900 4238
rect 144844 4134 144900 4172
rect 143948 4060 144228 4116
rect 143836 3780 143892 3790
rect 143836 3686 143892 3724
rect 144172 3778 144228 4060
rect 144172 3726 144174 3778
rect 144226 3726 144228 3778
rect 144172 3714 144228 3726
rect 145068 3556 145124 3566
rect 143500 3390 143502 3442
rect 143554 3390 143556 3442
rect 143500 3378 143556 3390
rect 144620 3554 145124 3556
rect 144620 3502 145070 3554
rect 145122 3502 145124 3554
rect 144620 3500 145124 3502
rect 144620 800 144676 3500
rect 145068 3444 145124 3500
rect 145068 3378 145124 3388
rect 144844 3332 144900 3342
rect 144844 3238 144900 3276
rect 145180 868 145236 4396
rect 145292 4340 145348 4350
rect 145292 4246 145348 4284
rect 145964 4226 146020 4238
rect 145964 4174 145966 4226
rect 146018 4174 146020 4226
rect 145964 3892 146020 4174
rect 146412 4228 146468 4238
rect 146412 4134 146468 4172
rect 145964 3826 146020 3836
rect 145628 3556 145684 3566
rect 145628 3462 145684 3500
rect 146076 3444 146132 3454
rect 146076 3350 146132 3388
rect 146524 3444 146580 5068
rect 147308 5122 147364 5134
rect 147308 5070 147310 5122
rect 147362 5070 147364 5122
rect 146860 4900 146916 4910
rect 147308 4900 147364 5070
rect 146860 4898 147252 4900
rect 146860 4846 146862 4898
rect 146914 4846 147252 4898
rect 146860 4844 147252 4846
rect 146860 4834 146916 4844
rect 146860 4452 146916 4462
rect 146860 4358 146916 4396
rect 146524 3378 146580 3388
rect 147084 4338 147140 4350
rect 147084 4286 147086 4338
rect 147138 4286 147140 4338
rect 147084 4228 147140 4286
rect 146860 3330 146916 3342
rect 146860 3278 146862 3330
rect 146914 3278 146916 3330
rect 146860 3220 146916 3278
rect 146860 3154 146916 3164
rect 147084 2996 147140 4172
rect 147084 2930 147140 2940
rect 147196 3442 147252 4844
rect 147308 4834 147364 4844
rect 147196 3390 147198 3442
rect 147250 3390 147252 3442
rect 147196 1204 147252 3390
rect 147644 3332 147700 6636
rect 147756 6466 147812 6478
rect 147756 6414 147758 6466
rect 147810 6414 147812 6466
rect 147756 6356 147812 6414
rect 147756 6290 147812 6300
rect 147756 6020 147812 6030
rect 147756 5926 147812 5964
rect 147756 4898 147812 4910
rect 147756 4846 147758 4898
rect 147810 4846 147812 4898
rect 147756 4788 147812 4846
rect 147756 4722 147812 4732
rect 147980 4676 148036 30156
rect 148492 29820 148756 29830
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148492 29754 148756 29764
rect 148492 28252 148756 28262
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148492 28186 148756 28196
rect 148204 27860 148260 27870
rect 148092 10610 148148 10622
rect 148092 10558 148094 10610
rect 148146 10558 148148 10610
rect 148092 10164 148148 10558
rect 148092 10098 148148 10108
rect 148092 9714 148148 9726
rect 148092 9662 148094 9714
rect 148146 9662 148148 9714
rect 148092 9268 148148 9662
rect 148092 9202 148148 9212
rect 148092 9044 148148 9054
rect 148092 8484 148148 8988
rect 148092 8418 148148 8428
rect 148092 8146 148148 8158
rect 148092 8094 148094 8146
rect 148146 8094 148148 8146
rect 148092 8036 148148 8094
rect 148092 7476 148148 7980
rect 148204 7588 148260 27804
rect 148492 26684 148756 26694
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148492 26618 148756 26628
rect 148492 25116 148756 25126
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148492 25050 148756 25060
rect 148492 23548 148756 23558
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148492 23482 148756 23492
rect 148492 21980 148756 21990
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148492 21914 148756 21924
rect 148492 20412 148756 20422
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148492 20346 148756 20356
rect 148492 18844 148756 18854
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148492 18778 148756 18788
rect 148492 17276 148756 17286
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148492 17210 148756 17220
rect 148492 15708 148756 15718
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148492 15642 148756 15652
rect 148492 14140 148756 14150
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148492 14074 148756 14084
rect 148492 12572 148756 12582
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148492 12506 148756 12516
rect 148492 11004 148756 11014
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148492 10938 148756 10948
rect 148492 9436 148756 9446
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148492 9370 148756 9380
rect 148492 7868 148756 7878
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148492 7802 148756 7812
rect 148204 7522 148260 7532
rect 148092 7410 148148 7420
rect 148092 6580 148148 6590
rect 148092 6486 148148 6524
rect 148492 6300 148756 6310
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148492 6234 148756 6244
rect 148092 5906 148148 5918
rect 148092 5854 148094 5906
rect 148146 5854 148148 5906
rect 148092 5684 148148 5854
rect 148092 5618 148148 5628
rect 148092 5010 148148 5022
rect 148092 4958 148094 5010
rect 148146 4958 148148 5010
rect 148092 4900 148148 4958
rect 148092 4834 148148 4844
rect 148492 4732 148756 4742
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148492 4666 148756 4676
rect 147980 4610 148036 4620
rect 147756 4564 147812 4574
rect 147756 4470 147812 4508
rect 148092 4338 148148 4350
rect 148092 4286 148094 4338
rect 148146 4286 148148 4338
rect 148092 3892 148148 4286
rect 148092 3826 148148 3836
rect 148092 3444 148148 3454
rect 147756 3332 147812 3342
rect 147644 3330 147812 3332
rect 147644 3278 147758 3330
rect 147810 3278 147812 3330
rect 147644 3276 147812 3278
rect 147756 3266 147812 3276
rect 148092 2100 148148 3388
rect 148492 3164 148756 3174
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148492 3098 148756 3108
rect 148092 2034 148148 2044
rect 147196 1138 147252 1148
rect 145180 802 145236 812
rect 133196 700 134260 756
rect 134512 0 134624 800
rect 136192 0 136304 800
rect 137872 0 137984 800
rect 139552 0 139664 800
rect 141232 0 141344 800
rect 142912 0 143024 800
rect 144592 0 144704 800
<< via2 >>
rect 146076 38780 146132 38836
rect 145964 37884 146020 37940
rect 145852 36988 145908 37044
rect 19622 36874 19678 36876
rect 19622 36822 19624 36874
rect 19624 36822 19676 36874
rect 19676 36822 19678 36874
rect 19622 36820 19678 36822
rect 19726 36874 19782 36876
rect 19726 36822 19728 36874
rect 19728 36822 19780 36874
rect 19780 36822 19782 36874
rect 19726 36820 19782 36822
rect 19830 36874 19886 36876
rect 19830 36822 19832 36874
rect 19832 36822 19884 36874
rect 19884 36822 19886 36874
rect 19830 36820 19886 36822
rect 56442 36874 56498 36876
rect 56442 36822 56444 36874
rect 56444 36822 56496 36874
rect 56496 36822 56498 36874
rect 56442 36820 56498 36822
rect 56546 36874 56602 36876
rect 56546 36822 56548 36874
rect 56548 36822 56600 36874
rect 56600 36822 56602 36874
rect 56546 36820 56602 36822
rect 56650 36874 56706 36876
rect 56650 36822 56652 36874
rect 56652 36822 56704 36874
rect 56704 36822 56706 36874
rect 56650 36820 56706 36822
rect 93262 36874 93318 36876
rect 93262 36822 93264 36874
rect 93264 36822 93316 36874
rect 93316 36822 93318 36874
rect 93262 36820 93318 36822
rect 93366 36874 93422 36876
rect 93366 36822 93368 36874
rect 93368 36822 93420 36874
rect 93420 36822 93422 36874
rect 93366 36820 93422 36822
rect 93470 36874 93526 36876
rect 93470 36822 93472 36874
rect 93472 36822 93524 36874
rect 93524 36822 93526 36874
rect 93470 36820 93526 36822
rect 130082 36874 130138 36876
rect 130082 36822 130084 36874
rect 130084 36822 130136 36874
rect 130136 36822 130138 36874
rect 130082 36820 130138 36822
rect 130186 36874 130242 36876
rect 130186 36822 130188 36874
rect 130188 36822 130240 36874
rect 130240 36822 130242 36874
rect 130186 36820 130242 36822
rect 130290 36874 130346 36876
rect 130290 36822 130292 36874
rect 130292 36822 130344 36874
rect 130344 36822 130346 36874
rect 130290 36820 130346 36822
rect 144284 36428 144340 36484
rect 141708 36204 141764 36260
rect 38032 36090 38088 36092
rect 38032 36038 38034 36090
rect 38034 36038 38086 36090
rect 38086 36038 38088 36090
rect 38032 36036 38088 36038
rect 38136 36090 38192 36092
rect 38136 36038 38138 36090
rect 38138 36038 38190 36090
rect 38190 36038 38192 36090
rect 38136 36036 38192 36038
rect 38240 36090 38296 36092
rect 38240 36038 38242 36090
rect 38242 36038 38294 36090
rect 38294 36038 38296 36090
rect 38240 36036 38296 36038
rect 74852 36090 74908 36092
rect 74852 36038 74854 36090
rect 74854 36038 74906 36090
rect 74906 36038 74908 36090
rect 74852 36036 74908 36038
rect 74956 36090 75012 36092
rect 74956 36038 74958 36090
rect 74958 36038 75010 36090
rect 75010 36038 75012 36090
rect 74956 36036 75012 36038
rect 75060 36090 75116 36092
rect 75060 36038 75062 36090
rect 75062 36038 75114 36090
rect 75114 36038 75116 36090
rect 75060 36036 75116 36038
rect 111672 36090 111728 36092
rect 111672 36038 111674 36090
rect 111674 36038 111726 36090
rect 111726 36038 111728 36090
rect 111672 36036 111728 36038
rect 111776 36090 111832 36092
rect 111776 36038 111778 36090
rect 111778 36038 111830 36090
rect 111830 36038 111832 36090
rect 111776 36036 111832 36038
rect 111880 36090 111936 36092
rect 111880 36038 111882 36090
rect 111882 36038 111934 36090
rect 111934 36038 111936 36090
rect 111880 36036 111936 36038
rect 19622 35306 19678 35308
rect 19622 35254 19624 35306
rect 19624 35254 19676 35306
rect 19676 35254 19678 35306
rect 19622 35252 19678 35254
rect 19726 35306 19782 35308
rect 19726 35254 19728 35306
rect 19728 35254 19780 35306
rect 19780 35254 19782 35306
rect 19726 35252 19782 35254
rect 19830 35306 19886 35308
rect 19830 35254 19832 35306
rect 19832 35254 19884 35306
rect 19884 35254 19886 35306
rect 19830 35252 19886 35254
rect 56442 35306 56498 35308
rect 56442 35254 56444 35306
rect 56444 35254 56496 35306
rect 56496 35254 56498 35306
rect 56442 35252 56498 35254
rect 56546 35306 56602 35308
rect 56546 35254 56548 35306
rect 56548 35254 56600 35306
rect 56600 35254 56602 35306
rect 56546 35252 56602 35254
rect 56650 35306 56706 35308
rect 56650 35254 56652 35306
rect 56652 35254 56704 35306
rect 56704 35254 56706 35306
rect 56650 35252 56706 35254
rect 93262 35306 93318 35308
rect 93262 35254 93264 35306
rect 93264 35254 93316 35306
rect 93316 35254 93318 35306
rect 93262 35252 93318 35254
rect 93366 35306 93422 35308
rect 93366 35254 93368 35306
rect 93368 35254 93420 35306
rect 93420 35254 93422 35306
rect 93366 35252 93422 35254
rect 93470 35306 93526 35308
rect 93470 35254 93472 35306
rect 93472 35254 93524 35306
rect 93524 35254 93526 35306
rect 93470 35252 93526 35254
rect 130082 35306 130138 35308
rect 130082 35254 130084 35306
rect 130084 35254 130136 35306
rect 130136 35254 130138 35306
rect 130082 35252 130138 35254
rect 130186 35306 130242 35308
rect 130186 35254 130188 35306
rect 130188 35254 130240 35306
rect 130240 35254 130242 35306
rect 130186 35252 130242 35254
rect 130290 35306 130346 35308
rect 130290 35254 130292 35306
rect 130292 35254 130344 35306
rect 130344 35254 130346 35306
rect 130290 35252 130346 35254
rect 38032 34522 38088 34524
rect 38032 34470 38034 34522
rect 38034 34470 38086 34522
rect 38086 34470 38088 34522
rect 38032 34468 38088 34470
rect 38136 34522 38192 34524
rect 38136 34470 38138 34522
rect 38138 34470 38190 34522
rect 38190 34470 38192 34522
rect 38136 34468 38192 34470
rect 38240 34522 38296 34524
rect 38240 34470 38242 34522
rect 38242 34470 38294 34522
rect 38294 34470 38296 34522
rect 38240 34468 38296 34470
rect 74852 34522 74908 34524
rect 74852 34470 74854 34522
rect 74854 34470 74906 34522
rect 74906 34470 74908 34522
rect 74852 34468 74908 34470
rect 74956 34522 75012 34524
rect 74956 34470 74958 34522
rect 74958 34470 75010 34522
rect 75010 34470 75012 34522
rect 74956 34468 75012 34470
rect 75060 34522 75116 34524
rect 75060 34470 75062 34522
rect 75062 34470 75114 34522
rect 75114 34470 75116 34522
rect 75060 34468 75116 34470
rect 111672 34522 111728 34524
rect 111672 34470 111674 34522
rect 111674 34470 111726 34522
rect 111726 34470 111728 34522
rect 111672 34468 111728 34470
rect 111776 34522 111832 34524
rect 111776 34470 111778 34522
rect 111778 34470 111830 34522
rect 111830 34470 111832 34522
rect 111776 34468 111832 34470
rect 111880 34522 111936 34524
rect 111880 34470 111882 34522
rect 111882 34470 111934 34522
rect 111934 34470 111936 34522
rect 111880 34468 111936 34470
rect 139356 33964 139412 34020
rect 19622 33738 19678 33740
rect 19622 33686 19624 33738
rect 19624 33686 19676 33738
rect 19676 33686 19678 33738
rect 19622 33684 19678 33686
rect 19726 33738 19782 33740
rect 19726 33686 19728 33738
rect 19728 33686 19780 33738
rect 19780 33686 19782 33738
rect 19726 33684 19782 33686
rect 19830 33738 19886 33740
rect 19830 33686 19832 33738
rect 19832 33686 19884 33738
rect 19884 33686 19886 33738
rect 19830 33684 19886 33686
rect 56442 33738 56498 33740
rect 56442 33686 56444 33738
rect 56444 33686 56496 33738
rect 56496 33686 56498 33738
rect 56442 33684 56498 33686
rect 56546 33738 56602 33740
rect 56546 33686 56548 33738
rect 56548 33686 56600 33738
rect 56600 33686 56602 33738
rect 56546 33684 56602 33686
rect 56650 33738 56706 33740
rect 56650 33686 56652 33738
rect 56652 33686 56704 33738
rect 56704 33686 56706 33738
rect 56650 33684 56706 33686
rect 93262 33738 93318 33740
rect 93262 33686 93264 33738
rect 93264 33686 93316 33738
rect 93316 33686 93318 33738
rect 93262 33684 93318 33686
rect 93366 33738 93422 33740
rect 93366 33686 93368 33738
rect 93368 33686 93420 33738
rect 93420 33686 93422 33738
rect 93366 33684 93422 33686
rect 93470 33738 93526 33740
rect 93470 33686 93472 33738
rect 93472 33686 93524 33738
rect 93524 33686 93526 33738
rect 93470 33684 93526 33686
rect 130082 33738 130138 33740
rect 130082 33686 130084 33738
rect 130084 33686 130136 33738
rect 130136 33686 130138 33738
rect 130082 33684 130138 33686
rect 130186 33738 130242 33740
rect 130186 33686 130188 33738
rect 130188 33686 130240 33738
rect 130240 33686 130242 33738
rect 130186 33684 130242 33686
rect 130290 33738 130346 33740
rect 130290 33686 130292 33738
rect 130292 33686 130344 33738
rect 130344 33686 130346 33738
rect 130290 33684 130346 33686
rect 134204 33292 134260 33348
rect 38032 32954 38088 32956
rect 38032 32902 38034 32954
rect 38034 32902 38086 32954
rect 38086 32902 38088 32954
rect 38032 32900 38088 32902
rect 38136 32954 38192 32956
rect 38136 32902 38138 32954
rect 38138 32902 38190 32954
rect 38190 32902 38192 32954
rect 38136 32900 38192 32902
rect 38240 32954 38296 32956
rect 38240 32902 38242 32954
rect 38242 32902 38294 32954
rect 38294 32902 38296 32954
rect 38240 32900 38296 32902
rect 74852 32954 74908 32956
rect 74852 32902 74854 32954
rect 74854 32902 74906 32954
rect 74906 32902 74908 32954
rect 74852 32900 74908 32902
rect 74956 32954 75012 32956
rect 74956 32902 74958 32954
rect 74958 32902 75010 32954
rect 75010 32902 75012 32954
rect 74956 32900 75012 32902
rect 75060 32954 75116 32956
rect 75060 32902 75062 32954
rect 75062 32902 75114 32954
rect 75114 32902 75116 32954
rect 75060 32900 75116 32902
rect 111672 32954 111728 32956
rect 111672 32902 111674 32954
rect 111674 32902 111726 32954
rect 111726 32902 111728 32954
rect 111672 32900 111728 32902
rect 111776 32954 111832 32956
rect 111776 32902 111778 32954
rect 111778 32902 111830 32954
rect 111830 32902 111832 32954
rect 111776 32900 111832 32902
rect 111880 32954 111936 32956
rect 111880 32902 111882 32954
rect 111882 32902 111934 32954
rect 111934 32902 111936 32954
rect 111880 32900 111936 32902
rect 19622 32170 19678 32172
rect 19622 32118 19624 32170
rect 19624 32118 19676 32170
rect 19676 32118 19678 32170
rect 19622 32116 19678 32118
rect 19726 32170 19782 32172
rect 19726 32118 19728 32170
rect 19728 32118 19780 32170
rect 19780 32118 19782 32170
rect 19726 32116 19782 32118
rect 19830 32170 19886 32172
rect 19830 32118 19832 32170
rect 19832 32118 19884 32170
rect 19884 32118 19886 32170
rect 19830 32116 19886 32118
rect 56442 32170 56498 32172
rect 56442 32118 56444 32170
rect 56444 32118 56496 32170
rect 56496 32118 56498 32170
rect 56442 32116 56498 32118
rect 56546 32170 56602 32172
rect 56546 32118 56548 32170
rect 56548 32118 56600 32170
rect 56600 32118 56602 32170
rect 56546 32116 56602 32118
rect 56650 32170 56706 32172
rect 56650 32118 56652 32170
rect 56652 32118 56704 32170
rect 56704 32118 56706 32170
rect 56650 32116 56706 32118
rect 93262 32170 93318 32172
rect 93262 32118 93264 32170
rect 93264 32118 93316 32170
rect 93316 32118 93318 32170
rect 93262 32116 93318 32118
rect 93366 32170 93422 32172
rect 93366 32118 93368 32170
rect 93368 32118 93420 32170
rect 93420 32118 93422 32170
rect 93366 32116 93422 32118
rect 93470 32170 93526 32172
rect 93470 32118 93472 32170
rect 93472 32118 93524 32170
rect 93524 32118 93526 32170
rect 93470 32116 93526 32118
rect 130082 32170 130138 32172
rect 130082 32118 130084 32170
rect 130084 32118 130136 32170
rect 130136 32118 130138 32170
rect 130082 32116 130138 32118
rect 130186 32170 130242 32172
rect 130186 32118 130188 32170
rect 130188 32118 130240 32170
rect 130240 32118 130242 32170
rect 130186 32116 130242 32118
rect 130290 32170 130346 32172
rect 130290 32118 130292 32170
rect 130292 32118 130344 32170
rect 130344 32118 130346 32170
rect 130290 32116 130346 32118
rect 38032 31386 38088 31388
rect 38032 31334 38034 31386
rect 38034 31334 38086 31386
rect 38086 31334 38088 31386
rect 38032 31332 38088 31334
rect 38136 31386 38192 31388
rect 38136 31334 38138 31386
rect 38138 31334 38190 31386
rect 38190 31334 38192 31386
rect 38136 31332 38192 31334
rect 38240 31386 38296 31388
rect 38240 31334 38242 31386
rect 38242 31334 38294 31386
rect 38294 31334 38296 31386
rect 38240 31332 38296 31334
rect 74852 31386 74908 31388
rect 74852 31334 74854 31386
rect 74854 31334 74906 31386
rect 74906 31334 74908 31386
rect 74852 31332 74908 31334
rect 74956 31386 75012 31388
rect 74956 31334 74958 31386
rect 74958 31334 75010 31386
rect 75010 31334 75012 31386
rect 74956 31332 75012 31334
rect 75060 31386 75116 31388
rect 75060 31334 75062 31386
rect 75062 31334 75114 31386
rect 75114 31334 75116 31386
rect 75060 31332 75116 31334
rect 111672 31386 111728 31388
rect 111672 31334 111674 31386
rect 111674 31334 111726 31386
rect 111726 31334 111728 31386
rect 111672 31332 111728 31334
rect 111776 31386 111832 31388
rect 111776 31334 111778 31386
rect 111778 31334 111830 31386
rect 111830 31334 111832 31386
rect 111776 31332 111832 31334
rect 111880 31386 111936 31388
rect 111880 31334 111882 31386
rect 111882 31334 111934 31386
rect 111934 31334 111936 31386
rect 111880 31332 111936 31334
rect 131404 30940 131460 30996
rect 19622 30602 19678 30604
rect 19622 30550 19624 30602
rect 19624 30550 19676 30602
rect 19676 30550 19678 30602
rect 19622 30548 19678 30550
rect 19726 30602 19782 30604
rect 19726 30550 19728 30602
rect 19728 30550 19780 30602
rect 19780 30550 19782 30602
rect 19726 30548 19782 30550
rect 19830 30602 19886 30604
rect 19830 30550 19832 30602
rect 19832 30550 19884 30602
rect 19884 30550 19886 30602
rect 19830 30548 19886 30550
rect 56442 30602 56498 30604
rect 56442 30550 56444 30602
rect 56444 30550 56496 30602
rect 56496 30550 56498 30602
rect 56442 30548 56498 30550
rect 56546 30602 56602 30604
rect 56546 30550 56548 30602
rect 56548 30550 56600 30602
rect 56600 30550 56602 30602
rect 56546 30548 56602 30550
rect 56650 30602 56706 30604
rect 56650 30550 56652 30602
rect 56652 30550 56704 30602
rect 56704 30550 56706 30602
rect 56650 30548 56706 30550
rect 93262 30602 93318 30604
rect 93262 30550 93264 30602
rect 93264 30550 93316 30602
rect 93316 30550 93318 30602
rect 93262 30548 93318 30550
rect 93366 30602 93422 30604
rect 93366 30550 93368 30602
rect 93368 30550 93420 30602
rect 93420 30550 93422 30602
rect 93366 30548 93422 30550
rect 93470 30602 93526 30604
rect 93470 30550 93472 30602
rect 93472 30550 93524 30602
rect 93524 30550 93526 30602
rect 93470 30548 93526 30550
rect 130082 30602 130138 30604
rect 130082 30550 130084 30602
rect 130084 30550 130136 30602
rect 130136 30550 130138 30602
rect 130082 30548 130138 30550
rect 130186 30602 130242 30604
rect 130186 30550 130188 30602
rect 130188 30550 130240 30602
rect 130240 30550 130242 30602
rect 130186 30548 130242 30550
rect 130290 30602 130346 30604
rect 130290 30550 130292 30602
rect 130292 30550 130344 30602
rect 130344 30550 130346 30602
rect 130290 30548 130346 30550
rect 38032 29818 38088 29820
rect 38032 29766 38034 29818
rect 38034 29766 38086 29818
rect 38086 29766 38088 29818
rect 38032 29764 38088 29766
rect 38136 29818 38192 29820
rect 38136 29766 38138 29818
rect 38138 29766 38190 29818
rect 38190 29766 38192 29818
rect 38136 29764 38192 29766
rect 38240 29818 38296 29820
rect 38240 29766 38242 29818
rect 38242 29766 38294 29818
rect 38294 29766 38296 29818
rect 38240 29764 38296 29766
rect 74852 29818 74908 29820
rect 74852 29766 74854 29818
rect 74854 29766 74906 29818
rect 74906 29766 74908 29818
rect 74852 29764 74908 29766
rect 74956 29818 75012 29820
rect 74956 29766 74958 29818
rect 74958 29766 75010 29818
rect 75010 29766 75012 29818
rect 74956 29764 75012 29766
rect 75060 29818 75116 29820
rect 75060 29766 75062 29818
rect 75062 29766 75114 29818
rect 75114 29766 75116 29818
rect 75060 29764 75116 29766
rect 111672 29818 111728 29820
rect 111672 29766 111674 29818
rect 111674 29766 111726 29818
rect 111726 29766 111728 29818
rect 111672 29764 111728 29766
rect 111776 29818 111832 29820
rect 111776 29766 111778 29818
rect 111778 29766 111830 29818
rect 111830 29766 111832 29818
rect 111776 29764 111832 29766
rect 111880 29818 111936 29820
rect 111880 29766 111882 29818
rect 111882 29766 111934 29818
rect 111934 29766 111936 29818
rect 111880 29764 111936 29766
rect 128268 29372 128324 29428
rect 19622 29034 19678 29036
rect 19622 28982 19624 29034
rect 19624 28982 19676 29034
rect 19676 28982 19678 29034
rect 19622 28980 19678 28982
rect 19726 29034 19782 29036
rect 19726 28982 19728 29034
rect 19728 28982 19780 29034
rect 19780 28982 19782 29034
rect 19726 28980 19782 28982
rect 19830 29034 19886 29036
rect 19830 28982 19832 29034
rect 19832 28982 19884 29034
rect 19884 28982 19886 29034
rect 19830 28980 19886 28982
rect 56442 29034 56498 29036
rect 56442 28982 56444 29034
rect 56444 28982 56496 29034
rect 56496 28982 56498 29034
rect 56442 28980 56498 28982
rect 56546 29034 56602 29036
rect 56546 28982 56548 29034
rect 56548 28982 56600 29034
rect 56600 28982 56602 29034
rect 56546 28980 56602 28982
rect 56650 29034 56706 29036
rect 56650 28982 56652 29034
rect 56652 28982 56704 29034
rect 56704 28982 56706 29034
rect 56650 28980 56706 28982
rect 93262 29034 93318 29036
rect 93262 28982 93264 29034
rect 93264 28982 93316 29034
rect 93316 28982 93318 29034
rect 93262 28980 93318 28982
rect 93366 29034 93422 29036
rect 93366 28982 93368 29034
rect 93368 28982 93420 29034
rect 93420 28982 93422 29034
rect 93366 28980 93422 28982
rect 93470 29034 93526 29036
rect 93470 28982 93472 29034
rect 93472 28982 93524 29034
rect 93524 28982 93526 29034
rect 93470 28980 93526 28982
rect 38032 28250 38088 28252
rect 38032 28198 38034 28250
rect 38034 28198 38086 28250
rect 38086 28198 38088 28250
rect 38032 28196 38088 28198
rect 38136 28250 38192 28252
rect 38136 28198 38138 28250
rect 38138 28198 38190 28250
rect 38190 28198 38192 28250
rect 38136 28196 38192 28198
rect 38240 28250 38296 28252
rect 38240 28198 38242 28250
rect 38242 28198 38294 28250
rect 38294 28198 38296 28250
rect 38240 28196 38296 28198
rect 74852 28250 74908 28252
rect 74852 28198 74854 28250
rect 74854 28198 74906 28250
rect 74906 28198 74908 28250
rect 74852 28196 74908 28198
rect 74956 28250 75012 28252
rect 74956 28198 74958 28250
rect 74958 28198 75010 28250
rect 75010 28198 75012 28250
rect 74956 28196 75012 28198
rect 75060 28250 75116 28252
rect 75060 28198 75062 28250
rect 75062 28198 75114 28250
rect 75114 28198 75116 28250
rect 75060 28196 75116 28198
rect 111672 28250 111728 28252
rect 111672 28198 111674 28250
rect 111674 28198 111726 28250
rect 111726 28198 111728 28250
rect 111672 28196 111728 28198
rect 111776 28250 111832 28252
rect 111776 28198 111778 28250
rect 111778 28198 111830 28250
rect 111830 28198 111832 28250
rect 111776 28196 111832 28198
rect 111880 28250 111936 28252
rect 111880 28198 111882 28250
rect 111882 28198 111934 28250
rect 111934 28198 111936 28250
rect 111880 28196 111936 28198
rect 126252 27692 126308 27748
rect 19622 27466 19678 27468
rect 19622 27414 19624 27466
rect 19624 27414 19676 27466
rect 19676 27414 19678 27466
rect 19622 27412 19678 27414
rect 19726 27466 19782 27468
rect 19726 27414 19728 27466
rect 19728 27414 19780 27466
rect 19780 27414 19782 27466
rect 19726 27412 19782 27414
rect 19830 27466 19886 27468
rect 19830 27414 19832 27466
rect 19832 27414 19884 27466
rect 19884 27414 19886 27466
rect 19830 27412 19886 27414
rect 56442 27466 56498 27468
rect 56442 27414 56444 27466
rect 56444 27414 56496 27466
rect 56496 27414 56498 27466
rect 56442 27412 56498 27414
rect 56546 27466 56602 27468
rect 56546 27414 56548 27466
rect 56548 27414 56600 27466
rect 56600 27414 56602 27466
rect 56546 27412 56602 27414
rect 56650 27466 56706 27468
rect 56650 27414 56652 27466
rect 56652 27414 56704 27466
rect 56704 27414 56706 27466
rect 56650 27412 56706 27414
rect 93262 27466 93318 27468
rect 93262 27414 93264 27466
rect 93264 27414 93316 27466
rect 93316 27414 93318 27466
rect 93262 27412 93318 27414
rect 93366 27466 93422 27468
rect 93366 27414 93368 27466
rect 93368 27414 93420 27466
rect 93420 27414 93422 27466
rect 93366 27412 93422 27414
rect 93470 27466 93526 27468
rect 93470 27414 93472 27466
rect 93472 27414 93524 27466
rect 93524 27414 93526 27466
rect 93470 27412 93526 27414
rect 38032 26682 38088 26684
rect 38032 26630 38034 26682
rect 38034 26630 38086 26682
rect 38086 26630 38088 26682
rect 38032 26628 38088 26630
rect 38136 26682 38192 26684
rect 38136 26630 38138 26682
rect 38138 26630 38190 26682
rect 38190 26630 38192 26682
rect 38136 26628 38192 26630
rect 38240 26682 38296 26684
rect 38240 26630 38242 26682
rect 38242 26630 38294 26682
rect 38294 26630 38296 26682
rect 38240 26628 38296 26630
rect 74852 26682 74908 26684
rect 74852 26630 74854 26682
rect 74854 26630 74906 26682
rect 74906 26630 74908 26682
rect 74852 26628 74908 26630
rect 74956 26682 75012 26684
rect 74956 26630 74958 26682
rect 74958 26630 75010 26682
rect 75010 26630 75012 26682
rect 74956 26628 75012 26630
rect 75060 26682 75116 26684
rect 75060 26630 75062 26682
rect 75062 26630 75114 26682
rect 75114 26630 75116 26682
rect 75060 26628 75116 26630
rect 111672 26682 111728 26684
rect 111672 26630 111674 26682
rect 111674 26630 111726 26682
rect 111726 26630 111728 26682
rect 111672 26628 111728 26630
rect 111776 26682 111832 26684
rect 111776 26630 111778 26682
rect 111778 26630 111830 26682
rect 111830 26630 111832 26682
rect 111776 26628 111832 26630
rect 111880 26682 111936 26684
rect 111880 26630 111882 26682
rect 111882 26630 111934 26682
rect 111934 26630 111936 26682
rect 111880 26628 111936 26630
rect 19622 25898 19678 25900
rect 19622 25846 19624 25898
rect 19624 25846 19676 25898
rect 19676 25846 19678 25898
rect 19622 25844 19678 25846
rect 19726 25898 19782 25900
rect 19726 25846 19728 25898
rect 19728 25846 19780 25898
rect 19780 25846 19782 25898
rect 19726 25844 19782 25846
rect 19830 25898 19886 25900
rect 19830 25846 19832 25898
rect 19832 25846 19884 25898
rect 19884 25846 19886 25898
rect 19830 25844 19886 25846
rect 56442 25898 56498 25900
rect 56442 25846 56444 25898
rect 56444 25846 56496 25898
rect 56496 25846 56498 25898
rect 56442 25844 56498 25846
rect 56546 25898 56602 25900
rect 56546 25846 56548 25898
rect 56548 25846 56600 25898
rect 56600 25846 56602 25898
rect 56546 25844 56602 25846
rect 56650 25898 56706 25900
rect 56650 25846 56652 25898
rect 56652 25846 56704 25898
rect 56704 25846 56706 25898
rect 56650 25844 56706 25846
rect 93262 25898 93318 25900
rect 93262 25846 93264 25898
rect 93264 25846 93316 25898
rect 93316 25846 93318 25898
rect 93262 25844 93318 25846
rect 93366 25898 93422 25900
rect 93366 25846 93368 25898
rect 93368 25846 93420 25898
rect 93420 25846 93422 25898
rect 93366 25844 93422 25846
rect 93470 25898 93526 25900
rect 93470 25846 93472 25898
rect 93472 25846 93524 25898
rect 93524 25846 93526 25898
rect 93470 25844 93526 25846
rect 123452 25228 123508 25284
rect 38032 25114 38088 25116
rect 38032 25062 38034 25114
rect 38034 25062 38086 25114
rect 38086 25062 38088 25114
rect 38032 25060 38088 25062
rect 38136 25114 38192 25116
rect 38136 25062 38138 25114
rect 38138 25062 38190 25114
rect 38190 25062 38192 25114
rect 38136 25060 38192 25062
rect 38240 25114 38296 25116
rect 38240 25062 38242 25114
rect 38242 25062 38294 25114
rect 38294 25062 38296 25114
rect 38240 25060 38296 25062
rect 74852 25114 74908 25116
rect 74852 25062 74854 25114
rect 74854 25062 74906 25114
rect 74906 25062 74908 25114
rect 74852 25060 74908 25062
rect 74956 25114 75012 25116
rect 74956 25062 74958 25114
rect 74958 25062 75010 25114
rect 75010 25062 75012 25114
rect 74956 25060 75012 25062
rect 75060 25114 75116 25116
rect 75060 25062 75062 25114
rect 75062 25062 75114 25114
rect 75114 25062 75116 25114
rect 75060 25060 75116 25062
rect 111672 25114 111728 25116
rect 111672 25062 111674 25114
rect 111674 25062 111726 25114
rect 111726 25062 111728 25114
rect 111672 25060 111728 25062
rect 111776 25114 111832 25116
rect 111776 25062 111778 25114
rect 111778 25062 111830 25114
rect 111830 25062 111832 25114
rect 111776 25060 111832 25062
rect 111880 25114 111936 25116
rect 111880 25062 111882 25114
rect 111882 25062 111934 25114
rect 111934 25062 111936 25114
rect 111880 25060 111936 25062
rect 19622 24330 19678 24332
rect 19622 24278 19624 24330
rect 19624 24278 19676 24330
rect 19676 24278 19678 24330
rect 19622 24276 19678 24278
rect 19726 24330 19782 24332
rect 19726 24278 19728 24330
rect 19728 24278 19780 24330
rect 19780 24278 19782 24330
rect 19726 24276 19782 24278
rect 19830 24330 19886 24332
rect 19830 24278 19832 24330
rect 19832 24278 19884 24330
rect 19884 24278 19886 24330
rect 19830 24276 19886 24278
rect 56442 24330 56498 24332
rect 56442 24278 56444 24330
rect 56444 24278 56496 24330
rect 56496 24278 56498 24330
rect 56442 24276 56498 24278
rect 56546 24330 56602 24332
rect 56546 24278 56548 24330
rect 56548 24278 56600 24330
rect 56600 24278 56602 24330
rect 56546 24276 56602 24278
rect 56650 24330 56706 24332
rect 56650 24278 56652 24330
rect 56652 24278 56704 24330
rect 56704 24278 56706 24330
rect 56650 24276 56706 24278
rect 93262 24330 93318 24332
rect 93262 24278 93264 24330
rect 93264 24278 93316 24330
rect 93316 24278 93318 24330
rect 93262 24276 93318 24278
rect 93366 24330 93422 24332
rect 93366 24278 93368 24330
rect 93368 24278 93420 24330
rect 93420 24278 93422 24330
rect 93366 24276 93422 24278
rect 93470 24330 93526 24332
rect 93470 24278 93472 24330
rect 93472 24278 93524 24330
rect 93524 24278 93526 24330
rect 93470 24276 93526 24278
rect 38032 23546 38088 23548
rect 38032 23494 38034 23546
rect 38034 23494 38086 23546
rect 38086 23494 38088 23546
rect 38032 23492 38088 23494
rect 38136 23546 38192 23548
rect 38136 23494 38138 23546
rect 38138 23494 38190 23546
rect 38190 23494 38192 23546
rect 38136 23492 38192 23494
rect 38240 23546 38296 23548
rect 38240 23494 38242 23546
rect 38242 23494 38294 23546
rect 38294 23494 38296 23546
rect 38240 23492 38296 23494
rect 74852 23546 74908 23548
rect 74852 23494 74854 23546
rect 74854 23494 74906 23546
rect 74906 23494 74908 23546
rect 74852 23492 74908 23494
rect 74956 23546 75012 23548
rect 74956 23494 74958 23546
rect 74958 23494 75010 23546
rect 75010 23494 75012 23546
rect 74956 23492 75012 23494
rect 75060 23546 75116 23548
rect 75060 23494 75062 23546
rect 75062 23494 75114 23546
rect 75114 23494 75116 23546
rect 75060 23492 75116 23494
rect 111672 23546 111728 23548
rect 111672 23494 111674 23546
rect 111674 23494 111726 23546
rect 111726 23494 111728 23546
rect 111672 23492 111728 23494
rect 111776 23546 111832 23548
rect 111776 23494 111778 23546
rect 111778 23494 111830 23546
rect 111830 23494 111832 23546
rect 111776 23492 111832 23494
rect 111880 23546 111936 23548
rect 111880 23494 111882 23546
rect 111882 23494 111934 23546
rect 111934 23494 111936 23546
rect 111880 23492 111936 23494
rect 121884 23100 121940 23156
rect 19622 22762 19678 22764
rect 19622 22710 19624 22762
rect 19624 22710 19676 22762
rect 19676 22710 19678 22762
rect 19622 22708 19678 22710
rect 19726 22762 19782 22764
rect 19726 22710 19728 22762
rect 19728 22710 19780 22762
rect 19780 22710 19782 22762
rect 19726 22708 19782 22710
rect 19830 22762 19886 22764
rect 19830 22710 19832 22762
rect 19832 22710 19884 22762
rect 19884 22710 19886 22762
rect 19830 22708 19886 22710
rect 56442 22762 56498 22764
rect 56442 22710 56444 22762
rect 56444 22710 56496 22762
rect 56496 22710 56498 22762
rect 56442 22708 56498 22710
rect 56546 22762 56602 22764
rect 56546 22710 56548 22762
rect 56548 22710 56600 22762
rect 56600 22710 56602 22762
rect 56546 22708 56602 22710
rect 56650 22762 56706 22764
rect 56650 22710 56652 22762
rect 56652 22710 56704 22762
rect 56704 22710 56706 22762
rect 56650 22708 56706 22710
rect 93262 22762 93318 22764
rect 93262 22710 93264 22762
rect 93264 22710 93316 22762
rect 93316 22710 93318 22762
rect 93262 22708 93318 22710
rect 93366 22762 93422 22764
rect 93366 22710 93368 22762
rect 93368 22710 93420 22762
rect 93420 22710 93422 22762
rect 93366 22708 93422 22710
rect 93470 22762 93526 22764
rect 93470 22710 93472 22762
rect 93472 22710 93524 22762
rect 93524 22710 93526 22762
rect 93470 22708 93526 22710
rect 115164 22316 115220 22372
rect 38032 21978 38088 21980
rect 38032 21926 38034 21978
rect 38034 21926 38086 21978
rect 38086 21926 38088 21978
rect 38032 21924 38088 21926
rect 38136 21978 38192 21980
rect 38136 21926 38138 21978
rect 38138 21926 38190 21978
rect 38190 21926 38192 21978
rect 38136 21924 38192 21926
rect 38240 21978 38296 21980
rect 38240 21926 38242 21978
rect 38242 21926 38294 21978
rect 38294 21926 38296 21978
rect 38240 21924 38296 21926
rect 74852 21978 74908 21980
rect 74852 21926 74854 21978
rect 74854 21926 74906 21978
rect 74906 21926 74908 21978
rect 74852 21924 74908 21926
rect 74956 21978 75012 21980
rect 74956 21926 74958 21978
rect 74958 21926 75010 21978
rect 75010 21926 75012 21978
rect 74956 21924 75012 21926
rect 75060 21978 75116 21980
rect 75060 21926 75062 21978
rect 75062 21926 75114 21978
rect 75114 21926 75116 21978
rect 75060 21924 75116 21926
rect 111672 21978 111728 21980
rect 111672 21926 111674 21978
rect 111674 21926 111726 21978
rect 111726 21926 111728 21978
rect 111672 21924 111728 21926
rect 111776 21978 111832 21980
rect 111776 21926 111778 21978
rect 111778 21926 111830 21978
rect 111830 21926 111832 21978
rect 111776 21924 111832 21926
rect 111880 21978 111936 21980
rect 111880 21926 111882 21978
rect 111882 21926 111934 21978
rect 111934 21926 111936 21978
rect 111880 21924 111936 21926
rect 19622 21194 19678 21196
rect 19622 21142 19624 21194
rect 19624 21142 19676 21194
rect 19676 21142 19678 21194
rect 19622 21140 19678 21142
rect 19726 21194 19782 21196
rect 19726 21142 19728 21194
rect 19728 21142 19780 21194
rect 19780 21142 19782 21194
rect 19726 21140 19782 21142
rect 19830 21194 19886 21196
rect 19830 21142 19832 21194
rect 19832 21142 19884 21194
rect 19884 21142 19886 21194
rect 19830 21140 19886 21142
rect 56442 21194 56498 21196
rect 56442 21142 56444 21194
rect 56444 21142 56496 21194
rect 56496 21142 56498 21194
rect 56442 21140 56498 21142
rect 56546 21194 56602 21196
rect 56546 21142 56548 21194
rect 56548 21142 56600 21194
rect 56600 21142 56602 21194
rect 56546 21140 56602 21142
rect 56650 21194 56706 21196
rect 56650 21142 56652 21194
rect 56652 21142 56704 21194
rect 56704 21142 56706 21194
rect 56650 21140 56706 21142
rect 93262 21194 93318 21196
rect 93262 21142 93264 21194
rect 93264 21142 93316 21194
rect 93316 21142 93318 21194
rect 93262 21140 93318 21142
rect 93366 21194 93422 21196
rect 93366 21142 93368 21194
rect 93368 21142 93420 21194
rect 93420 21142 93422 21194
rect 93366 21140 93422 21142
rect 93470 21194 93526 21196
rect 93470 21142 93472 21194
rect 93472 21142 93524 21194
rect 93524 21142 93526 21194
rect 93470 21140 93526 21142
rect 114044 20748 114100 20804
rect 38032 20410 38088 20412
rect 38032 20358 38034 20410
rect 38034 20358 38086 20410
rect 38086 20358 38088 20410
rect 38032 20356 38088 20358
rect 38136 20410 38192 20412
rect 38136 20358 38138 20410
rect 38138 20358 38190 20410
rect 38190 20358 38192 20410
rect 38136 20356 38192 20358
rect 38240 20410 38296 20412
rect 38240 20358 38242 20410
rect 38242 20358 38294 20410
rect 38294 20358 38296 20410
rect 38240 20356 38296 20358
rect 74852 20410 74908 20412
rect 74852 20358 74854 20410
rect 74854 20358 74906 20410
rect 74906 20358 74908 20410
rect 74852 20356 74908 20358
rect 74956 20410 75012 20412
rect 74956 20358 74958 20410
rect 74958 20358 75010 20410
rect 75010 20358 75012 20410
rect 74956 20356 75012 20358
rect 75060 20410 75116 20412
rect 75060 20358 75062 20410
rect 75062 20358 75114 20410
rect 75114 20358 75116 20410
rect 75060 20356 75116 20358
rect 111672 20410 111728 20412
rect 111672 20358 111674 20410
rect 111674 20358 111726 20410
rect 111726 20358 111728 20410
rect 111672 20356 111728 20358
rect 111776 20410 111832 20412
rect 111776 20358 111778 20410
rect 111778 20358 111830 20410
rect 111830 20358 111832 20410
rect 111776 20356 111832 20358
rect 111880 20410 111936 20412
rect 111880 20358 111882 20410
rect 111882 20358 111934 20410
rect 111934 20358 111936 20410
rect 111880 20356 111936 20358
rect 19622 19626 19678 19628
rect 19622 19574 19624 19626
rect 19624 19574 19676 19626
rect 19676 19574 19678 19626
rect 19622 19572 19678 19574
rect 19726 19626 19782 19628
rect 19726 19574 19728 19626
rect 19728 19574 19780 19626
rect 19780 19574 19782 19626
rect 19726 19572 19782 19574
rect 19830 19626 19886 19628
rect 19830 19574 19832 19626
rect 19832 19574 19884 19626
rect 19884 19574 19886 19626
rect 19830 19572 19886 19574
rect 56442 19626 56498 19628
rect 56442 19574 56444 19626
rect 56444 19574 56496 19626
rect 56496 19574 56498 19626
rect 56442 19572 56498 19574
rect 56546 19626 56602 19628
rect 56546 19574 56548 19626
rect 56548 19574 56600 19626
rect 56600 19574 56602 19626
rect 56546 19572 56602 19574
rect 56650 19626 56706 19628
rect 56650 19574 56652 19626
rect 56652 19574 56704 19626
rect 56704 19574 56706 19626
rect 56650 19572 56706 19574
rect 93262 19626 93318 19628
rect 93262 19574 93264 19626
rect 93264 19574 93316 19626
rect 93316 19574 93318 19626
rect 93262 19572 93318 19574
rect 93366 19626 93422 19628
rect 93366 19574 93368 19626
rect 93368 19574 93420 19626
rect 93420 19574 93422 19626
rect 93366 19572 93422 19574
rect 93470 19626 93526 19628
rect 93470 19574 93472 19626
rect 93472 19574 93524 19626
rect 93524 19574 93526 19626
rect 93470 19572 93526 19574
rect 110348 19180 110404 19236
rect 38032 18842 38088 18844
rect 38032 18790 38034 18842
rect 38034 18790 38086 18842
rect 38086 18790 38088 18842
rect 38032 18788 38088 18790
rect 38136 18842 38192 18844
rect 38136 18790 38138 18842
rect 38138 18790 38190 18842
rect 38190 18790 38192 18842
rect 38136 18788 38192 18790
rect 38240 18842 38296 18844
rect 38240 18790 38242 18842
rect 38242 18790 38294 18842
rect 38294 18790 38296 18842
rect 38240 18788 38296 18790
rect 74852 18842 74908 18844
rect 74852 18790 74854 18842
rect 74854 18790 74906 18842
rect 74906 18790 74908 18842
rect 74852 18788 74908 18790
rect 74956 18842 75012 18844
rect 74956 18790 74958 18842
rect 74958 18790 75010 18842
rect 75010 18790 75012 18842
rect 74956 18788 75012 18790
rect 75060 18842 75116 18844
rect 75060 18790 75062 18842
rect 75062 18790 75114 18842
rect 75114 18790 75116 18842
rect 75060 18788 75116 18790
rect 106764 18284 106820 18340
rect 19622 18058 19678 18060
rect 19622 18006 19624 18058
rect 19624 18006 19676 18058
rect 19676 18006 19678 18058
rect 19622 18004 19678 18006
rect 19726 18058 19782 18060
rect 19726 18006 19728 18058
rect 19728 18006 19780 18058
rect 19780 18006 19782 18058
rect 19726 18004 19782 18006
rect 19830 18058 19886 18060
rect 19830 18006 19832 18058
rect 19832 18006 19884 18058
rect 19884 18006 19886 18058
rect 19830 18004 19886 18006
rect 56442 18058 56498 18060
rect 56442 18006 56444 18058
rect 56444 18006 56496 18058
rect 56496 18006 56498 18058
rect 56442 18004 56498 18006
rect 56546 18058 56602 18060
rect 56546 18006 56548 18058
rect 56548 18006 56600 18058
rect 56600 18006 56602 18058
rect 56546 18004 56602 18006
rect 56650 18058 56706 18060
rect 56650 18006 56652 18058
rect 56652 18006 56704 18058
rect 56704 18006 56706 18058
rect 56650 18004 56706 18006
rect 93262 18058 93318 18060
rect 93262 18006 93264 18058
rect 93264 18006 93316 18058
rect 93316 18006 93318 18058
rect 93262 18004 93318 18006
rect 93366 18058 93422 18060
rect 93366 18006 93368 18058
rect 93368 18006 93420 18058
rect 93420 18006 93422 18058
rect 93366 18004 93422 18006
rect 93470 18058 93526 18060
rect 93470 18006 93472 18058
rect 93472 18006 93524 18058
rect 93524 18006 93526 18058
rect 93470 18004 93526 18006
rect 38032 17274 38088 17276
rect 38032 17222 38034 17274
rect 38034 17222 38086 17274
rect 38086 17222 38088 17274
rect 38032 17220 38088 17222
rect 38136 17274 38192 17276
rect 38136 17222 38138 17274
rect 38138 17222 38190 17274
rect 38190 17222 38192 17274
rect 38136 17220 38192 17222
rect 38240 17274 38296 17276
rect 38240 17222 38242 17274
rect 38242 17222 38294 17274
rect 38294 17222 38296 17274
rect 38240 17220 38296 17222
rect 74852 17274 74908 17276
rect 74852 17222 74854 17274
rect 74854 17222 74906 17274
rect 74906 17222 74908 17274
rect 74852 17220 74908 17222
rect 74956 17274 75012 17276
rect 74956 17222 74958 17274
rect 74958 17222 75010 17274
rect 75010 17222 75012 17274
rect 74956 17220 75012 17222
rect 75060 17274 75116 17276
rect 75060 17222 75062 17274
rect 75062 17222 75114 17274
rect 75114 17222 75116 17274
rect 75060 17220 75116 17222
rect 19622 16490 19678 16492
rect 19622 16438 19624 16490
rect 19624 16438 19676 16490
rect 19676 16438 19678 16490
rect 19622 16436 19678 16438
rect 19726 16490 19782 16492
rect 19726 16438 19728 16490
rect 19728 16438 19780 16490
rect 19780 16438 19782 16490
rect 19726 16436 19782 16438
rect 19830 16490 19886 16492
rect 19830 16438 19832 16490
rect 19832 16438 19884 16490
rect 19884 16438 19886 16490
rect 19830 16436 19886 16438
rect 56442 16490 56498 16492
rect 56442 16438 56444 16490
rect 56444 16438 56496 16490
rect 56496 16438 56498 16490
rect 56442 16436 56498 16438
rect 56546 16490 56602 16492
rect 56546 16438 56548 16490
rect 56548 16438 56600 16490
rect 56600 16438 56602 16490
rect 56546 16436 56602 16438
rect 56650 16490 56706 16492
rect 56650 16438 56652 16490
rect 56652 16438 56704 16490
rect 56704 16438 56706 16490
rect 56650 16436 56706 16438
rect 93262 16490 93318 16492
rect 93262 16438 93264 16490
rect 93264 16438 93316 16490
rect 93316 16438 93318 16490
rect 93262 16436 93318 16438
rect 93366 16490 93422 16492
rect 93366 16438 93368 16490
rect 93368 16438 93420 16490
rect 93420 16438 93422 16490
rect 93366 16436 93422 16438
rect 93470 16490 93526 16492
rect 93470 16438 93472 16490
rect 93472 16438 93524 16490
rect 93524 16438 93526 16490
rect 93470 16436 93526 16438
rect 38032 15706 38088 15708
rect 38032 15654 38034 15706
rect 38034 15654 38086 15706
rect 38086 15654 38088 15706
rect 38032 15652 38088 15654
rect 38136 15706 38192 15708
rect 38136 15654 38138 15706
rect 38138 15654 38190 15706
rect 38190 15654 38192 15706
rect 38136 15652 38192 15654
rect 38240 15706 38296 15708
rect 38240 15654 38242 15706
rect 38242 15654 38294 15706
rect 38294 15654 38296 15706
rect 38240 15652 38296 15654
rect 74852 15706 74908 15708
rect 74852 15654 74854 15706
rect 74854 15654 74906 15706
rect 74906 15654 74908 15706
rect 74852 15652 74908 15654
rect 74956 15706 75012 15708
rect 74956 15654 74958 15706
rect 74958 15654 75010 15706
rect 75010 15654 75012 15706
rect 74956 15652 75012 15654
rect 75060 15706 75116 15708
rect 75060 15654 75062 15706
rect 75062 15654 75114 15706
rect 75114 15654 75116 15706
rect 75060 15652 75116 15654
rect 101836 15372 101892 15428
rect 19622 14922 19678 14924
rect 19622 14870 19624 14922
rect 19624 14870 19676 14922
rect 19676 14870 19678 14922
rect 19622 14868 19678 14870
rect 19726 14922 19782 14924
rect 19726 14870 19728 14922
rect 19728 14870 19780 14922
rect 19780 14870 19782 14922
rect 19726 14868 19782 14870
rect 19830 14922 19886 14924
rect 19830 14870 19832 14922
rect 19832 14870 19884 14922
rect 19884 14870 19886 14922
rect 19830 14868 19886 14870
rect 56442 14922 56498 14924
rect 56442 14870 56444 14922
rect 56444 14870 56496 14922
rect 56496 14870 56498 14922
rect 56442 14868 56498 14870
rect 56546 14922 56602 14924
rect 56546 14870 56548 14922
rect 56548 14870 56600 14922
rect 56600 14870 56602 14922
rect 56546 14868 56602 14870
rect 56650 14922 56706 14924
rect 56650 14870 56652 14922
rect 56652 14870 56704 14922
rect 56704 14870 56706 14922
rect 56650 14868 56706 14870
rect 93262 14922 93318 14924
rect 93262 14870 93264 14922
rect 93264 14870 93316 14922
rect 93316 14870 93318 14922
rect 93262 14868 93318 14870
rect 93366 14922 93422 14924
rect 93366 14870 93368 14922
rect 93368 14870 93420 14922
rect 93420 14870 93422 14922
rect 93366 14868 93422 14870
rect 93470 14922 93526 14924
rect 93470 14870 93472 14922
rect 93472 14870 93524 14922
rect 93524 14870 93526 14922
rect 93470 14868 93526 14870
rect 100716 14476 100772 14532
rect 38032 14138 38088 14140
rect 38032 14086 38034 14138
rect 38034 14086 38086 14138
rect 38086 14086 38088 14138
rect 38032 14084 38088 14086
rect 38136 14138 38192 14140
rect 38136 14086 38138 14138
rect 38138 14086 38190 14138
rect 38190 14086 38192 14138
rect 38136 14084 38192 14086
rect 38240 14138 38296 14140
rect 38240 14086 38242 14138
rect 38242 14086 38294 14138
rect 38294 14086 38296 14138
rect 38240 14084 38296 14086
rect 74852 14138 74908 14140
rect 74852 14086 74854 14138
rect 74854 14086 74906 14138
rect 74906 14086 74908 14138
rect 74852 14084 74908 14086
rect 74956 14138 75012 14140
rect 74956 14086 74958 14138
rect 74958 14086 75010 14138
rect 75010 14086 75012 14138
rect 74956 14084 75012 14086
rect 75060 14138 75116 14140
rect 75060 14086 75062 14138
rect 75062 14086 75114 14138
rect 75114 14086 75116 14138
rect 75060 14084 75116 14086
rect 19622 13354 19678 13356
rect 19622 13302 19624 13354
rect 19624 13302 19676 13354
rect 19676 13302 19678 13354
rect 19622 13300 19678 13302
rect 19726 13354 19782 13356
rect 19726 13302 19728 13354
rect 19728 13302 19780 13354
rect 19780 13302 19782 13354
rect 19726 13300 19782 13302
rect 19830 13354 19886 13356
rect 19830 13302 19832 13354
rect 19832 13302 19884 13354
rect 19884 13302 19886 13354
rect 19830 13300 19886 13302
rect 56442 13354 56498 13356
rect 56442 13302 56444 13354
rect 56444 13302 56496 13354
rect 56496 13302 56498 13354
rect 56442 13300 56498 13302
rect 56546 13354 56602 13356
rect 56546 13302 56548 13354
rect 56548 13302 56600 13354
rect 56600 13302 56602 13354
rect 56546 13300 56602 13302
rect 56650 13354 56706 13356
rect 56650 13302 56652 13354
rect 56652 13302 56704 13354
rect 56704 13302 56706 13354
rect 56650 13300 56706 13302
rect 93262 13354 93318 13356
rect 93262 13302 93264 13354
rect 93264 13302 93316 13354
rect 93316 13302 93318 13354
rect 93262 13300 93318 13302
rect 93366 13354 93422 13356
rect 93366 13302 93368 13354
rect 93368 13302 93420 13354
rect 93420 13302 93422 13354
rect 93366 13300 93422 13302
rect 93470 13354 93526 13356
rect 93470 13302 93472 13354
rect 93472 13302 93524 13354
rect 93524 13302 93526 13354
rect 93470 13300 93526 13302
rect 99820 12908 99876 12964
rect 38032 12570 38088 12572
rect 38032 12518 38034 12570
rect 38034 12518 38086 12570
rect 38086 12518 38088 12570
rect 38032 12516 38088 12518
rect 38136 12570 38192 12572
rect 38136 12518 38138 12570
rect 38138 12518 38190 12570
rect 38190 12518 38192 12570
rect 38136 12516 38192 12518
rect 38240 12570 38296 12572
rect 38240 12518 38242 12570
rect 38242 12518 38294 12570
rect 38294 12518 38296 12570
rect 38240 12516 38296 12518
rect 74852 12570 74908 12572
rect 74852 12518 74854 12570
rect 74854 12518 74906 12570
rect 74906 12518 74908 12570
rect 74852 12516 74908 12518
rect 74956 12570 75012 12572
rect 74956 12518 74958 12570
rect 74958 12518 75010 12570
rect 75010 12518 75012 12570
rect 74956 12516 75012 12518
rect 75060 12570 75116 12572
rect 75060 12518 75062 12570
rect 75062 12518 75114 12570
rect 75114 12518 75116 12570
rect 75060 12516 75116 12518
rect 19622 11786 19678 11788
rect 19622 11734 19624 11786
rect 19624 11734 19676 11786
rect 19676 11734 19678 11786
rect 19622 11732 19678 11734
rect 19726 11786 19782 11788
rect 19726 11734 19728 11786
rect 19728 11734 19780 11786
rect 19780 11734 19782 11786
rect 19726 11732 19782 11734
rect 19830 11786 19886 11788
rect 19830 11734 19832 11786
rect 19832 11734 19884 11786
rect 19884 11734 19886 11786
rect 19830 11732 19886 11734
rect 56442 11786 56498 11788
rect 56442 11734 56444 11786
rect 56444 11734 56496 11786
rect 56496 11734 56498 11786
rect 56442 11732 56498 11734
rect 56546 11786 56602 11788
rect 56546 11734 56548 11786
rect 56548 11734 56600 11786
rect 56600 11734 56602 11786
rect 56546 11732 56602 11734
rect 56650 11786 56706 11788
rect 56650 11734 56652 11786
rect 56652 11734 56704 11786
rect 56704 11734 56706 11786
rect 56650 11732 56706 11734
rect 93262 11786 93318 11788
rect 93262 11734 93264 11786
rect 93264 11734 93316 11786
rect 93316 11734 93318 11786
rect 93262 11732 93318 11734
rect 93366 11786 93422 11788
rect 93366 11734 93368 11786
rect 93368 11734 93420 11786
rect 93420 11734 93422 11786
rect 93366 11732 93422 11734
rect 93470 11786 93526 11788
rect 93470 11734 93472 11786
rect 93472 11734 93524 11786
rect 93524 11734 93526 11786
rect 93470 11732 93526 11734
rect 98924 11228 98980 11284
rect 38032 11002 38088 11004
rect 38032 10950 38034 11002
rect 38034 10950 38086 11002
rect 38086 10950 38088 11002
rect 38032 10948 38088 10950
rect 38136 11002 38192 11004
rect 38136 10950 38138 11002
rect 38138 10950 38190 11002
rect 38190 10950 38192 11002
rect 38136 10948 38192 10950
rect 38240 11002 38296 11004
rect 38240 10950 38242 11002
rect 38242 10950 38294 11002
rect 38294 10950 38296 11002
rect 38240 10948 38296 10950
rect 74852 11002 74908 11004
rect 74852 10950 74854 11002
rect 74854 10950 74906 11002
rect 74906 10950 74908 11002
rect 74852 10948 74908 10950
rect 74956 11002 75012 11004
rect 74956 10950 74958 11002
rect 74958 10950 75010 11002
rect 75010 10950 75012 11002
rect 74956 10948 75012 10950
rect 75060 11002 75116 11004
rect 75060 10950 75062 11002
rect 75062 10950 75114 11002
rect 75114 10950 75116 11002
rect 75060 10948 75116 10950
rect 59500 10444 59556 10500
rect 42700 10332 42756 10388
rect 19622 10218 19678 10220
rect 19622 10166 19624 10218
rect 19624 10166 19676 10218
rect 19676 10166 19678 10218
rect 19622 10164 19678 10166
rect 19726 10218 19782 10220
rect 19726 10166 19728 10218
rect 19728 10166 19780 10218
rect 19780 10166 19782 10218
rect 19726 10164 19782 10166
rect 19830 10218 19886 10220
rect 19830 10166 19832 10218
rect 19832 10166 19884 10218
rect 19884 10166 19886 10218
rect 19830 10164 19886 10166
rect 38032 9434 38088 9436
rect 38032 9382 38034 9434
rect 38034 9382 38086 9434
rect 38086 9382 38088 9434
rect 38032 9380 38088 9382
rect 38136 9434 38192 9436
rect 38136 9382 38138 9434
rect 38138 9382 38190 9434
rect 38190 9382 38192 9434
rect 38136 9380 38192 9382
rect 38240 9434 38296 9436
rect 38240 9382 38242 9434
rect 38242 9382 38294 9434
rect 38294 9382 38296 9434
rect 38240 9380 38296 9382
rect 41356 8988 41412 9044
rect 15148 8876 15204 8932
rect 13468 7308 13524 7364
rect 11788 5852 11844 5908
rect 10108 5740 10164 5796
rect 9660 5068 9716 5124
rect 8316 4338 8372 4340
rect 8316 4286 8318 4338
rect 8318 4286 8370 4338
rect 8370 4286 8372 4338
rect 8316 4284 8372 4286
rect 8876 4338 8932 4340
rect 8876 4286 8878 4338
rect 8878 4286 8930 4338
rect 8930 4286 8932 4338
rect 8876 4284 8932 4286
rect 9660 4284 9716 4340
rect 11004 4508 11060 4564
rect 6636 4226 6692 4228
rect 6636 4174 6638 4226
rect 6638 4174 6690 4226
rect 6690 4174 6692 4226
rect 6636 4172 6692 4174
rect 5180 3388 5236 3444
rect 6076 3442 6132 3444
rect 6076 3390 6078 3442
rect 6078 3390 6130 3442
rect 6130 3390 6132 3442
rect 6076 3388 6132 3390
rect 8876 3554 8932 3556
rect 8876 3502 8878 3554
rect 8878 3502 8930 3554
rect 8930 3502 8932 3554
rect 8876 3500 8932 3502
rect 9772 3500 9828 3556
rect 11340 4562 11396 4564
rect 11340 4510 11342 4562
rect 11342 4510 11394 4562
rect 11394 4510 11396 4562
rect 11340 4508 11396 4510
rect 11788 4508 11844 4564
rect 13020 4562 13076 4564
rect 13020 4510 13022 4562
rect 13022 4510 13074 4562
rect 13074 4510 13076 4562
rect 13020 4508 13076 4510
rect 13468 4508 13524 4564
rect 17500 8764 17556 8820
rect 16940 4172 16996 4228
rect 16716 3554 16772 3556
rect 16716 3502 16718 3554
rect 16718 3502 16770 3554
rect 16770 3502 16772 3554
rect 16716 3500 16772 3502
rect 15260 3388 15316 3444
rect 15820 3442 15876 3444
rect 15820 3390 15822 3442
rect 15822 3390 15874 3442
rect 15874 3390 15876 3442
rect 15820 3388 15876 3390
rect 19622 8650 19678 8652
rect 19622 8598 19624 8650
rect 19624 8598 19676 8650
rect 19676 8598 19678 8650
rect 19622 8596 19678 8598
rect 19726 8650 19782 8652
rect 19726 8598 19728 8650
rect 19728 8598 19780 8650
rect 19780 8598 19782 8650
rect 19726 8596 19782 8598
rect 19830 8650 19886 8652
rect 19830 8598 19832 8650
rect 19832 8598 19884 8650
rect 19884 8598 19886 8650
rect 19830 8596 19886 8598
rect 38032 7866 38088 7868
rect 38032 7814 38034 7866
rect 38034 7814 38086 7866
rect 38086 7814 38088 7866
rect 38032 7812 38088 7814
rect 38136 7866 38192 7868
rect 38136 7814 38138 7866
rect 38138 7814 38190 7866
rect 38190 7814 38192 7866
rect 38136 7812 38192 7814
rect 38240 7866 38296 7868
rect 38240 7814 38242 7866
rect 38242 7814 38294 7866
rect 38294 7814 38296 7866
rect 38240 7812 38296 7814
rect 39116 7532 39172 7588
rect 21644 7196 21700 7252
rect 19622 7082 19678 7084
rect 19622 7030 19624 7082
rect 19624 7030 19676 7082
rect 19676 7030 19678 7082
rect 19622 7028 19678 7030
rect 19726 7082 19782 7084
rect 19726 7030 19728 7082
rect 19728 7030 19780 7082
rect 19780 7030 19782 7082
rect 19726 7028 19782 7030
rect 19830 7082 19886 7084
rect 19830 7030 19832 7082
rect 19832 7030 19884 7082
rect 19884 7030 19886 7082
rect 19830 7028 19886 7030
rect 19622 5514 19678 5516
rect 19622 5462 19624 5514
rect 19624 5462 19676 5514
rect 19676 5462 19678 5514
rect 19622 5460 19678 5462
rect 19726 5514 19782 5516
rect 19726 5462 19728 5514
rect 19728 5462 19780 5514
rect 19780 5462 19782 5514
rect 19726 5460 19782 5462
rect 19830 5514 19886 5516
rect 19830 5462 19832 5514
rect 19832 5462 19884 5514
rect 19884 5462 19886 5514
rect 19830 5460 19886 5462
rect 18956 4396 19012 4452
rect 19404 4450 19460 4452
rect 19404 4398 19406 4450
rect 19406 4398 19458 4450
rect 19458 4398 19460 4450
rect 19404 4396 19460 4398
rect 17948 4226 18004 4228
rect 17948 4174 17950 4226
rect 17950 4174 18002 4226
rect 18002 4174 18004 4226
rect 17948 4172 18004 4174
rect 19622 3946 19678 3948
rect 19622 3894 19624 3946
rect 19624 3894 19676 3946
rect 19676 3894 19678 3946
rect 19622 3892 19678 3894
rect 19726 3946 19782 3948
rect 19726 3894 19728 3946
rect 19728 3894 19780 3946
rect 19780 3894 19782 3946
rect 19726 3892 19782 3894
rect 19830 3946 19886 3948
rect 19830 3894 19832 3946
rect 19832 3894 19884 3946
rect 19884 3894 19886 3946
rect 19830 3892 19886 3894
rect 17500 3500 17556 3556
rect 20076 3554 20132 3556
rect 20076 3502 20078 3554
rect 20078 3502 20130 3554
rect 20130 3502 20132 3554
rect 20076 3500 20132 3502
rect 20636 3554 20692 3556
rect 20636 3502 20638 3554
rect 20638 3502 20690 3554
rect 20690 3502 20692 3554
rect 20636 3500 20692 3502
rect 22540 6748 22596 6804
rect 35980 6524 36036 6580
rect 30716 5628 30772 5684
rect 21644 3500 21700 3556
rect 18620 3388 18676 3444
rect 19180 3442 19236 3444
rect 19180 3390 19182 3442
rect 19182 3390 19234 3442
rect 19234 3390 19236 3442
rect 19180 3388 19236 3390
rect 20300 3388 20356 3444
rect 21756 3442 21812 3444
rect 21756 3390 21758 3442
rect 21758 3390 21810 3442
rect 21810 3390 21812 3442
rect 21756 3388 21812 3390
rect 22652 3612 22708 3668
rect 22988 3612 23044 3668
rect 24220 1484 24276 1540
rect 25900 3330 25956 3332
rect 25900 3278 25902 3330
rect 25902 3278 25954 3330
rect 25954 3278 25956 3330
rect 25900 3276 25956 3278
rect 28700 3388 28756 3444
rect 27580 2940 27636 2996
rect 29260 3442 29316 3444
rect 29260 3390 29262 3442
rect 29262 3390 29314 3442
rect 29314 3390 29316 3442
rect 29260 3388 29316 3390
rect 29596 2828 29652 2884
rect 32060 4172 32116 4228
rect 32620 4226 32676 4228
rect 32620 4174 32622 4226
rect 32622 4174 32674 4226
rect 32674 4174 32676 4226
rect 32620 4172 32676 4174
rect 30716 3276 30772 3332
rect 30940 2716 30996 2772
rect 32396 2492 32452 2548
rect 34300 2380 34356 2436
rect 38032 6298 38088 6300
rect 38032 6246 38034 6298
rect 38034 6246 38086 6298
rect 38086 6246 38088 6298
rect 38032 6244 38088 6246
rect 38136 6298 38192 6300
rect 38136 6246 38138 6298
rect 38138 6246 38190 6298
rect 38190 6246 38192 6298
rect 38136 6244 38192 6246
rect 38240 6298 38296 6300
rect 38240 6246 38242 6298
rect 38242 6246 38294 6298
rect 38294 6246 38296 6298
rect 38240 6244 38296 6246
rect 38032 4730 38088 4732
rect 38032 4678 38034 4730
rect 38034 4678 38086 4730
rect 38086 4678 38088 4730
rect 38032 4676 38088 4678
rect 38136 4730 38192 4732
rect 38136 4678 38138 4730
rect 38138 4678 38190 4730
rect 38190 4678 38192 4730
rect 38136 4676 38192 4678
rect 38240 4730 38296 4732
rect 38240 4678 38242 4730
rect 38242 4678 38294 4730
rect 38294 4678 38296 4730
rect 38240 4676 38296 4678
rect 37660 3330 37716 3332
rect 37660 3278 37662 3330
rect 37662 3278 37714 3330
rect 37714 3278 37716 3330
rect 37660 3276 37716 3278
rect 38032 3162 38088 3164
rect 38032 3110 38034 3162
rect 38034 3110 38086 3162
rect 38086 3110 38088 3162
rect 38032 3108 38088 3110
rect 38136 3162 38192 3164
rect 38136 3110 38138 3162
rect 38138 3110 38190 3162
rect 38190 3110 38192 3162
rect 38136 3108 38192 3110
rect 38240 3162 38296 3164
rect 38240 3110 38242 3162
rect 38242 3110 38294 3162
rect 38294 3110 38296 3162
rect 38240 3108 38296 3110
rect 40460 3388 40516 3444
rect 39116 3276 39172 3332
rect 39340 3330 39396 3332
rect 39340 3278 39342 3330
rect 39342 3278 39394 3330
rect 39394 3278 39396 3330
rect 39340 3276 39396 3278
rect 41020 3442 41076 3444
rect 41020 3390 41022 3442
rect 41022 3390 41074 3442
rect 41074 3390 41076 3442
rect 41020 3388 41076 3390
rect 42476 4508 42532 4564
rect 42476 3276 42532 3332
rect 56442 10218 56498 10220
rect 56442 10166 56444 10218
rect 56444 10166 56496 10218
rect 56496 10166 56498 10218
rect 56442 10164 56498 10166
rect 56546 10218 56602 10220
rect 56546 10166 56548 10218
rect 56548 10166 56600 10218
rect 56600 10166 56602 10218
rect 56546 10164 56602 10166
rect 56650 10218 56706 10220
rect 56650 10166 56652 10218
rect 56652 10166 56704 10218
rect 56704 10166 56706 10218
rect 56650 10164 56706 10166
rect 56442 8650 56498 8652
rect 56442 8598 56444 8650
rect 56444 8598 56496 8650
rect 56496 8598 56498 8650
rect 56442 8596 56498 8598
rect 56546 8650 56602 8652
rect 56546 8598 56548 8650
rect 56548 8598 56600 8650
rect 56600 8598 56602 8650
rect 56546 8596 56602 8598
rect 56650 8650 56706 8652
rect 56650 8598 56652 8650
rect 56652 8598 56704 8650
rect 56704 8598 56706 8650
rect 56650 8596 56706 8598
rect 53116 8428 53172 8484
rect 51100 7644 51156 7700
rect 43820 4172 43876 4228
rect 44380 4226 44436 4228
rect 44380 4174 44382 4226
rect 44382 4174 44434 4226
rect 44434 4174 44436 4226
rect 44380 4172 44436 4174
rect 44156 1148 44212 1204
rect 46060 1260 46116 1316
rect 47740 812 47796 868
rect 49420 1372 49476 1428
rect 52220 3388 52276 3444
rect 52780 3442 52836 3444
rect 52780 3390 52782 3442
rect 52782 3390 52834 3442
rect 52834 3390 52836 3442
rect 52780 3388 52836 3390
rect 57260 7420 57316 7476
rect 56442 7082 56498 7084
rect 56442 7030 56444 7082
rect 56444 7030 56496 7082
rect 56496 7030 56498 7082
rect 56442 7028 56498 7030
rect 56546 7082 56602 7084
rect 56546 7030 56548 7082
rect 56548 7030 56600 7082
rect 56600 7030 56602 7082
rect 56546 7028 56602 7030
rect 56650 7082 56706 7084
rect 56650 7030 56652 7082
rect 56652 7030 56704 7082
rect 56704 7030 56706 7082
rect 56650 7028 56706 7030
rect 56442 5514 56498 5516
rect 56442 5462 56444 5514
rect 56444 5462 56496 5514
rect 56496 5462 56498 5514
rect 56442 5460 56498 5462
rect 56546 5514 56602 5516
rect 56546 5462 56548 5514
rect 56548 5462 56600 5514
rect 56600 5462 56602 5514
rect 56546 5460 56602 5462
rect 56650 5514 56706 5516
rect 56650 5462 56652 5514
rect 56652 5462 56704 5514
rect 56704 5462 56706 5514
rect 56650 5460 56706 5462
rect 55916 5292 55972 5348
rect 55580 4172 55636 4228
rect 54236 4060 54292 4116
rect 54460 3330 54516 3332
rect 54460 3278 54462 3330
rect 54462 3278 54514 3330
rect 54514 3278 54516 3330
rect 54460 3276 54516 3278
rect 54236 2940 54292 2996
rect 56140 4226 56196 4228
rect 56140 4174 56142 4226
rect 56142 4174 56194 4226
rect 56194 4174 56196 4226
rect 56140 4172 56196 4174
rect 56442 3946 56498 3948
rect 56442 3894 56444 3946
rect 56444 3894 56496 3946
rect 56496 3894 56498 3946
rect 56442 3892 56498 3894
rect 56546 3946 56602 3948
rect 56546 3894 56548 3946
rect 56548 3894 56600 3946
rect 56600 3894 56602 3946
rect 56546 3892 56602 3894
rect 56650 3946 56706 3948
rect 56650 3894 56652 3946
rect 56652 3894 56704 3946
rect 56704 3894 56706 3946
rect 56650 3892 56706 3894
rect 57260 3612 57316 3668
rect 56924 3276 56980 3332
rect 56924 1036 56980 1092
rect 57820 3330 57876 3332
rect 57820 3278 57822 3330
rect 57822 3278 57874 3330
rect 57874 3278 57876 3330
rect 57820 3276 57876 3278
rect 93262 10218 93318 10220
rect 93262 10166 93264 10218
rect 93264 10166 93316 10218
rect 93316 10166 93318 10218
rect 93262 10164 93318 10166
rect 93366 10218 93422 10220
rect 93366 10166 93368 10218
rect 93368 10166 93420 10218
rect 93420 10166 93422 10218
rect 93366 10164 93422 10166
rect 93470 10218 93526 10220
rect 93470 10166 93472 10218
rect 93472 10166 93524 10218
rect 93524 10166 93526 10218
rect 93470 10164 93526 10166
rect 74852 9434 74908 9436
rect 74852 9382 74854 9434
rect 74854 9382 74906 9434
rect 74906 9382 74908 9434
rect 74852 9380 74908 9382
rect 74956 9434 75012 9436
rect 74956 9382 74958 9434
rect 74958 9382 75010 9434
rect 75010 9382 75012 9434
rect 74956 9380 75012 9382
rect 75060 9434 75116 9436
rect 75060 9382 75062 9434
rect 75062 9382 75114 9434
rect 75114 9382 75116 9434
rect 75060 9380 75116 9382
rect 90748 9100 90804 9156
rect 82908 8876 82964 8932
rect 74852 7866 74908 7868
rect 74852 7814 74854 7866
rect 74854 7814 74906 7866
rect 74906 7814 74908 7866
rect 74852 7812 74908 7814
rect 74956 7866 75012 7868
rect 74956 7814 74958 7866
rect 74958 7814 75010 7866
rect 75010 7814 75012 7866
rect 74956 7812 75012 7814
rect 75060 7866 75116 7868
rect 75060 7814 75062 7866
rect 75062 7814 75114 7866
rect 75114 7814 75116 7866
rect 75060 7812 75116 7814
rect 80556 7308 80612 7364
rect 71260 6860 71316 6916
rect 61292 5180 61348 5236
rect 60396 4844 60452 4900
rect 61292 4396 61348 4452
rect 60396 2828 60452 2884
rect 67340 4172 67396 4228
rect 66220 3948 66276 4004
rect 62636 3612 62692 3668
rect 61180 2604 61236 2660
rect 63980 3388 64036 3444
rect 62860 2940 62916 2996
rect 62636 2492 62692 2548
rect 64540 3442 64596 3444
rect 64540 3390 64542 3442
rect 64542 3390 64594 3442
rect 64594 3390 64596 3442
rect 64540 3388 64596 3390
rect 64092 3276 64148 3332
rect 64876 2492 64932 2548
rect 64092 924 64148 980
rect 67900 4226 67956 4228
rect 67900 4174 67902 4226
rect 67902 4174 67954 4226
rect 67954 4174 67956 4226
rect 67900 4172 67956 4174
rect 67676 2044 67732 2100
rect 69580 2156 69636 2212
rect 77644 6636 77700 6692
rect 74852 6298 74908 6300
rect 74852 6246 74854 6298
rect 74854 6246 74906 6298
rect 74906 6246 74908 6298
rect 74852 6244 74908 6246
rect 74956 6298 75012 6300
rect 74956 6246 74958 6298
rect 74958 6246 75010 6298
rect 75010 6246 75012 6298
rect 74956 6244 75012 6246
rect 75060 6298 75116 6300
rect 75060 6246 75062 6298
rect 75062 6246 75114 6298
rect 75114 6246 75116 6298
rect 75060 6244 75116 6246
rect 76076 6188 76132 6244
rect 75180 5068 75236 5124
rect 74852 4730 74908 4732
rect 74852 4678 74854 4730
rect 74854 4678 74906 4730
rect 74906 4678 74908 4730
rect 74852 4676 74908 4678
rect 74956 4730 75012 4732
rect 74956 4678 74958 4730
rect 74958 4678 75010 4730
rect 75010 4678 75012 4730
rect 74956 4676 75012 4678
rect 75060 4730 75116 4732
rect 75060 4678 75062 4730
rect 75062 4678 75114 4730
rect 75114 4678 75116 4730
rect 75060 4676 75116 4678
rect 73948 4450 74004 4452
rect 73948 4398 73950 4450
rect 73950 4398 74002 4450
rect 74002 4398 74004 4450
rect 73948 4396 74004 4398
rect 73388 4284 73444 4340
rect 72492 4172 72548 4228
rect 73276 4226 73332 4228
rect 73276 4174 73278 4226
rect 73278 4174 73330 4226
rect 73330 4174 73332 4226
rect 73276 4172 73332 4174
rect 72828 3724 72884 3780
rect 75852 5122 75908 5124
rect 75852 5070 75854 5122
rect 75854 5070 75906 5122
rect 75906 5070 75908 5122
rect 75852 5068 75908 5070
rect 75516 4956 75572 5012
rect 75292 4450 75348 4452
rect 75292 4398 75294 4450
rect 75294 4398 75346 4450
rect 75346 4398 75348 4450
rect 75292 4396 75348 4398
rect 79660 5852 79716 5908
rect 76076 4396 76132 4452
rect 76972 5068 77028 5124
rect 77644 5068 77700 5124
rect 77868 5740 77924 5796
rect 78204 5068 78260 5124
rect 78540 5122 78596 5124
rect 78540 5070 78542 5122
rect 78542 5070 78594 5122
rect 78594 5070 78596 5122
rect 78540 5068 78596 5070
rect 78876 5068 78932 5124
rect 79436 5122 79492 5124
rect 79436 5070 79438 5122
rect 79438 5070 79490 5122
rect 79490 5070 79492 5122
rect 79436 5068 79492 5070
rect 82236 7308 82292 7364
rect 80892 4732 80948 4788
rect 81340 4732 81396 4788
rect 82124 4732 82180 4788
rect 75740 3388 75796 3444
rect 74852 3162 74908 3164
rect 74852 3110 74854 3162
rect 74854 3110 74906 3162
rect 74906 3110 74908 3162
rect 74852 3108 74908 3110
rect 74956 3162 75012 3164
rect 74956 3110 74958 3162
rect 74958 3110 75010 3162
rect 75010 3110 75012 3162
rect 74956 3108 75012 3110
rect 75060 3162 75116 3164
rect 75060 3110 75062 3162
rect 75062 3110 75114 3162
rect 75114 3110 75116 3162
rect 75060 3108 75116 3110
rect 74620 2828 74676 2884
rect 77196 3442 77252 3444
rect 77196 3390 77198 3442
rect 77198 3390 77250 3442
rect 77250 3390 77252 3442
rect 77196 3388 77252 3390
rect 78764 3388 78820 3444
rect 77420 3276 77476 3332
rect 79996 4450 80052 4452
rect 79996 4398 79998 4450
rect 79998 4398 80050 4450
rect 80050 4398 80052 4450
rect 79996 4396 80052 4398
rect 80444 4450 80500 4452
rect 80444 4398 80446 4450
rect 80446 4398 80498 4450
rect 80498 4398 80500 4450
rect 80444 4396 80500 4398
rect 81340 4450 81396 4452
rect 81340 4398 81342 4450
rect 81342 4398 81394 4450
rect 81394 4398 81396 4450
rect 81340 4396 81396 4398
rect 80780 3500 80836 3556
rect 82124 4396 82180 4452
rect 83916 8764 83972 8820
rect 83244 5122 83300 5124
rect 83244 5070 83246 5122
rect 83246 5070 83298 5122
rect 83298 5070 83300 5122
rect 83244 5068 83300 5070
rect 83580 5068 83636 5124
rect 90524 8764 90580 8820
rect 88956 7420 89012 7476
rect 87276 7196 87332 7252
rect 84476 6300 84532 6356
rect 86940 6300 86996 6356
rect 85372 5964 85428 6020
rect 84588 5068 84644 5124
rect 82684 4732 82740 4788
rect 85372 5068 85428 5124
rect 85596 5180 85652 5236
rect 85932 4844 85988 4900
rect 86380 4898 86436 4900
rect 86380 4846 86382 4898
rect 86382 4846 86434 4898
rect 86434 4846 86436 4898
rect 86380 4844 86436 4846
rect 78876 812 78932 868
rect 79100 3388 79156 3444
rect 82684 3500 82740 3556
rect 81116 3442 81172 3444
rect 81116 3390 81118 3442
rect 81118 3390 81170 3442
rect 81170 3390 81172 3442
rect 81116 3388 81172 3390
rect 82460 3388 82516 3444
rect 85820 4172 85876 4228
rect 83356 3388 83412 3444
rect 84140 3388 84196 3444
rect 84700 3442 84756 3444
rect 84700 3390 84702 3442
rect 84702 3390 84754 3442
rect 84754 3390 84756 3442
rect 84700 3388 84756 3390
rect 86716 4226 86772 4228
rect 86716 4174 86718 4226
rect 86718 4174 86770 4226
rect 86770 4174 86772 4226
rect 86716 4172 86772 4174
rect 88396 7196 88452 7252
rect 87612 5180 87668 5236
rect 88060 5234 88116 5236
rect 88060 5182 88062 5234
rect 88062 5182 88114 5234
rect 88114 5182 88116 5234
rect 88060 5180 88116 5182
rect 89404 5180 89460 5236
rect 87948 4844 88004 4900
rect 89292 4844 89348 4900
rect 90188 5234 90244 5236
rect 90188 5182 90190 5234
rect 90190 5182 90242 5234
rect 90242 5182 90244 5234
rect 90188 5180 90244 5182
rect 89740 4898 89796 4900
rect 89740 4846 89742 4898
rect 89742 4846 89794 4898
rect 89794 4846 89796 4898
rect 89740 4844 89796 4846
rect 93262 8650 93318 8652
rect 93262 8598 93264 8650
rect 93264 8598 93316 8650
rect 93316 8598 93318 8650
rect 93262 8596 93318 8598
rect 93366 8650 93422 8652
rect 93366 8598 93368 8650
rect 93368 8598 93420 8650
rect 93420 8598 93422 8650
rect 93366 8596 93422 8598
rect 93470 8650 93526 8652
rect 93470 8598 93472 8650
rect 93472 8598 93524 8650
rect 93524 8598 93526 8650
rect 93470 8596 93526 8598
rect 93262 7082 93318 7084
rect 93262 7030 93264 7082
rect 93264 7030 93316 7082
rect 93316 7030 93318 7082
rect 93262 7028 93318 7030
rect 93366 7082 93422 7084
rect 93366 7030 93368 7082
rect 93368 7030 93420 7082
rect 93420 7030 93422 7082
rect 93366 7028 93422 7030
rect 93470 7082 93526 7084
rect 93470 7030 93472 7082
rect 93472 7030 93524 7082
rect 93524 7030 93526 7082
rect 93470 7028 93526 7030
rect 97132 5628 97188 5684
rect 93262 5514 93318 5516
rect 93262 5462 93264 5514
rect 93264 5462 93316 5514
rect 93316 5462 93318 5514
rect 93262 5460 93318 5462
rect 93366 5514 93422 5516
rect 93366 5462 93368 5514
rect 93368 5462 93420 5514
rect 93420 5462 93422 5514
rect 93366 5460 93422 5462
rect 93470 5514 93526 5516
rect 93470 5462 93472 5514
rect 93472 5462 93524 5514
rect 93524 5462 93526 5514
rect 93470 5460 93526 5462
rect 90748 5180 90804 5236
rect 90524 4844 90580 4900
rect 90524 4396 90580 4452
rect 87500 3388 87556 3444
rect 88956 3442 89012 3444
rect 88956 3390 88958 3442
rect 88958 3390 89010 3442
rect 89010 3390 89012 3442
rect 88956 3388 89012 3390
rect 89180 3388 89236 3444
rect 91308 4450 91364 4452
rect 91308 4398 91310 4450
rect 91310 4398 91362 4450
rect 91362 4398 91364 4450
rect 91308 4396 91364 4398
rect 93262 3946 93318 3948
rect 93262 3894 93264 3946
rect 93264 3894 93316 3946
rect 93316 3894 93318 3946
rect 93262 3892 93318 3894
rect 93366 3946 93422 3948
rect 93366 3894 93368 3946
rect 93368 3894 93420 3946
rect 93420 3894 93422 3946
rect 93366 3892 93422 3894
rect 93470 3946 93526 3948
rect 93470 3894 93472 3946
rect 93472 3894 93524 3946
rect 93524 3894 93526 3946
rect 93470 3892 93526 3894
rect 92540 3500 92596 3556
rect 93772 3554 93828 3556
rect 93772 3502 93774 3554
rect 93774 3502 93826 3554
rect 93826 3502 93828 3554
rect 93772 3500 93828 3502
rect 90524 3388 90580 3444
rect 90860 3276 90916 3332
rect 92876 3442 92932 3444
rect 92876 3390 92878 3442
rect 92878 3390 92930 3442
rect 92930 3390 92932 3442
rect 92876 3388 92932 3390
rect 94108 2268 94164 2324
rect 97580 4844 97636 4900
rect 97692 4450 97748 4452
rect 97692 4398 97694 4450
rect 97694 4398 97746 4450
rect 97746 4398 97748 4450
rect 97692 4396 97748 4398
rect 98364 4844 98420 4900
rect 96460 3500 96516 3556
rect 95004 3330 95060 3332
rect 95004 3278 95006 3330
rect 95006 3278 95058 3330
rect 95058 3278 95060 3330
rect 95004 3276 95060 3278
rect 95676 2716 95732 2772
rect 95676 1596 95732 1652
rect 97132 3388 97188 3444
rect 98364 4172 98420 4228
rect 97804 3442 97860 3444
rect 97804 3390 97806 3442
rect 97806 3390 97858 3442
rect 97858 3390 97860 3442
rect 97804 3388 97860 3390
rect 98700 4172 98756 4228
rect 99484 11282 99540 11284
rect 99484 11230 99486 11282
rect 99486 11230 99538 11282
rect 99538 11230 99540 11282
rect 99484 11228 99540 11230
rect 99596 10108 99652 10164
rect 99260 5068 99316 5124
rect 98588 3554 98644 3556
rect 98588 3502 98590 3554
rect 98590 3502 98642 3554
rect 98642 3502 98644 3554
rect 98588 3500 98644 3502
rect 99148 3276 99204 3332
rect 98476 1484 98532 1540
rect 99484 5068 99540 5124
rect 100380 5010 100436 5012
rect 100380 4958 100382 5010
rect 100382 4958 100434 5010
rect 100434 4958 100436 5010
rect 100380 4956 100436 4958
rect 100604 4956 100660 5012
rect 99820 4284 99876 4340
rect 100716 4396 100772 4452
rect 100492 4172 100548 4228
rect 99596 4060 99652 4116
rect 99932 4060 99988 4116
rect 105532 14252 105588 14308
rect 102844 12012 102900 12068
rect 102844 10108 102900 10164
rect 101052 4338 101108 4340
rect 101052 4286 101054 4338
rect 101054 4286 101106 4338
rect 101106 4286 101108 4338
rect 101052 4284 101108 4286
rect 103068 5852 103124 5908
rect 102060 5010 102116 5012
rect 102060 4958 102062 5010
rect 102062 4958 102114 5010
rect 102114 4958 102116 5010
rect 102060 4956 102116 4958
rect 102620 5122 102676 5124
rect 102620 5070 102622 5122
rect 102622 5070 102674 5122
rect 102674 5070 102676 5122
rect 102620 5068 102676 5070
rect 103964 5906 104020 5908
rect 103964 5854 103966 5906
rect 103966 5854 104018 5906
rect 104018 5854 104020 5906
rect 103964 5852 104020 5854
rect 103068 5068 103124 5124
rect 102844 4956 102900 5012
rect 102060 4060 102116 4116
rect 101612 1596 101668 1652
rect 102732 4284 102788 4340
rect 103740 5010 103796 5012
rect 103740 4958 103742 5010
rect 103742 4958 103794 5010
rect 103794 4958 103796 5010
rect 103740 4956 103796 4958
rect 103516 4508 103572 4564
rect 102956 4114 103012 4116
rect 102956 4062 102958 4114
rect 102958 4062 103010 4114
rect 103010 4062 103012 4114
rect 102956 4060 103012 4062
rect 105868 10108 105924 10164
rect 105644 6524 105700 6580
rect 104412 5906 104468 5908
rect 104412 5854 104414 5906
rect 104414 5854 104466 5906
rect 104466 5854 104468 5906
rect 104412 5852 104468 5854
rect 104300 5068 104356 5124
rect 104076 3612 104132 3668
rect 102956 3500 103012 3556
rect 104188 4284 104244 4340
rect 104412 3388 104468 3444
rect 105644 4508 105700 4564
rect 108332 15820 108388 15876
rect 109564 10332 109620 10388
rect 108332 5068 108388 5124
rect 109004 7532 109060 7588
rect 106988 4562 107044 4564
rect 106988 4510 106990 4562
rect 106990 4510 107042 4562
rect 107042 4510 107044 4562
rect 106988 4508 107044 4510
rect 109564 5234 109620 5236
rect 109564 5182 109566 5234
rect 109566 5182 109618 5234
rect 109618 5182 109620 5234
rect 109564 5180 109620 5182
rect 105308 4338 105364 4340
rect 105308 4286 105310 4338
rect 105310 4286 105362 4338
rect 105362 4286 105364 4338
rect 105308 4284 105364 4286
rect 104636 3554 104692 3556
rect 104636 3502 104638 3554
rect 104638 3502 104690 3554
rect 104690 3502 104692 3554
rect 104636 3500 104692 3502
rect 106092 3500 106148 3556
rect 105980 3442 106036 3444
rect 105980 3390 105982 3442
rect 105982 3390 106034 3442
rect 106034 3390 106036 3442
rect 105980 3388 106036 3390
rect 102844 2380 102900 2436
rect 106764 3554 106820 3556
rect 106764 3502 106766 3554
rect 106766 3502 106818 3554
rect 106818 3502 106820 3554
rect 106764 3500 106820 3502
rect 108556 4226 108612 4228
rect 108556 4174 108558 4226
rect 108558 4174 108610 4226
rect 108610 4174 108612 4226
rect 108556 4172 108612 4174
rect 107884 3612 107940 3668
rect 108220 3500 108276 3556
rect 107436 3388 107492 3444
rect 107884 3442 107940 3444
rect 107884 3390 107886 3442
rect 107886 3390 107938 3442
rect 107938 3390 107940 3442
rect 107884 3388 107940 3390
rect 108668 3442 108724 3444
rect 108668 3390 108670 3442
rect 108670 3390 108722 3442
rect 108722 3390 108724 3442
rect 108668 3388 108724 3390
rect 109900 4620 109956 4676
rect 109788 4450 109844 4452
rect 109788 4398 109790 4450
rect 109790 4398 109842 4450
rect 109842 4398 109844 4450
rect 109788 4396 109844 4398
rect 109004 3388 109060 3444
rect 109340 4172 109396 4228
rect 109900 3612 109956 3668
rect 110012 4284 110068 4340
rect 109452 3442 109508 3444
rect 109452 3390 109454 3442
rect 109454 3390 109506 3442
rect 109506 3390 109508 3442
rect 109452 3388 109508 3390
rect 111672 18842 111728 18844
rect 111672 18790 111674 18842
rect 111674 18790 111726 18842
rect 111726 18790 111728 18842
rect 111672 18788 111728 18790
rect 111776 18842 111832 18844
rect 111776 18790 111778 18842
rect 111778 18790 111830 18842
rect 111830 18790 111832 18842
rect 111776 18788 111832 18790
rect 111880 18842 111936 18844
rect 111880 18790 111882 18842
rect 111882 18790 111934 18842
rect 111934 18790 111936 18842
rect 111880 18788 111936 18790
rect 111672 17274 111728 17276
rect 111672 17222 111674 17274
rect 111674 17222 111726 17274
rect 111726 17222 111728 17274
rect 111672 17220 111728 17222
rect 111776 17274 111832 17276
rect 111776 17222 111778 17274
rect 111778 17222 111830 17274
rect 111830 17222 111832 17274
rect 111776 17220 111832 17222
rect 111880 17274 111936 17276
rect 111880 17222 111882 17274
rect 111882 17222 111934 17274
rect 111934 17222 111936 17274
rect 111880 17220 111936 17222
rect 111672 15706 111728 15708
rect 111672 15654 111674 15706
rect 111674 15654 111726 15706
rect 111726 15654 111728 15706
rect 111672 15652 111728 15654
rect 111776 15706 111832 15708
rect 111776 15654 111778 15706
rect 111778 15654 111830 15706
rect 111830 15654 111832 15706
rect 111776 15652 111832 15654
rect 111880 15706 111936 15708
rect 111880 15654 111882 15706
rect 111882 15654 111934 15706
rect 111934 15654 111936 15706
rect 111880 15652 111936 15654
rect 111672 14138 111728 14140
rect 111672 14086 111674 14138
rect 111674 14086 111726 14138
rect 111726 14086 111728 14138
rect 111672 14084 111728 14086
rect 111776 14138 111832 14140
rect 111776 14086 111778 14138
rect 111778 14086 111830 14138
rect 111830 14086 111832 14138
rect 111776 14084 111832 14086
rect 111880 14138 111936 14140
rect 111880 14086 111882 14138
rect 111882 14086 111934 14138
rect 111934 14086 111936 14138
rect 111880 14084 111936 14086
rect 111672 12570 111728 12572
rect 111672 12518 111674 12570
rect 111674 12518 111726 12570
rect 111726 12518 111728 12570
rect 111672 12516 111728 12518
rect 111776 12570 111832 12572
rect 111776 12518 111778 12570
rect 111778 12518 111830 12570
rect 111830 12518 111832 12570
rect 111776 12516 111832 12518
rect 111880 12570 111936 12572
rect 111880 12518 111882 12570
rect 111882 12518 111934 12570
rect 111934 12518 111936 12570
rect 111880 12516 111936 12518
rect 111672 11002 111728 11004
rect 111672 10950 111674 11002
rect 111674 10950 111726 11002
rect 111726 10950 111728 11002
rect 111672 10948 111728 10950
rect 111776 11002 111832 11004
rect 111776 10950 111778 11002
rect 111778 10950 111830 11002
rect 111830 10950 111832 11002
rect 111776 10948 111832 10950
rect 111880 11002 111936 11004
rect 111880 10950 111882 11002
rect 111882 10950 111934 11002
rect 111934 10950 111936 11002
rect 111880 10948 111936 10950
rect 111672 9434 111728 9436
rect 111672 9382 111674 9434
rect 111674 9382 111726 9434
rect 111726 9382 111728 9434
rect 111672 9380 111728 9382
rect 111776 9434 111832 9436
rect 111776 9382 111778 9434
rect 111778 9382 111830 9434
rect 111830 9382 111832 9434
rect 111776 9380 111832 9382
rect 111880 9434 111936 9436
rect 111880 9382 111882 9434
rect 111882 9382 111934 9434
rect 111934 9382 111936 9434
rect 111880 9380 111936 9382
rect 112140 9212 112196 9268
rect 110572 8988 110628 9044
rect 111672 7866 111728 7868
rect 111672 7814 111674 7866
rect 111674 7814 111726 7866
rect 111726 7814 111728 7866
rect 111672 7812 111728 7814
rect 111776 7866 111832 7868
rect 111776 7814 111778 7866
rect 111778 7814 111830 7866
rect 111830 7814 111832 7866
rect 111776 7812 111832 7814
rect 111880 7866 111936 7868
rect 111880 7814 111882 7866
rect 111882 7814 111934 7866
rect 111934 7814 111936 7866
rect 111880 7812 111936 7814
rect 111244 5906 111300 5908
rect 111244 5854 111246 5906
rect 111246 5854 111298 5906
rect 111298 5854 111300 5906
rect 111244 5852 111300 5854
rect 111672 6298 111728 6300
rect 111672 6246 111674 6298
rect 111674 6246 111726 6298
rect 111726 6246 111728 6298
rect 111672 6244 111728 6246
rect 111776 6298 111832 6300
rect 111776 6246 111778 6298
rect 111778 6246 111830 6298
rect 111830 6246 111832 6298
rect 111776 6244 111832 6246
rect 111880 6298 111936 6300
rect 111880 6246 111882 6298
rect 111882 6246 111934 6298
rect 111934 6246 111936 6298
rect 111880 6244 111936 6246
rect 111468 5852 111524 5908
rect 110572 4508 110628 4564
rect 110460 4338 110516 4340
rect 110460 4286 110462 4338
rect 110462 4286 110514 4338
rect 110514 4286 110516 4338
rect 110460 4284 110516 4286
rect 111020 5180 111076 5236
rect 111804 5122 111860 5124
rect 111804 5070 111806 5122
rect 111806 5070 111858 5122
rect 111858 5070 111860 5122
rect 111804 5068 111860 5070
rect 110796 4284 110852 4340
rect 111672 4730 111728 4732
rect 111672 4678 111674 4730
rect 111674 4678 111726 4730
rect 111726 4678 111728 4730
rect 111672 4676 111728 4678
rect 111776 4730 111832 4732
rect 111776 4678 111778 4730
rect 111778 4678 111830 4730
rect 111830 4678 111832 4730
rect 111776 4676 111832 4678
rect 111880 4730 111936 4732
rect 111880 4678 111882 4730
rect 111882 4678 111934 4730
rect 111934 4678 111936 4730
rect 111880 4676 111936 4678
rect 112252 5068 112308 5124
rect 112140 5010 112196 5012
rect 112140 4958 112142 5010
rect 112142 4958 112194 5010
rect 112194 4958 112196 5010
rect 112140 4956 112196 4958
rect 112140 4562 112196 4564
rect 112140 4510 112142 4562
rect 112142 4510 112194 4562
rect 112194 4510 112196 4562
rect 112140 4508 112196 4510
rect 111468 4284 111524 4340
rect 111804 4284 111860 4340
rect 110236 3554 110292 3556
rect 110236 3502 110238 3554
rect 110238 3502 110290 3554
rect 110290 3502 110292 3554
rect 110236 3500 110292 3502
rect 111020 3388 111076 3444
rect 111692 3612 111748 3668
rect 112252 3836 112308 3892
rect 112476 4396 112532 4452
rect 113484 7756 113540 7812
rect 114268 6748 114324 6804
rect 112812 5010 112868 5012
rect 112812 4958 112814 5010
rect 112814 4958 112866 5010
rect 112866 4958 112868 5010
rect 112812 4956 112868 4958
rect 113148 5010 113204 5012
rect 113148 4958 113150 5010
rect 113150 4958 113202 5010
rect 113202 4958 113204 5010
rect 113148 4956 113204 4958
rect 112812 3500 112868 3556
rect 111244 3276 111300 3332
rect 111672 3162 111728 3164
rect 111672 3110 111674 3162
rect 111674 3110 111726 3162
rect 111726 3110 111728 3162
rect 111672 3108 111728 3110
rect 111776 3162 111832 3164
rect 111776 3110 111778 3162
rect 111778 3110 111830 3162
rect 111830 3110 111832 3162
rect 111776 3108 111832 3110
rect 111880 3162 111936 3164
rect 111880 3110 111882 3162
rect 111882 3110 111934 3162
rect 111934 3110 111936 3162
rect 111880 3108 111936 3110
rect 112476 2492 112532 2548
rect 112476 1484 112532 1540
rect 113372 3388 113428 3444
rect 113484 3330 113540 3332
rect 113484 3278 113486 3330
rect 113486 3278 113538 3330
rect 113538 3278 113540 3330
rect 113484 3276 113540 3278
rect 113820 3442 113876 3444
rect 113820 3390 113822 3442
rect 113822 3390 113874 3442
rect 113874 3390 113876 3442
rect 113820 3388 113876 3390
rect 113596 2268 113652 2324
rect 114044 5180 114100 5236
rect 114156 4898 114212 4900
rect 114156 4846 114158 4898
rect 114158 4846 114210 4898
rect 114210 4846 114212 4898
rect 114156 4844 114212 4846
rect 114044 3836 114100 3892
rect 114044 3388 114100 3444
rect 118412 21420 118468 21476
rect 116620 16940 116676 16996
rect 115948 11340 116004 11396
rect 116620 10108 116676 10164
rect 119420 19292 119476 19348
rect 119196 17388 119252 17444
rect 119196 14252 119252 14308
rect 118412 9212 118468 9268
rect 115948 7756 116004 7812
rect 118524 6748 118580 6804
rect 117852 5852 117908 5908
rect 115388 5234 115444 5236
rect 115388 5182 115390 5234
rect 115390 5182 115442 5234
rect 115442 5182 115444 5234
rect 115388 5180 115444 5182
rect 115164 4956 115220 5012
rect 115612 4956 115668 5012
rect 114604 4844 114660 4900
rect 115052 3836 115108 3892
rect 115948 5010 116004 5012
rect 115948 4958 115950 5010
rect 115950 4958 116002 5010
rect 116002 4958 116004 5010
rect 115948 4956 116004 4958
rect 114604 3554 114660 3556
rect 114604 3502 114606 3554
rect 114606 3502 114658 3554
rect 114658 3502 114660 3554
rect 114604 3500 114660 3502
rect 115948 3836 116004 3892
rect 116284 5010 116340 5012
rect 116284 4958 116286 5010
rect 116286 4958 116338 5010
rect 116338 4958 116340 5010
rect 116284 4956 116340 4958
rect 117068 4562 117124 4564
rect 117068 4510 117070 4562
rect 117070 4510 117122 4562
rect 117122 4510 117124 4562
rect 117068 4508 117124 4510
rect 116172 3612 116228 3668
rect 116508 3612 116564 3668
rect 113932 3276 113988 3332
rect 112812 1148 112868 1204
rect 114380 3388 114436 3444
rect 115948 1260 116004 1316
rect 116060 3388 116116 3444
rect 116732 3554 116788 3556
rect 116732 3502 116734 3554
rect 116734 3502 116786 3554
rect 116786 3502 116788 3554
rect 116732 3500 116788 3502
rect 117628 5122 117684 5124
rect 117628 5070 117630 5122
rect 117630 5070 117682 5122
rect 117682 5070 117684 5122
rect 117628 5068 117684 5070
rect 117852 5068 117908 5124
rect 118188 4508 118244 4564
rect 117180 3388 117236 3444
rect 117740 3442 117796 3444
rect 117740 3390 117742 3442
rect 117742 3390 117794 3442
rect 117794 3390 117796 3442
rect 117740 3388 117796 3390
rect 118412 3500 118468 3556
rect 117852 1148 117908 1204
rect 120316 11676 120372 11732
rect 121436 7644 121492 7700
rect 119196 3388 119252 3444
rect 119644 4338 119700 4340
rect 119644 4286 119646 4338
rect 119646 4286 119698 4338
rect 119698 4286 119700 4338
rect 119644 4284 119700 4286
rect 120988 4338 121044 4340
rect 120988 4286 120990 4338
rect 120990 4286 121042 4338
rect 121042 4286 121044 4338
rect 120988 4284 121044 4286
rect 120988 3612 121044 3668
rect 119644 3554 119700 3556
rect 119644 3502 119646 3554
rect 119646 3502 119698 3554
rect 119698 3502 119700 3554
rect 119644 3500 119700 3502
rect 119532 3442 119588 3444
rect 119532 3390 119534 3442
rect 119534 3390 119586 3442
rect 119586 3390 119588 3442
rect 119532 3388 119588 3390
rect 120988 2604 121044 2660
rect 123452 11676 123508 11732
rect 125132 23660 125188 23716
rect 124012 10892 124068 10948
rect 123676 8428 123732 8484
rect 121884 4956 121940 5012
rect 122668 4450 122724 4452
rect 122668 4398 122670 4450
rect 122670 4398 122722 4450
rect 122722 4398 122724 4450
rect 122668 4396 122724 4398
rect 121660 4060 121716 4116
rect 119532 1372 119588 1428
rect 122556 3500 122612 3556
rect 122220 3442 122276 3444
rect 122220 3390 122222 3442
rect 122222 3390 122274 3442
rect 122274 3390 122276 3442
rect 122220 3388 122276 3390
rect 122892 4114 122948 4116
rect 122892 4062 122894 4114
rect 122894 4062 122946 4114
rect 122946 4062 122948 4114
rect 122892 4060 122948 4062
rect 122780 3388 122836 3444
rect 123900 5794 123956 5796
rect 123900 5742 123902 5794
rect 123902 5742 123954 5794
rect 123954 5742 123956 5794
rect 123900 5740 123956 5742
rect 125132 6748 125188 6804
rect 125356 7532 125412 7588
rect 124348 5740 124404 5796
rect 123676 3836 123732 3892
rect 124012 4396 124068 4452
rect 124236 3554 124292 3556
rect 124236 3502 124238 3554
rect 124238 3502 124290 3554
rect 124290 3502 124292 3554
rect 124236 3500 124292 3502
rect 125916 5292 125972 5348
rect 124796 4450 124852 4452
rect 124796 4398 124798 4450
rect 124798 4398 124850 4450
rect 124850 4398 124852 4450
rect 124796 4396 124852 4398
rect 127708 10444 127764 10500
rect 127596 8092 127652 8148
rect 130082 29034 130138 29036
rect 130082 28982 130084 29034
rect 130084 28982 130136 29034
rect 130136 28982 130138 29034
rect 130082 28980 130138 28982
rect 130186 29034 130242 29036
rect 130186 28982 130188 29034
rect 130188 28982 130240 29034
rect 130240 28982 130242 29034
rect 130186 28980 130242 28982
rect 130290 29034 130346 29036
rect 130290 28982 130292 29034
rect 130292 28982 130344 29034
rect 130344 28982 130346 29034
rect 130290 28980 130346 28982
rect 130082 27466 130138 27468
rect 130082 27414 130084 27466
rect 130084 27414 130136 27466
rect 130136 27414 130138 27466
rect 130082 27412 130138 27414
rect 130186 27466 130242 27468
rect 130186 27414 130188 27466
rect 130188 27414 130240 27466
rect 130240 27414 130242 27466
rect 130186 27412 130242 27414
rect 130290 27466 130346 27468
rect 130290 27414 130292 27466
rect 130292 27414 130344 27466
rect 130344 27414 130346 27466
rect 130290 27412 130346 27414
rect 130082 25898 130138 25900
rect 130082 25846 130084 25898
rect 130084 25846 130136 25898
rect 130136 25846 130138 25898
rect 130082 25844 130138 25846
rect 130186 25898 130242 25900
rect 130186 25846 130188 25898
rect 130188 25846 130240 25898
rect 130240 25846 130242 25898
rect 130186 25844 130242 25846
rect 130290 25898 130346 25900
rect 130290 25846 130292 25898
rect 130292 25846 130344 25898
rect 130344 25846 130346 25898
rect 130290 25844 130346 25846
rect 130082 24330 130138 24332
rect 130082 24278 130084 24330
rect 130084 24278 130136 24330
rect 130136 24278 130138 24330
rect 130082 24276 130138 24278
rect 130186 24330 130242 24332
rect 130186 24278 130188 24330
rect 130188 24278 130240 24330
rect 130240 24278 130242 24330
rect 130186 24276 130242 24278
rect 130290 24330 130346 24332
rect 130290 24278 130292 24330
rect 130292 24278 130344 24330
rect 130344 24278 130346 24330
rect 130290 24276 130346 24278
rect 130082 22762 130138 22764
rect 130082 22710 130084 22762
rect 130084 22710 130136 22762
rect 130136 22710 130138 22762
rect 130082 22708 130138 22710
rect 130186 22762 130242 22764
rect 130186 22710 130188 22762
rect 130188 22710 130240 22762
rect 130240 22710 130242 22762
rect 130186 22708 130242 22710
rect 130290 22762 130346 22764
rect 130290 22710 130292 22762
rect 130292 22710 130344 22762
rect 130344 22710 130346 22762
rect 130290 22708 130346 22710
rect 130082 21194 130138 21196
rect 130082 21142 130084 21194
rect 130084 21142 130136 21194
rect 130136 21142 130138 21194
rect 130082 21140 130138 21142
rect 130186 21194 130242 21196
rect 130186 21142 130188 21194
rect 130188 21142 130240 21194
rect 130240 21142 130242 21194
rect 130186 21140 130242 21142
rect 130290 21194 130346 21196
rect 130290 21142 130292 21194
rect 130292 21142 130344 21194
rect 130344 21142 130346 21194
rect 130290 21140 130346 21142
rect 130082 19626 130138 19628
rect 130082 19574 130084 19626
rect 130084 19574 130136 19626
rect 130136 19574 130138 19626
rect 130082 19572 130138 19574
rect 130186 19626 130242 19628
rect 130186 19574 130188 19626
rect 130188 19574 130240 19626
rect 130240 19574 130242 19626
rect 130186 19572 130242 19574
rect 130290 19626 130346 19628
rect 130290 19574 130292 19626
rect 130292 19574 130344 19626
rect 130344 19574 130346 19626
rect 130290 19572 130346 19574
rect 130082 18058 130138 18060
rect 130082 18006 130084 18058
rect 130084 18006 130136 18058
rect 130136 18006 130138 18058
rect 130082 18004 130138 18006
rect 130186 18058 130242 18060
rect 130186 18006 130188 18058
rect 130188 18006 130240 18058
rect 130240 18006 130242 18058
rect 130186 18004 130242 18006
rect 130290 18058 130346 18060
rect 130290 18006 130292 18058
rect 130292 18006 130344 18058
rect 130344 18006 130346 18058
rect 130290 18004 130346 18006
rect 130082 16490 130138 16492
rect 130082 16438 130084 16490
rect 130084 16438 130136 16490
rect 130136 16438 130138 16490
rect 130082 16436 130138 16438
rect 130186 16490 130242 16492
rect 130186 16438 130188 16490
rect 130188 16438 130240 16490
rect 130240 16438 130242 16490
rect 130186 16436 130242 16438
rect 130290 16490 130346 16492
rect 130290 16438 130292 16490
rect 130292 16438 130344 16490
rect 130344 16438 130346 16490
rect 130290 16436 130346 16438
rect 130082 14922 130138 14924
rect 130082 14870 130084 14922
rect 130084 14870 130136 14922
rect 130136 14870 130138 14922
rect 130082 14868 130138 14870
rect 130186 14922 130242 14924
rect 130186 14870 130188 14922
rect 130188 14870 130240 14922
rect 130240 14870 130242 14922
rect 130186 14868 130242 14870
rect 130290 14922 130346 14924
rect 130290 14870 130292 14922
rect 130292 14870 130344 14922
rect 130344 14870 130346 14922
rect 130290 14868 130346 14870
rect 130082 13354 130138 13356
rect 130082 13302 130084 13354
rect 130084 13302 130136 13354
rect 130136 13302 130138 13354
rect 130082 13300 130138 13302
rect 130186 13354 130242 13356
rect 130186 13302 130188 13354
rect 130188 13302 130240 13354
rect 130240 13302 130242 13354
rect 130186 13300 130242 13302
rect 130290 13354 130346 13356
rect 130290 13302 130292 13354
rect 130292 13302 130344 13354
rect 130344 13302 130346 13354
rect 130290 13300 130346 13302
rect 130082 11786 130138 11788
rect 130082 11734 130084 11786
rect 130084 11734 130136 11786
rect 130136 11734 130138 11786
rect 130082 11732 130138 11734
rect 130186 11786 130242 11788
rect 130186 11734 130188 11786
rect 130188 11734 130240 11786
rect 130240 11734 130242 11786
rect 130186 11732 130242 11734
rect 130290 11786 130346 11788
rect 130290 11734 130292 11786
rect 130292 11734 130344 11786
rect 130344 11734 130346 11786
rect 130290 11732 130346 11734
rect 130082 10218 130138 10220
rect 130082 10166 130084 10218
rect 130084 10166 130136 10218
rect 130136 10166 130138 10218
rect 130082 10164 130138 10166
rect 130186 10218 130242 10220
rect 130186 10166 130188 10218
rect 130188 10166 130240 10218
rect 130240 10166 130242 10218
rect 130186 10164 130242 10166
rect 130290 10218 130346 10220
rect 130290 10166 130292 10218
rect 130292 10166 130344 10218
rect 130344 10166 130346 10218
rect 130290 10164 130346 10166
rect 130082 8650 130138 8652
rect 130082 8598 130084 8650
rect 130084 8598 130136 8650
rect 130136 8598 130138 8650
rect 130082 8596 130138 8598
rect 130186 8650 130242 8652
rect 130186 8598 130188 8650
rect 130188 8598 130240 8650
rect 130240 8598 130242 8650
rect 130186 8596 130242 8598
rect 130290 8650 130346 8652
rect 130290 8598 130292 8650
rect 130292 8598 130344 8650
rect 130344 8598 130346 8650
rect 130290 8596 130346 8598
rect 127708 6524 127764 6580
rect 127036 5068 127092 5124
rect 126700 4956 126756 5012
rect 124348 1148 124404 1204
rect 124460 3388 124516 3444
rect 126028 3836 126084 3892
rect 127260 4562 127316 4564
rect 127260 4510 127262 4562
rect 127262 4510 127314 4562
rect 127314 4510 127316 4562
rect 127260 4508 127316 4510
rect 130082 7082 130138 7084
rect 130082 7030 130084 7082
rect 130084 7030 130136 7082
rect 130136 7030 130138 7082
rect 130082 7028 130138 7030
rect 130186 7082 130242 7084
rect 130186 7030 130188 7082
rect 130188 7030 130240 7082
rect 130240 7030 130242 7082
rect 130186 7028 130242 7030
rect 130290 7082 130346 7084
rect 130290 7030 130292 7082
rect 130292 7030 130344 7082
rect 130344 7030 130346 7082
rect 130290 7028 130346 7030
rect 129276 6578 129332 6580
rect 129276 6526 129278 6578
rect 129278 6526 129330 6578
rect 129330 6526 129332 6578
rect 129276 6524 129332 6526
rect 129836 6524 129892 6580
rect 127932 4508 127988 4564
rect 126700 4450 126756 4452
rect 126700 4398 126702 4450
rect 126702 4398 126754 4450
rect 126754 4398 126756 4450
rect 126700 4396 126756 4398
rect 126140 3500 126196 3556
rect 125580 3442 125636 3444
rect 125580 3390 125582 3442
rect 125582 3390 125634 3442
rect 125634 3390 125636 3442
rect 125580 3388 125636 3390
rect 127484 3554 127540 3556
rect 127484 3502 127486 3554
rect 127486 3502 127538 3554
rect 127538 3502 127540 3554
rect 127484 3500 127540 3502
rect 128268 3836 128324 3892
rect 128044 3442 128100 3444
rect 128044 3390 128046 3442
rect 128046 3390 128098 3442
rect 128098 3390 128100 3442
rect 128044 3388 128100 3390
rect 129052 5010 129108 5012
rect 129052 4958 129054 5010
rect 129054 4958 129106 5010
rect 129106 4958 129108 5010
rect 129052 4956 129108 4958
rect 129388 4284 129444 4340
rect 128828 3500 128884 3556
rect 129388 3500 129444 3556
rect 128940 924 128996 980
rect 129612 4898 129668 4900
rect 129612 4846 129614 4898
rect 129614 4846 129666 4898
rect 129666 4846 129668 4898
rect 129612 4844 129668 4846
rect 130082 5514 130138 5516
rect 130082 5462 130084 5514
rect 130084 5462 130136 5514
rect 130136 5462 130138 5514
rect 130082 5460 130138 5462
rect 130186 5514 130242 5516
rect 130186 5462 130188 5514
rect 130188 5462 130240 5514
rect 130240 5462 130242 5514
rect 130186 5460 130242 5462
rect 130290 5514 130346 5516
rect 130290 5462 130292 5514
rect 130292 5462 130344 5514
rect 130344 5462 130346 5514
rect 130290 5460 130346 5462
rect 129612 4338 129668 4340
rect 129612 4286 129614 4338
rect 129614 4286 129666 4338
rect 129666 4286 129668 4338
rect 129612 4284 129668 4286
rect 129724 3836 129780 3892
rect 130620 4844 130676 4900
rect 130508 4620 130564 4676
rect 130082 3946 130138 3948
rect 130082 3894 130084 3946
rect 130084 3894 130136 3946
rect 130136 3894 130138 3946
rect 130082 3892 130138 3894
rect 130186 3946 130242 3948
rect 130186 3894 130188 3946
rect 130188 3894 130240 3946
rect 130240 3894 130242 3946
rect 130186 3892 130242 3894
rect 130290 3946 130346 3948
rect 130290 3894 130292 3946
rect 130292 3894 130344 3946
rect 130344 3894 130346 3946
rect 130290 3892 130346 3894
rect 131628 4898 131684 4900
rect 131628 4846 131630 4898
rect 131630 4846 131682 4898
rect 131682 4846 131684 4898
rect 131628 4844 131684 4846
rect 132412 4956 132468 5012
rect 132076 4898 132132 4900
rect 132076 4846 132078 4898
rect 132078 4846 132130 4898
rect 132130 4846 132132 4898
rect 132076 4844 132132 4846
rect 131292 3612 131348 3668
rect 131068 3500 131124 3556
rect 131180 3388 131236 3444
rect 131404 3554 131460 3556
rect 131404 3502 131406 3554
rect 131406 3502 131458 3554
rect 131458 3502 131460 3554
rect 131404 3500 131460 3502
rect 131740 3500 131796 3556
rect 132076 3276 132132 3332
rect 133084 5180 133140 5236
rect 132972 5010 133028 5012
rect 132972 4958 132974 5010
rect 132974 4958 133026 5010
rect 133026 4958 133028 5010
rect 132972 4956 133028 4958
rect 133308 5180 133364 5236
rect 132860 4562 132916 4564
rect 132860 4510 132862 4562
rect 132862 4510 132914 4562
rect 132914 4510 132916 4562
rect 132860 4508 132916 4510
rect 133868 4508 133924 4564
rect 134092 4956 134148 5012
rect 136892 31500 136948 31556
rect 135212 27132 135268 27188
rect 135324 24556 135380 24612
rect 135324 19292 135380 19348
rect 135212 10892 135268 10948
rect 134876 8146 134932 8148
rect 134876 8094 134878 8146
rect 134878 8094 134930 8146
rect 134930 8094 134932 8146
rect 134876 8092 134932 8094
rect 135324 8146 135380 8148
rect 135324 8094 135326 8146
rect 135326 8094 135378 8146
rect 135378 8094 135380 8146
rect 135324 8092 135380 8094
rect 136556 6188 136612 6244
rect 134652 4956 134708 5012
rect 135548 5010 135604 5012
rect 135548 4958 135550 5010
rect 135550 4958 135602 5010
rect 135602 4958 135604 5010
rect 135548 4956 135604 4958
rect 135100 4450 135156 4452
rect 135100 4398 135102 4450
rect 135102 4398 135154 4450
rect 135154 4398 135156 4450
rect 135100 4396 135156 4398
rect 132748 3388 132804 3444
rect 133420 3442 133476 3444
rect 133420 3390 133422 3442
rect 133422 3390 133474 3442
rect 133474 3390 133476 3442
rect 133420 3388 133476 3390
rect 133084 3330 133140 3332
rect 133084 3278 133086 3330
rect 133086 3278 133138 3330
rect 133138 3278 133140 3330
rect 133084 3276 133140 3278
rect 132524 3164 132580 3220
rect 133980 3164 134036 3220
rect 131852 2940 131908 2996
rect 136332 4396 136388 4452
rect 136108 4284 136164 4340
rect 136444 3612 136500 3668
rect 136220 3388 136276 3444
rect 135548 1484 135604 1540
rect 139244 28588 139300 28644
rect 139244 27692 139300 27748
rect 136892 5180 136948 5236
rect 137788 6748 137844 6804
rect 136780 4396 136836 4452
rect 140812 33852 140868 33908
rect 138236 4620 138292 4676
rect 137228 4450 137284 4452
rect 137228 4398 137230 4450
rect 137230 4398 137282 4450
rect 137282 4398 137284 4450
rect 137228 4396 137284 4398
rect 137116 4338 137172 4340
rect 137116 4286 137118 4338
rect 137118 4286 137170 4338
rect 137170 4286 137172 4338
rect 137116 4284 137172 4286
rect 139132 4620 139188 4676
rect 137228 4060 137284 4116
rect 137340 3442 137396 3444
rect 137340 3390 137342 3442
rect 137342 3390 137394 3442
rect 137394 3390 137396 3442
rect 137340 3388 137396 3390
rect 137900 3500 137956 3556
rect 136556 3164 136612 3220
rect 136444 2044 136500 2100
rect 138124 3442 138180 3444
rect 138124 3390 138126 3442
rect 138126 3390 138178 3442
rect 138178 3390 138180 3442
rect 138124 3388 138180 3390
rect 140140 5852 140196 5908
rect 139916 5794 139972 5796
rect 139916 5742 139918 5794
rect 139918 5742 139970 5794
rect 139970 5742 139972 5794
rect 139916 5740 139972 5742
rect 139356 3612 139412 3668
rect 139692 4844 139748 4900
rect 139580 4450 139636 4452
rect 139580 4398 139582 4450
rect 139582 4398 139634 4450
rect 139634 4398 139636 4450
rect 139580 4396 139636 4398
rect 140252 4844 140308 4900
rect 139692 3836 139748 3892
rect 139692 3388 139748 3444
rect 139468 3276 139524 3332
rect 139468 3052 139524 3108
rect 140924 5740 140980 5796
rect 140924 5068 140980 5124
rect 141148 4844 141204 4900
rect 140028 3276 140084 3332
rect 144844 36482 144900 36484
rect 144844 36430 144846 36482
rect 144846 36430 144898 36482
rect 144898 36430 144900 36482
rect 144844 36428 144900 36430
rect 143836 36258 143892 36260
rect 143836 36206 143838 36258
rect 143838 36206 143890 36258
rect 143890 36206 143892 36258
rect 143836 36204 143892 36206
rect 142604 35532 142660 35588
rect 143164 33516 143220 33572
rect 141372 5906 141428 5908
rect 141372 5854 141374 5906
rect 141374 5854 141426 5906
rect 141426 5854 141428 5906
rect 141372 5852 141428 5854
rect 141596 5068 141652 5124
rect 141820 4620 141876 4676
rect 142156 4562 142212 4564
rect 142156 4510 142158 4562
rect 142158 4510 142210 4562
rect 142210 4510 142212 4562
rect 142156 4508 142212 4510
rect 142828 4508 142884 4564
rect 141148 3554 141204 3556
rect 141148 3502 141150 3554
rect 141150 3502 141202 3554
rect 141202 3502 141204 3554
rect 141148 3500 141204 3502
rect 141372 4172 141428 4228
rect 142828 4172 142884 4228
rect 142940 4284 142996 4340
rect 141820 3330 141876 3332
rect 141820 3278 141822 3330
rect 141822 3278 141874 3330
rect 141874 3278 141876 3330
rect 141820 3276 141876 3278
rect 142156 3442 142212 3444
rect 142156 3390 142158 3442
rect 142158 3390 142210 3442
rect 142210 3390 142212 3442
rect 142156 3388 142212 3390
rect 142044 3276 142100 3332
rect 141036 3052 141092 3108
rect 138684 2156 138740 2212
rect 143276 6860 143332 6916
rect 143052 4172 143108 4228
rect 143164 3724 143220 3780
rect 143276 4172 143332 4228
rect 143500 5068 143556 5124
rect 143724 4620 143780 4676
rect 144284 35586 144340 35588
rect 144284 35534 144286 35586
rect 144286 35534 144338 35586
rect 144338 35534 144340 35586
rect 144284 35532 144340 35534
rect 145068 35532 145124 35588
rect 146860 36204 146916 36260
rect 147756 36204 147812 36260
rect 148492 36090 148548 36092
rect 148492 36038 148494 36090
rect 148494 36038 148546 36090
rect 148546 36038 148548 36090
rect 148492 36036 148548 36038
rect 148596 36090 148652 36092
rect 148596 36038 148598 36090
rect 148598 36038 148650 36090
rect 148650 36038 148652 36090
rect 148596 36036 148652 36038
rect 148700 36090 148756 36092
rect 148700 36038 148702 36090
rect 148702 36038 148754 36090
rect 148754 36038 148756 36090
rect 148700 36036 148756 36038
rect 146412 34130 146468 34132
rect 146412 34078 146414 34130
rect 146414 34078 146466 34130
rect 146466 34078 146468 34130
rect 146412 34076 146468 34078
rect 145852 34018 145908 34020
rect 145852 33966 145854 34018
rect 145854 33966 145906 34018
rect 145906 33966 145908 34018
rect 145852 33964 145908 33966
rect 146860 33964 146916 34020
rect 145404 33852 145460 33908
rect 147756 35308 147812 35364
rect 148492 34522 148548 34524
rect 148492 34470 148494 34522
rect 148494 34470 148546 34522
rect 148546 34470 148548 34522
rect 148492 34468 148548 34470
rect 148596 34522 148652 34524
rect 148596 34470 148598 34522
rect 148598 34470 148650 34522
rect 148650 34470 148652 34522
rect 148596 34468 148652 34470
rect 148700 34522 148756 34524
rect 148700 34470 148702 34522
rect 148702 34470 148754 34522
rect 148754 34470 148756 34522
rect 148700 34468 148756 34470
rect 147756 34300 147812 34356
rect 147084 34130 147140 34132
rect 147084 34078 147086 34130
rect 147086 34078 147138 34130
rect 147138 34078 147140 34130
rect 147084 34076 147140 34078
rect 147868 34076 147924 34132
rect 146972 33852 147028 33908
rect 147756 33628 147812 33684
rect 144508 33516 144564 33572
rect 146300 33346 146356 33348
rect 146300 33294 146302 33346
rect 146302 33294 146354 33346
rect 146354 33294 146356 33346
rect 146300 33292 146356 33294
rect 146860 33346 146916 33348
rect 146860 33294 146862 33346
rect 146862 33294 146914 33346
rect 146914 33294 146916 33346
rect 146860 33292 146916 33294
rect 147756 32508 147812 32564
rect 146300 31554 146356 31556
rect 146300 31502 146302 31554
rect 146302 31502 146354 31554
rect 146354 31502 146356 31554
rect 146300 31500 146356 31502
rect 147756 31666 147812 31668
rect 147756 31614 147758 31666
rect 147758 31614 147810 31666
rect 147810 31614 147812 31666
rect 147756 31612 147812 31614
rect 146860 31500 146916 31556
rect 146412 30994 146468 30996
rect 146412 30942 146414 30994
rect 146414 30942 146466 30994
rect 146466 30942 146468 30994
rect 146412 30940 146468 30942
rect 146860 30994 146916 30996
rect 146860 30942 146862 30994
rect 146862 30942 146914 30994
rect 146914 30942 146916 30994
rect 146860 30940 146916 30942
rect 147756 30716 147812 30772
rect 146300 30210 146356 30212
rect 146300 30158 146302 30210
rect 146302 30158 146354 30210
rect 146354 30158 146356 30210
rect 146300 30156 146356 30158
rect 147084 30210 147140 30212
rect 147084 30158 147086 30210
rect 147086 30158 147138 30210
rect 147138 30158 147140 30210
rect 147084 30156 147140 30158
rect 147756 29932 147812 29988
rect 146412 29426 146468 29428
rect 146412 29374 146414 29426
rect 146414 29374 146466 29426
rect 146466 29374 146468 29426
rect 146412 29372 146468 29374
rect 146860 29426 146916 29428
rect 146860 29374 146862 29426
rect 146862 29374 146914 29426
rect 146914 29374 146916 29426
rect 146860 29372 146916 29374
rect 147756 28924 147812 28980
rect 146300 28642 146356 28644
rect 146300 28590 146302 28642
rect 146302 28590 146354 28642
rect 146354 28590 146356 28642
rect 146300 28588 146356 28590
rect 146860 28642 146916 28644
rect 146860 28590 146862 28642
rect 146862 28590 146914 28642
rect 146914 28590 146916 28642
rect 146860 28588 146916 28590
rect 147756 28028 147812 28084
rect 146412 27858 146468 27860
rect 146412 27806 146414 27858
rect 146414 27806 146466 27858
rect 146466 27806 146468 27858
rect 146412 27804 146468 27806
rect 147084 27858 147140 27860
rect 147084 27806 147086 27858
rect 147086 27806 147138 27858
rect 147138 27806 147140 27858
rect 147084 27804 147140 27806
rect 146300 27186 146356 27188
rect 146300 27134 146302 27186
rect 146302 27134 146354 27186
rect 146354 27134 146356 27186
rect 146300 27132 146356 27134
rect 146860 27132 146916 27188
rect 147756 27132 147812 27188
rect 147756 26236 147812 26292
rect 146300 25282 146356 25284
rect 146300 25230 146302 25282
rect 146302 25230 146354 25282
rect 146354 25230 146356 25282
rect 146300 25228 146356 25230
rect 147756 25394 147812 25396
rect 147756 25342 147758 25394
rect 147758 25342 147810 25394
rect 147810 25342 147812 25394
rect 147756 25340 147812 25342
rect 146860 25228 146916 25284
rect 146412 24610 146468 24612
rect 146412 24558 146414 24610
rect 146414 24558 146466 24610
rect 146466 24558 146468 24610
rect 146412 24556 146468 24558
rect 146860 24556 146916 24612
rect 147756 24444 147812 24500
rect 146300 23714 146356 23716
rect 146300 23662 146302 23714
rect 146302 23662 146354 23714
rect 146354 23662 146356 23714
rect 146300 23660 146356 23662
rect 146860 23660 146916 23716
rect 147756 23660 147812 23716
rect 146412 23154 146468 23156
rect 146412 23102 146414 23154
rect 146414 23102 146466 23154
rect 146466 23102 146468 23154
rect 146412 23100 146468 23102
rect 146860 23154 146916 23156
rect 146860 23102 146862 23154
rect 146862 23102 146914 23154
rect 146914 23102 146916 23154
rect 146860 23100 146916 23102
rect 147756 22652 147812 22708
rect 146300 22370 146356 22372
rect 146300 22318 146302 22370
rect 146302 22318 146354 22370
rect 146354 22318 146356 22370
rect 146300 22316 146356 22318
rect 146860 22370 146916 22372
rect 146860 22318 146862 22370
rect 146862 22318 146914 22370
rect 146914 22318 146916 22370
rect 146860 22316 146916 22318
rect 147756 21868 147812 21924
rect 146412 21474 146468 21476
rect 146412 21422 146414 21474
rect 146414 21422 146466 21474
rect 146466 21422 146468 21474
rect 146412 21420 146468 21422
rect 146860 21420 146916 21476
rect 147756 20860 147812 20916
rect 146300 20802 146356 20804
rect 146300 20750 146302 20802
rect 146302 20750 146354 20802
rect 146354 20750 146356 20802
rect 146300 20748 146356 20750
rect 146860 20802 146916 20804
rect 146860 20750 146862 20802
rect 146862 20750 146914 20802
rect 146914 20750 146916 20802
rect 146860 20748 146916 20750
rect 147756 20188 147812 20244
rect 146300 19234 146356 19236
rect 146300 19182 146302 19234
rect 146302 19182 146354 19234
rect 146354 19182 146356 19234
rect 146300 19180 146356 19182
rect 146860 19234 146916 19236
rect 146860 19182 146862 19234
rect 146862 19182 146914 19234
rect 146914 19182 146916 19234
rect 146860 19180 146916 19182
rect 147756 19122 147812 19124
rect 147756 19070 147758 19122
rect 147758 19070 147810 19122
rect 147810 19070 147812 19122
rect 147756 19068 147812 19070
rect 146412 18338 146468 18340
rect 146412 18286 146414 18338
rect 146414 18286 146466 18338
rect 146466 18286 146468 18338
rect 146412 18284 146468 18286
rect 146860 18284 146916 18340
rect 147756 18172 147812 18228
rect 146300 17442 146356 17444
rect 146300 17390 146302 17442
rect 146302 17390 146354 17442
rect 146354 17390 146356 17442
rect 146300 17388 146356 17390
rect 146860 17388 146916 17444
rect 147756 17388 147812 17444
rect 146412 16994 146468 16996
rect 146412 16942 146414 16994
rect 146414 16942 146466 16994
rect 146466 16942 146468 16994
rect 146412 16940 146468 16942
rect 146860 16940 146916 16996
rect 147756 16380 147812 16436
rect 146300 15874 146356 15876
rect 146300 15822 146302 15874
rect 146302 15822 146354 15874
rect 146354 15822 146356 15874
rect 146300 15820 146356 15822
rect 146860 15820 146916 15876
rect 147756 15484 147812 15540
rect 146412 15426 146468 15428
rect 146412 15374 146414 15426
rect 146414 15374 146466 15426
rect 146466 15374 146468 15426
rect 146412 15372 146468 15374
rect 146860 15372 146916 15428
rect 147756 14588 147812 14644
rect 146300 14530 146356 14532
rect 146300 14478 146302 14530
rect 146302 14478 146354 14530
rect 146354 14478 146356 14530
rect 146300 14476 146356 14478
rect 146860 14530 146916 14532
rect 146860 14478 146862 14530
rect 146862 14478 146914 14530
rect 146914 14478 146916 14530
rect 146860 14476 146916 14478
rect 147756 13692 147812 13748
rect 146300 12962 146356 12964
rect 146300 12910 146302 12962
rect 146302 12910 146354 12962
rect 146354 12910 146356 12962
rect 146300 12908 146356 12910
rect 146860 12962 146916 12964
rect 146860 12910 146862 12962
rect 146862 12910 146914 12962
rect 146914 12910 146916 12962
rect 146860 12908 146916 12910
rect 147756 12850 147812 12852
rect 147756 12798 147758 12850
rect 147758 12798 147810 12850
rect 147810 12798 147812 12850
rect 147756 12796 147812 12798
rect 146412 12066 146468 12068
rect 146412 12014 146414 12066
rect 146414 12014 146466 12066
rect 146466 12014 146468 12066
rect 146412 12012 146468 12014
rect 146860 12012 146916 12068
rect 147756 11900 147812 11956
rect 146300 11394 146356 11396
rect 146300 11342 146302 11394
rect 146302 11342 146354 11394
rect 146354 11342 146356 11394
rect 146300 11340 146356 11342
rect 146860 11394 146916 11396
rect 146860 11342 146862 11394
rect 146862 11342 146914 11394
rect 146914 11342 146916 11394
rect 146860 11340 146916 11342
rect 147756 11116 147812 11172
rect 147308 10108 147364 10164
rect 147308 9212 147364 9268
rect 147308 9042 147364 9044
rect 147308 8990 147310 9042
rect 147310 8990 147362 9042
rect 147362 8990 147364 9042
rect 147308 8988 147364 8990
rect 147756 9154 147812 9156
rect 147756 9102 147758 9154
rect 147758 9102 147810 9154
rect 147810 9102 147812 9154
rect 147756 9100 147812 9102
rect 147644 8764 147700 8820
rect 147532 8092 147588 8148
rect 147308 8034 147364 8036
rect 147308 7982 147310 8034
rect 147310 7982 147362 8034
rect 147362 7982 147364 8034
rect 147308 7980 147364 7982
rect 146076 7308 146132 7364
rect 147756 7196 147812 7252
rect 148492 32954 148548 32956
rect 148492 32902 148494 32954
rect 148494 32902 148546 32954
rect 148546 32902 148548 32954
rect 148492 32900 148548 32902
rect 148596 32954 148652 32956
rect 148596 32902 148598 32954
rect 148598 32902 148650 32954
rect 148650 32902 148652 32954
rect 148596 32900 148652 32902
rect 148700 32954 148756 32956
rect 148700 32902 148702 32954
rect 148702 32902 148754 32954
rect 148754 32902 148756 32954
rect 148700 32900 148756 32902
rect 148492 31386 148548 31388
rect 148492 31334 148494 31386
rect 148494 31334 148546 31386
rect 148546 31334 148548 31386
rect 148492 31332 148548 31334
rect 148596 31386 148652 31388
rect 148596 31334 148598 31386
rect 148598 31334 148650 31386
rect 148650 31334 148652 31386
rect 148596 31332 148652 31334
rect 148700 31386 148756 31388
rect 148700 31334 148702 31386
rect 148702 31334 148754 31386
rect 148754 31334 148756 31386
rect 148700 31332 148756 31334
rect 147868 6748 147924 6804
rect 147980 30156 148036 30212
rect 147644 6636 147700 6692
rect 147308 6578 147364 6580
rect 147308 6526 147310 6578
rect 147310 6526 147362 6578
rect 147362 6526 147364 6578
rect 147308 6524 147364 6526
rect 147308 5628 147364 5684
rect 146076 4508 146132 4564
rect 145180 4396 145236 4452
rect 144060 4338 144116 4340
rect 144060 4286 144062 4338
rect 144062 4286 144114 4338
rect 144114 4286 144116 4338
rect 144060 4284 144116 4286
rect 144844 4226 144900 4228
rect 144844 4174 144846 4226
rect 144846 4174 144898 4226
rect 144898 4174 144900 4226
rect 144844 4172 144900 4174
rect 143836 3778 143892 3780
rect 143836 3726 143838 3778
rect 143838 3726 143890 3778
rect 143890 3726 143892 3778
rect 143836 3724 143892 3726
rect 145068 3388 145124 3444
rect 144844 3330 144900 3332
rect 144844 3278 144846 3330
rect 144846 3278 144898 3330
rect 144898 3278 144900 3330
rect 144844 3276 144900 3278
rect 145292 4338 145348 4340
rect 145292 4286 145294 4338
rect 145294 4286 145346 4338
rect 145346 4286 145348 4338
rect 145292 4284 145348 4286
rect 146412 4226 146468 4228
rect 146412 4174 146414 4226
rect 146414 4174 146466 4226
rect 146466 4174 146468 4226
rect 146412 4172 146468 4174
rect 145964 3836 146020 3892
rect 145628 3554 145684 3556
rect 145628 3502 145630 3554
rect 145630 3502 145682 3554
rect 145682 3502 145684 3554
rect 145628 3500 145684 3502
rect 146076 3442 146132 3444
rect 146076 3390 146078 3442
rect 146078 3390 146130 3442
rect 146130 3390 146132 3442
rect 146076 3388 146132 3390
rect 146860 4450 146916 4452
rect 146860 4398 146862 4450
rect 146862 4398 146914 4450
rect 146914 4398 146916 4450
rect 146860 4396 146916 4398
rect 146524 3388 146580 3444
rect 147084 4172 147140 4228
rect 146860 3164 146916 3220
rect 147084 2940 147140 2996
rect 147308 4844 147364 4900
rect 147756 6300 147812 6356
rect 147756 6018 147812 6020
rect 147756 5966 147758 6018
rect 147758 5966 147810 6018
rect 147810 5966 147812 6018
rect 147756 5964 147812 5966
rect 147756 4732 147812 4788
rect 148492 29818 148548 29820
rect 148492 29766 148494 29818
rect 148494 29766 148546 29818
rect 148546 29766 148548 29818
rect 148492 29764 148548 29766
rect 148596 29818 148652 29820
rect 148596 29766 148598 29818
rect 148598 29766 148650 29818
rect 148650 29766 148652 29818
rect 148596 29764 148652 29766
rect 148700 29818 148756 29820
rect 148700 29766 148702 29818
rect 148702 29766 148754 29818
rect 148754 29766 148756 29818
rect 148700 29764 148756 29766
rect 148492 28250 148548 28252
rect 148492 28198 148494 28250
rect 148494 28198 148546 28250
rect 148546 28198 148548 28250
rect 148492 28196 148548 28198
rect 148596 28250 148652 28252
rect 148596 28198 148598 28250
rect 148598 28198 148650 28250
rect 148650 28198 148652 28250
rect 148596 28196 148652 28198
rect 148700 28250 148756 28252
rect 148700 28198 148702 28250
rect 148702 28198 148754 28250
rect 148754 28198 148756 28250
rect 148700 28196 148756 28198
rect 148204 27804 148260 27860
rect 148092 10108 148148 10164
rect 148092 9212 148148 9268
rect 148092 9042 148148 9044
rect 148092 8990 148094 9042
rect 148094 8990 148146 9042
rect 148146 8990 148148 9042
rect 148092 8988 148148 8990
rect 148092 8428 148148 8484
rect 148092 7980 148148 8036
rect 148492 26682 148548 26684
rect 148492 26630 148494 26682
rect 148494 26630 148546 26682
rect 148546 26630 148548 26682
rect 148492 26628 148548 26630
rect 148596 26682 148652 26684
rect 148596 26630 148598 26682
rect 148598 26630 148650 26682
rect 148650 26630 148652 26682
rect 148596 26628 148652 26630
rect 148700 26682 148756 26684
rect 148700 26630 148702 26682
rect 148702 26630 148754 26682
rect 148754 26630 148756 26682
rect 148700 26628 148756 26630
rect 148492 25114 148548 25116
rect 148492 25062 148494 25114
rect 148494 25062 148546 25114
rect 148546 25062 148548 25114
rect 148492 25060 148548 25062
rect 148596 25114 148652 25116
rect 148596 25062 148598 25114
rect 148598 25062 148650 25114
rect 148650 25062 148652 25114
rect 148596 25060 148652 25062
rect 148700 25114 148756 25116
rect 148700 25062 148702 25114
rect 148702 25062 148754 25114
rect 148754 25062 148756 25114
rect 148700 25060 148756 25062
rect 148492 23546 148548 23548
rect 148492 23494 148494 23546
rect 148494 23494 148546 23546
rect 148546 23494 148548 23546
rect 148492 23492 148548 23494
rect 148596 23546 148652 23548
rect 148596 23494 148598 23546
rect 148598 23494 148650 23546
rect 148650 23494 148652 23546
rect 148596 23492 148652 23494
rect 148700 23546 148756 23548
rect 148700 23494 148702 23546
rect 148702 23494 148754 23546
rect 148754 23494 148756 23546
rect 148700 23492 148756 23494
rect 148492 21978 148548 21980
rect 148492 21926 148494 21978
rect 148494 21926 148546 21978
rect 148546 21926 148548 21978
rect 148492 21924 148548 21926
rect 148596 21978 148652 21980
rect 148596 21926 148598 21978
rect 148598 21926 148650 21978
rect 148650 21926 148652 21978
rect 148596 21924 148652 21926
rect 148700 21978 148756 21980
rect 148700 21926 148702 21978
rect 148702 21926 148754 21978
rect 148754 21926 148756 21978
rect 148700 21924 148756 21926
rect 148492 20410 148548 20412
rect 148492 20358 148494 20410
rect 148494 20358 148546 20410
rect 148546 20358 148548 20410
rect 148492 20356 148548 20358
rect 148596 20410 148652 20412
rect 148596 20358 148598 20410
rect 148598 20358 148650 20410
rect 148650 20358 148652 20410
rect 148596 20356 148652 20358
rect 148700 20410 148756 20412
rect 148700 20358 148702 20410
rect 148702 20358 148754 20410
rect 148754 20358 148756 20410
rect 148700 20356 148756 20358
rect 148492 18842 148548 18844
rect 148492 18790 148494 18842
rect 148494 18790 148546 18842
rect 148546 18790 148548 18842
rect 148492 18788 148548 18790
rect 148596 18842 148652 18844
rect 148596 18790 148598 18842
rect 148598 18790 148650 18842
rect 148650 18790 148652 18842
rect 148596 18788 148652 18790
rect 148700 18842 148756 18844
rect 148700 18790 148702 18842
rect 148702 18790 148754 18842
rect 148754 18790 148756 18842
rect 148700 18788 148756 18790
rect 148492 17274 148548 17276
rect 148492 17222 148494 17274
rect 148494 17222 148546 17274
rect 148546 17222 148548 17274
rect 148492 17220 148548 17222
rect 148596 17274 148652 17276
rect 148596 17222 148598 17274
rect 148598 17222 148650 17274
rect 148650 17222 148652 17274
rect 148596 17220 148652 17222
rect 148700 17274 148756 17276
rect 148700 17222 148702 17274
rect 148702 17222 148754 17274
rect 148754 17222 148756 17274
rect 148700 17220 148756 17222
rect 148492 15706 148548 15708
rect 148492 15654 148494 15706
rect 148494 15654 148546 15706
rect 148546 15654 148548 15706
rect 148492 15652 148548 15654
rect 148596 15706 148652 15708
rect 148596 15654 148598 15706
rect 148598 15654 148650 15706
rect 148650 15654 148652 15706
rect 148596 15652 148652 15654
rect 148700 15706 148756 15708
rect 148700 15654 148702 15706
rect 148702 15654 148754 15706
rect 148754 15654 148756 15706
rect 148700 15652 148756 15654
rect 148492 14138 148548 14140
rect 148492 14086 148494 14138
rect 148494 14086 148546 14138
rect 148546 14086 148548 14138
rect 148492 14084 148548 14086
rect 148596 14138 148652 14140
rect 148596 14086 148598 14138
rect 148598 14086 148650 14138
rect 148650 14086 148652 14138
rect 148596 14084 148652 14086
rect 148700 14138 148756 14140
rect 148700 14086 148702 14138
rect 148702 14086 148754 14138
rect 148754 14086 148756 14138
rect 148700 14084 148756 14086
rect 148492 12570 148548 12572
rect 148492 12518 148494 12570
rect 148494 12518 148546 12570
rect 148546 12518 148548 12570
rect 148492 12516 148548 12518
rect 148596 12570 148652 12572
rect 148596 12518 148598 12570
rect 148598 12518 148650 12570
rect 148650 12518 148652 12570
rect 148596 12516 148652 12518
rect 148700 12570 148756 12572
rect 148700 12518 148702 12570
rect 148702 12518 148754 12570
rect 148754 12518 148756 12570
rect 148700 12516 148756 12518
rect 148492 11002 148548 11004
rect 148492 10950 148494 11002
rect 148494 10950 148546 11002
rect 148546 10950 148548 11002
rect 148492 10948 148548 10950
rect 148596 11002 148652 11004
rect 148596 10950 148598 11002
rect 148598 10950 148650 11002
rect 148650 10950 148652 11002
rect 148596 10948 148652 10950
rect 148700 11002 148756 11004
rect 148700 10950 148702 11002
rect 148702 10950 148754 11002
rect 148754 10950 148756 11002
rect 148700 10948 148756 10950
rect 148492 9434 148548 9436
rect 148492 9382 148494 9434
rect 148494 9382 148546 9434
rect 148546 9382 148548 9434
rect 148492 9380 148548 9382
rect 148596 9434 148652 9436
rect 148596 9382 148598 9434
rect 148598 9382 148650 9434
rect 148650 9382 148652 9434
rect 148596 9380 148652 9382
rect 148700 9434 148756 9436
rect 148700 9382 148702 9434
rect 148702 9382 148754 9434
rect 148754 9382 148756 9434
rect 148700 9380 148756 9382
rect 148492 7866 148548 7868
rect 148492 7814 148494 7866
rect 148494 7814 148546 7866
rect 148546 7814 148548 7866
rect 148492 7812 148548 7814
rect 148596 7866 148652 7868
rect 148596 7814 148598 7866
rect 148598 7814 148650 7866
rect 148650 7814 148652 7866
rect 148596 7812 148652 7814
rect 148700 7866 148756 7868
rect 148700 7814 148702 7866
rect 148702 7814 148754 7866
rect 148754 7814 148756 7866
rect 148700 7812 148756 7814
rect 148204 7532 148260 7588
rect 148092 7420 148148 7476
rect 148092 6578 148148 6580
rect 148092 6526 148094 6578
rect 148094 6526 148146 6578
rect 148146 6526 148148 6578
rect 148092 6524 148148 6526
rect 148492 6298 148548 6300
rect 148492 6246 148494 6298
rect 148494 6246 148546 6298
rect 148546 6246 148548 6298
rect 148492 6244 148548 6246
rect 148596 6298 148652 6300
rect 148596 6246 148598 6298
rect 148598 6246 148650 6298
rect 148650 6246 148652 6298
rect 148596 6244 148652 6246
rect 148700 6298 148756 6300
rect 148700 6246 148702 6298
rect 148702 6246 148754 6298
rect 148754 6246 148756 6298
rect 148700 6244 148756 6246
rect 148092 5628 148148 5684
rect 148092 4844 148148 4900
rect 147980 4620 148036 4676
rect 148492 4730 148548 4732
rect 148492 4678 148494 4730
rect 148494 4678 148546 4730
rect 148546 4678 148548 4730
rect 148492 4676 148548 4678
rect 148596 4730 148652 4732
rect 148596 4678 148598 4730
rect 148598 4678 148650 4730
rect 148650 4678 148652 4730
rect 148596 4676 148652 4678
rect 148700 4730 148756 4732
rect 148700 4678 148702 4730
rect 148702 4678 148754 4730
rect 148754 4678 148756 4730
rect 148700 4676 148756 4678
rect 147756 4562 147812 4564
rect 147756 4510 147758 4562
rect 147758 4510 147810 4562
rect 147810 4510 147812 4562
rect 147756 4508 147812 4510
rect 148092 3836 148148 3892
rect 148092 3442 148148 3444
rect 148092 3390 148094 3442
rect 148094 3390 148146 3442
rect 148146 3390 148148 3442
rect 148092 3388 148148 3390
rect 148492 3162 148548 3164
rect 148492 3110 148494 3162
rect 148494 3110 148546 3162
rect 148546 3110 148548 3162
rect 148492 3108 148548 3110
rect 148596 3162 148652 3164
rect 148596 3110 148598 3162
rect 148598 3110 148650 3162
rect 148650 3110 148652 3162
rect 148596 3108 148652 3110
rect 148700 3162 148756 3164
rect 148700 3110 148702 3162
rect 148702 3110 148754 3162
rect 148754 3110 148756 3162
rect 148700 3108 148756 3110
rect 148092 2044 148148 2100
rect 147196 1148 147252 1204
rect 145180 812 145236 868
<< metal3 >>
rect 149200 38836 150000 38864
rect 146066 38780 146076 38836
rect 146132 38780 150000 38836
rect 149200 38752 150000 38780
rect 149200 37940 150000 37968
rect 145954 37884 145964 37940
rect 146020 37884 150000 37940
rect 149200 37856 150000 37884
rect 149200 37044 150000 37072
rect 145842 36988 145852 37044
rect 145908 36988 150000 37044
rect 149200 36960 150000 36988
rect 19612 36820 19622 36876
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19886 36820 19896 36876
rect 56432 36820 56442 36876
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56706 36820 56716 36876
rect 93252 36820 93262 36876
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93526 36820 93536 36876
rect 130072 36820 130082 36876
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130346 36820 130356 36876
rect 144274 36428 144284 36484
rect 144340 36428 144844 36484
rect 144900 36428 144910 36484
rect 141698 36204 141708 36260
rect 141764 36204 143836 36260
rect 143892 36204 146860 36260
rect 146916 36204 146926 36260
rect 147746 36204 147756 36260
rect 147812 36204 148932 36260
rect 148876 36148 148932 36204
rect 149200 36148 150000 36176
rect 148876 36092 150000 36148
rect 38022 36036 38032 36092
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38296 36036 38306 36092
rect 74842 36036 74852 36092
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 75116 36036 75126 36092
rect 111662 36036 111672 36092
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111936 36036 111946 36092
rect 148482 36036 148492 36092
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148756 36036 148766 36092
rect 149200 36064 150000 36092
rect 142594 35532 142604 35588
rect 142660 35532 144284 35588
rect 144340 35532 145068 35588
rect 145124 35532 145134 35588
rect 147746 35308 147756 35364
rect 147812 35308 147822 35364
rect 19612 35252 19622 35308
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19886 35252 19896 35308
rect 56432 35252 56442 35308
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56706 35252 56716 35308
rect 93252 35252 93262 35308
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93526 35252 93536 35308
rect 130072 35252 130082 35308
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130346 35252 130356 35308
rect 147756 35252 147812 35308
rect 149200 35252 150000 35280
rect 147756 35196 150000 35252
rect 149200 35168 150000 35196
rect 38022 34468 38032 34524
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38296 34468 38306 34524
rect 74842 34468 74852 34524
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 75116 34468 75126 34524
rect 111662 34468 111672 34524
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111936 34468 111946 34524
rect 148482 34468 148492 34524
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148756 34468 148766 34524
rect 149200 34356 150000 34384
rect 147746 34300 147756 34356
rect 147812 34300 150000 34356
rect 149200 34272 150000 34300
rect 146402 34076 146412 34132
rect 146468 34076 147084 34132
rect 147140 34076 147868 34132
rect 147924 34076 147934 34132
rect 139346 33964 139356 34020
rect 139412 33964 145852 34020
rect 145908 33964 146860 34020
rect 146916 33964 146926 34020
rect 140802 33852 140812 33908
rect 140868 33852 145404 33908
rect 145460 33852 146972 33908
rect 147028 33852 147038 33908
rect 19612 33684 19622 33740
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19886 33684 19896 33740
rect 56432 33684 56442 33740
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56706 33684 56716 33740
rect 93252 33684 93262 33740
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93526 33684 93536 33740
rect 130072 33684 130082 33740
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130346 33684 130356 33740
rect 147746 33628 147756 33684
rect 147812 33628 147822 33684
rect 147756 33572 147812 33628
rect 143154 33516 143164 33572
rect 143220 33516 144508 33572
rect 144564 33516 144574 33572
rect 147756 33516 147924 33572
rect 147868 33460 147924 33516
rect 149200 33460 150000 33488
rect 147868 33404 150000 33460
rect 149200 33376 150000 33404
rect 134194 33292 134204 33348
rect 134260 33292 146300 33348
rect 146356 33292 146860 33348
rect 146916 33292 146926 33348
rect 38022 32900 38032 32956
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38296 32900 38306 32956
rect 74842 32900 74852 32956
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 75116 32900 75126 32956
rect 111662 32900 111672 32956
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111936 32900 111946 32956
rect 148482 32900 148492 32956
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148756 32900 148766 32956
rect 149200 32564 150000 32592
rect 147746 32508 147756 32564
rect 147812 32508 150000 32564
rect 149200 32480 150000 32508
rect 19612 32116 19622 32172
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19886 32116 19896 32172
rect 56432 32116 56442 32172
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56706 32116 56716 32172
rect 93252 32116 93262 32172
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93526 32116 93536 32172
rect 130072 32116 130082 32172
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130346 32116 130356 32172
rect 149200 31668 150000 31696
rect 147746 31612 147756 31668
rect 147812 31612 150000 31668
rect 149200 31584 150000 31612
rect 136882 31500 136892 31556
rect 136948 31500 146300 31556
rect 146356 31500 146860 31556
rect 146916 31500 146926 31556
rect 38022 31332 38032 31388
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38296 31332 38306 31388
rect 74842 31332 74852 31388
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 75116 31332 75126 31388
rect 111662 31332 111672 31388
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111936 31332 111946 31388
rect 148482 31332 148492 31388
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148756 31332 148766 31388
rect 131394 30940 131404 30996
rect 131460 30940 146412 30996
rect 146468 30940 146860 30996
rect 146916 30940 146926 30996
rect 149200 30772 150000 30800
rect 147746 30716 147756 30772
rect 147812 30716 150000 30772
rect 149200 30688 150000 30716
rect 19612 30548 19622 30604
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19886 30548 19896 30604
rect 56432 30548 56442 30604
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56706 30548 56716 30604
rect 93252 30548 93262 30604
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93526 30548 93536 30604
rect 130072 30548 130082 30604
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130346 30548 130356 30604
rect 146290 30156 146300 30212
rect 146356 30156 147084 30212
rect 147140 30156 147980 30212
rect 148036 30156 148046 30212
rect 147746 29932 147756 29988
rect 147812 29932 148932 29988
rect 148876 29876 148932 29932
rect 149200 29876 150000 29904
rect 148876 29820 150000 29876
rect 38022 29764 38032 29820
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38296 29764 38306 29820
rect 74842 29764 74852 29820
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 75116 29764 75126 29820
rect 111662 29764 111672 29820
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111936 29764 111946 29820
rect 148482 29764 148492 29820
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148756 29764 148766 29820
rect 149200 29792 150000 29820
rect 128258 29372 128268 29428
rect 128324 29372 146412 29428
rect 146468 29372 146860 29428
rect 146916 29372 146926 29428
rect 19612 28980 19622 29036
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19886 28980 19896 29036
rect 56432 28980 56442 29036
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56706 28980 56716 29036
rect 93252 28980 93262 29036
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93526 28980 93536 29036
rect 130072 28980 130082 29036
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130346 28980 130356 29036
rect 149200 28980 150000 29008
rect 147746 28924 147756 28980
rect 147812 28924 150000 28980
rect 149200 28896 150000 28924
rect 139234 28588 139244 28644
rect 139300 28588 146300 28644
rect 146356 28588 146860 28644
rect 146916 28588 146926 28644
rect 38022 28196 38032 28252
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38296 28196 38306 28252
rect 74842 28196 74852 28252
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 75116 28196 75126 28252
rect 111662 28196 111672 28252
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111936 28196 111946 28252
rect 148482 28196 148492 28252
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148756 28196 148766 28252
rect 149200 28084 150000 28112
rect 147746 28028 147756 28084
rect 147812 28028 150000 28084
rect 149200 28000 150000 28028
rect 146402 27804 146412 27860
rect 146468 27804 147084 27860
rect 147140 27804 148204 27860
rect 148260 27804 148270 27860
rect 126242 27692 126252 27748
rect 126308 27692 139244 27748
rect 139300 27692 139310 27748
rect 19612 27412 19622 27468
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19886 27412 19896 27468
rect 56432 27412 56442 27468
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56706 27412 56716 27468
rect 93252 27412 93262 27468
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93526 27412 93536 27468
rect 130072 27412 130082 27468
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130346 27412 130356 27468
rect 149200 27188 150000 27216
rect 135202 27132 135212 27188
rect 135268 27132 146300 27188
rect 146356 27132 146860 27188
rect 146916 27132 146926 27188
rect 147746 27132 147756 27188
rect 147812 27132 150000 27188
rect 149200 27104 150000 27132
rect 38022 26628 38032 26684
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38296 26628 38306 26684
rect 74842 26628 74852 26684
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 75116 26628 75126 26684
rect 111662 26628 111672 26684
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111936 26628 111946 26684
rect 148482 26628 148492 26684
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148756 26628 148766 26684
rect 149200 26292 150000 26320
rect 147746 26236 147756 26292
rect 147812 26236 150000 26292
rect 149200 26208 150000 26236
rect 19612 25844 19622 25900
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19886 25844 19896 25900
rect 56432 25844 56442 25900
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56706 25844 56716 25900
rect 93252 25844 93262 25900
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93526 25844 93536 25900
rect 130072 25844 130082 25900
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130346 25844 130356 25900
rect 149200 25396 150000 25424
rect 147746 25340 147756 25396
rect 147812 25340 150000 25396
rect 149200 25312 150000 25340
rect 123442 25228 123452 25284
rect 123508 25228 146300 25284
rect 146356 25228 146860 25284
rect 146916 25228 146926 25284
rect 38022 25060 38032 25116
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38296 25060 38306 25116
rect 74842 25060 74852 25116
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 75116 25060 75126 25116
rect 111662 25060 111672 25116
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111936 25060 111946 25116
rect 148482 25060 148492 25116
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148756 25060 148766 25116
rect 135314 24556 135324 24612
rect 135380 24556 146412 24612
rect 146468 24556 146860 24612
rect 146916 24556 146926 24612
rect 149200 24500 150000 24528
rect 147746 24444 147756 24500
rect 147812 24444 150000 24500
rect 149200 24416 150000 24444
rect 19612 24276 19622 24332
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19886 24276 19896 24332
rect 56432 24276 56442 24332
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56706 24276 56716 24332
rect 93252 24276 93262 24332
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93526 24276 93536 24332
rect 130072 24276 130082 24332
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130346 24276 130356 24332
rect 125122 23660 125132 23716
rect 125188 23660 146300 23716
rect 146356 23660 146860 23716
rect 146916 23660 146926 23716
rect 147746 23660 147756 23716
rect 147812 23660 148932 23716
rect 148876 23604 148932 23660
rect 149200 23604 150000 23632
rect 148876 23548 150000 23604
rect 38022 23492 38032 23548
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38296 23492 38306 23548
rect 74842 23492 74852 23548
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 75116 23492 75126 23548
rect 111662 23492 111672 23548
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111936 23492 111946 23548
rect 148482 23492 148492 23548
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148756 23492 148766 23548
rect 149200 23520 150000 23548
rect 121874 23100 121884 23156
rect 121940 23100 146412 23156
rect 146468 23100 146860 23156
rect 146916 23100 146926 23156
rect 19612 22708 19622 22764
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19886 22708 19896 22764
rect 56432 22708 56442 22764
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56706 22708 56716 22764
rect 93252 22708 93262 22764
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93526 22708 93536 22764
rect 130072 22708 130082 22764
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130346 22708 130356 22764
rect 149200 22708 150000 22736
rect 147746 22652 147756 22708
rect 147812 22652 150000 22708
rect 149200 22624 150000 22652
rect 115154 22316 115164 22372
rect 115220 22316 146300 22372
rect 146356 22316 146860 22372
rect 146916 22316 146926 22372
rect 38022 21924 38032 21980
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38296 21924 38306 21980
rect 74842 21924 74852 21980
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 75116 21924 75126 21980
rect 111662 21924 111672 21980
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111936 21924 111946 21980
rect 148482 21924 148492 21980
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148756 21924 148766 21980
rect 147746 21868 147756 21924
rect 147812 21868 147822 21924
rect 147756 21812 147812 21868
rect 149200 21812 150000 21840
rect 147756 21756 150000 21812
rect 149200 21728 150000 21756
rect 118402 21420 118412 21476
rect 118468 21420 146412 21476
rect 146468 21420 146860 21476
rect 146916 21420 146926 21476
rect 19612 21140 19622 21196
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19886 21140 19896 21196
rect 56432 21140 56442 21196
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56706 21140 56716 21196
rect 93252 21140 93262 21196
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93526 21140 93536 21196
rect 130072 21140 130082 21196
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130346 21140 130356 21196
rect 149200 20916 150000 20944
rect 147746 20860 147756 20916
rect 147812 20860 150000 20916
rect 149200 20832 150000 20860
rect 114034 20748 114044 20804
rect 114100 20748 146300 20804
rect 146356 20748 146860 20804
rect 146916 20748 146926 20804
rect 38022 20356 38032 20412
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38296 20356 38306 20412
rect 74842 20356 74852 20412
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 75116 20356 75126 20412
rect 111662 20356 111672 20412
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111936 20356 111946 20412
rect 148482 20356 148492 20412
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148756 20356 148766 20412
rect 147746 20188 147756 20244
rect 147812 20188 147822 20244
rect 147756 20020 147812 20188
rect 149200 20020 150000 20048
rect 147756 19964 150000 20020
rect 149200 19936 150000 19964
rect 19612 19572 19622 19628
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19886 19572 19896 19628
rect 56432 19572 56442 19628
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56706 19572 56716 19628
rect 93252 19572 93262 19628
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93526 19572 93536 19628
rect 130072 19572 130082 19628
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130346 19572 130356 19628
rect 119410 19292 119420 19348
rect 119476 19292 135324 19348
rect 135380 19292 135390 19348
rect 110338 19180 110348 19236
rect 110404 19180 146300 19236
rect 146356 19180 146860 19236
rect 146916 19180 146926 19236
rect 149200 19124 150000 19152
rect 147746 19068 147756 19124
rect 147812 19068 150000 19124
rect 149200 19040 150000 19068
rect 38022 18788 38032 18844
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38296 18788 38306 18844
rect 74842 18788 74852 18844
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 75116 18788 75126 18844
rect 111662 18788 111672 18844
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111936 18788 111946 18844
rect 148482 18788 148492 18844
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148756 18788 148766 18844
rect 106754 18284 106764 18340
rect 106820 18284 146412 18340
rect 146468 18284 146860 18340
rect 146916 18284 146926 18340
rect 149200 18228 150000 18256
rect 147746 18172 147756 18228
rect 147812 18172 150000 18228
rect 149200 18144 150000 18172
rect 19612 18004 19622 18060
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19886 18004 19896 18060
rect 56432 18004 56442 18060
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56706 18004 56716 18060
rect 93252 18004 93262 18060
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93526 18004 93536 18060
rect 130072 18004 130082 18060
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130346 18004 130356 18060
rect 119186 17388 119196 17444
rect 119252 17388 146300 17444
rect 146356 17388 146860 17444
rect 146916 17388 146926 17444
rect 147746 17388 147756 17444
rect 147812 17388 148932 17444
rect 148876 17332 148932 17388
rect 149200 17332 150000 17360
rect 148876 17276 150000 17332
rect 38022 17220 38032 17276
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38296 17220 38306 17276
rect 74842 17220 74852 17276
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 75116 17220 75126 17276
rect 111662 17220 111672 17276
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111936 17220 111946 17276
rect 148482 17220 148492 17276
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148756 17220 148766 17276
rect 149200 17248 150000 17276
rect 116610 16940 116620 16996
rect 116676 16940 146412 16996
rect 146468 16940 146860 16996
rect 146916 16940 146926 16996
rect 19612 16436 19622 16492
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19886 16436 19896 16492
rect 56432 16436 56442 16492
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56706 16436 56716 16492
rect 93252 16436 93262 16492
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93526 16436 93536 16492
rect 130072 16436 130082 16492
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130346 16436 130356 16492
rect 149200 16436 150000 16464
rect 147746 16380 147756 16436
rect 147812 16380 150000 16436
rect 149200 16352 150000 16380
rect 108322 15820 108332 15876
rect 108388 15820 146300 15876
rect 146356 15820 146860 15876
rect 146916 15820 146926 15876
rect 38022 15652 38032 15708
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38296 15652 38306 15708
rect 74842 15652 74852 15708
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 75116 15652 75126 15708
rect 111662 15652 111672 15708
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111936 15652 111946 15708
rect 148482 15652 148492 15708
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148756 15652 148766 15708
rect 149200 15540 150000 15568
rect 147746 15484 147756 15540
rect 147812 15484 150000 15540
rect 149200 15456 150000 15484
rect 101826 15372 101836 15428
rect 101892 15372 146412 15428
rect 146468 15372 146860 15428
rect 146916 15372 146926 15428
rect 19612 14868 19622 14924
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19886 14868 19896 14924
rect 56432 14868 56442 14924
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56706 14868 56716 14924
rect 93252 14868 93262 14924
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93526 14868 93536 14924
rect 130072 14868 130082 14924
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130346 14868 130356 14924
rect 149200 14644 150000 14672
rect 147746 14588 147756 14644
rect 147812 14588 150000 14644
rect 149200 14560 150000 14588
rect 100706 14476 100716 14532
rect 100772 14476 146300 14532
rect 146356 14476 146860 14532
rect 146916 14476 146926 14532
rect 105522 14252 105532 14308
rect 105588 14252 119196 14308
rect 119252 14252 119262 14308
rect 38022 14084 38032 14140
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38296 14084 38306 14140
rect 74842 14084 74852 14140
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 75116 14084 75126 14140
rect 111662 14084 111672 14140
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111936 14084 111946 14140
rect 148482 14084 148492 14140
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148756 14084 148766 14140
rect 149200 13748 150000 13776
rect 147746 13692 147756 13748
rect 147812 13692 150000 13748
rect 149200 13664 150000 13692
rect 19612 13300 19622 13356
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19886 13300 19896 13356
rect 56432 13300 56442 13356
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56706 13300 56716 13356
rect 93252 13300 93262 13356
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93526 13300 93536 13356
rect 130072 13300 130082 13356
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130346 13300 130356 13356
rect 99810 12908 99820 12964
rect 99876 12908 146300 12964
rect 146356 12908 146860 12964
rect 146916 12908 146926 12964
rect 149200 12852 150000 12880
rect 147746 12796 147756 12852
rect 147812 12796 150000 12852
rect 149200 12768 150000 12796
rect 38022 12516 38032 12572
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38296 12516 38306 12572
rect 74842 12516 74852 12572
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 75116 12516 75126 12572
rect 111662 12516 111672 12572
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111936 12516 111946 12572
rect 148482 12516 148492 12572
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148756 12516 148766 12572
rect 102834 12012 102844 12068
rect 102900 12012 146412 12068
rect 146468 12012 146860 12068
rect 146916 12012 146926 12068
rect 149200 11956 150000 11984
rect 147746 11900 147756 11956
rect 147812 11900 150000 11956
rect 149200 11872 150000 11900
rect 19612 11732 19622 11788
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19886 11732 19896 11788
rect 56432 11732 56442 11788
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56706 11732 56716 11788
rect 93252 11732 93262 11788
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93526 11732 93536 11788
rect 130072 11732 130082 11788
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130346 11732 130356 11788
rect 120306 11676 120316 11732
rect 120372 11676 123452 11732
rect 123508 11676 123518 11732
rect 115938 11340 115948 11396
rect 116004 11340 146300 11396
rect 146356 11340 146860 11396
rect 146916 11340 146926 11396
rect 98914 11228 98924 11284
rect 98980 11228 99484 11284
rect 99540 11228 99550 11284
rect 147746 11116 147756 11172
rect 147812 11116 148932 11172
rect 148876 11060 148932 11116
rect 149200 11060 150000 11088
rect 148876 11004 150000 11060
rect 38022 10948 38032 11004
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38296 10948 38306 11004
rect 74842 10948 74852 11004
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 75116 10948 75126 11004
rect 111662 10948 111672 11004
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111936 10948 111946 11004
rect 148482 10948 148492 11004
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148756 10948 148766 11004
rect 149200 10976 150000 11004
rect 124002 10892 124012 10948
rect 124068 10892 135212 10948
rect 135268 10892 135278 10948
rect 59490 10444 59500 10500
rect 59556 10444 127708 10500
rect 127764 10444 127774 10500
rect 42690 10332 42700 10388
rect 42756 10332 109564 10388
rect 109620 10332 109630 10388
rect 19612 10164 19622 10220
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19886 10164 19896 10220
rect 56432 10164 56442 10220
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56706 10164 56716 10220
rect 93252 10164 93262 10220
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93526 10164 93536 10220
rect 130072 10164 130082 10220
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130346 10164 130356 10220
rect 149200 10164 150000 10192
rect 99586 10108 99596 10164
rect 99652 10108 102844 10164
rect 102900 10108 102910 10164
rect 105858 10108 105868 10164
rect 105924 10108 116620 10164
rect 116676 10108 116686 10164
rect 147298 10108 147308 10164
rect 147364 10108 148092 10164
rect 148148 10108 150000 10164
rect 149200 10080 150000 10108
rect 38022 9380 38032 9436
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38296 9380 38306 9436
rect 74842 9380 74852 9436
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 75116 9380 75126 9436
rect 111662 9380 111672 9436
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111936 9380 111946 9436
rect 148482 9380 148492 9436
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148756 9380 148766 9436
rect 149200 9268 150000 9296
rect 112130 9212 112140 9268
rect 112196 9212 118412 9268
rect 118468 9212 118478 9268
rect 147298 9212 147308 9268
rect 147364 9212 148092 9268
rect 148148 9212 150000 9268
rect 149200 9184 150000 9212
rect 90738 9100 90748 9156
rect 90804 9100 147756 9156
rect 147812 9100 147822 9156
rect 41346 8988 41356 9044
rect 41412 8988 110572 9044
rect 110628 8988 110638 9044
rect 147298 8988 147308 9044
rect 147364 8988 148092 9044
rect 148148 8988 148158 9044
rect 15138 8876 15148 8932
rect 15204 8876 82908 8932
rect 82964 8876 82974 8932
rect 17490 8764 17500 8820
rect 17556 8764 83916 8820
rect 83972 8764 83982 8820
rect 90514 8764 90524 8820
rect 90580 8764 147644 8820
rect 147700 8764 147710 8820
rect 19612 8596 19622 8652
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19886 8596 19896 8652
rect 56432 8596 56442 8652
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56706 8596 56716 8652
rect 93252 8596 93262 8652
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93526 8596 93536 8652
rect 130072 8596 130082 8652
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130346 8596 130356 8652
rect 53106 8428 53116 8484
rect 53172 8428 123676 8484
rect 123732 8428 123742 8484
rect 148082 8428 148092 8484
rect 148148 8428 148158 8484
rect 148092 8372 148148 8428
rect 149200 8372 150000 8400
rect 148092 8316 150000 8372
rect 149200 8288 150000 8316
rect 127586 8092 127596 8148
rect 127652 8092 134876 8148
rect 134932 8092 135324 8148
rect 135380 8092 147532 8148
rect 147588 8092 147598 8148
rect 147298 7980 147308 8036
rect 147364 7980 148092 8036
rect 148148 7980 148158 8036
rect 38022 7812 38032 7868
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38296 7812 38306 7868
rect 74842 7812 74852 7868
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 75116 7812 75126 7868
rect 111662 7812 111672 7868
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111936 7812 111946 7868
rect 148482 7812 148492 7868
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148756 7812 148766 7868
rect 113474 7756 113484 7812
rect 113540 7756 115948 7812
rect 116004 7756 116014 7812
rect 51090 7644 51100 7700
rect 51156 7644 121436 7700
rect 121492 7644 121502 7700
rect 39106 7532 39116 7588
rect 39172 7532 109004 7588
rect 109060 7532 109070 7588
rect 125346 7532 125356 7588
rect 125412 7532 148204 7588
rect 148260 7532 148270 7588
rect 149200 7476 150000 7504
rect 57250 7420 57260 7476
rect 57316 7420 88956 7476
rect 89012 7420 89022 7476
rect 148082 7420 148092 7476
rect 148148 7420 150000 7476
rect 149200 7392 150000 7420
rect 13458 7308 13468 7364
rect 13524 7308 80556 7364
rect 80612 7308 80622 7364
rect 82226 7308 82236 7364
rect 82292 7308 146076 7364
rect 146132 7308 146142 7364
rect 21634 7196 21644 7252
rect 21700 7196 87276 7252
rect 87332 7196 87342 7252
rect 88386 7196 88396 7252
rect 88452 7196 147756 7252
rect 147812 7196 147822 7252
rect 19612 7028 19622 7084
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19886 7028 19896 7084
rect 56432 7028 56442 7084
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56706 7028 56716 7084
rect 93252 7028 93262 7084
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93526 7028 93536 7084
rect 130072 7028 130082 7084
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130346 7028 130356 7084
rect 71250 6860 71260 6916
rect 71316 6860 143276 6916
rect 143332 6860 143342 6916
rect 22530 6748 22540 6804
rect 22596 6748 114268 6804
rect 114324 6748 114334 6804
rect 118514 6748 118524 6804
rect 118580 6748 125132 6804
rect 125188 6748 125198 6804
rect 137778 6748 137788 6804
rect 137844 6748 147868 6804
rect 147924 6748 147934 6804
rect 77634 6636 77644 6692
rect 77700 6636 147644 6692
rect 147700 6636 147710 6692
rect 149200 6580 150000 6608
rect 35970 6524 35980 6580
rect 36036 6524 105644 6580
rect 105700 6524 105710 6580
rect 127698 6524 127708 6580
rect 127764 6524 129276 6580
rect 129332 6524 129836 6580
rect 129892 6524 129902 6580
rect 147298 6524 147308 6580
rect 147364 6524 148092 6580
rect 148148 6524 150000 6580
rect 149200 6496 150000 6524
rect 102452 6412 114268 6468
rect 102452 6356 102508 6412
rect 84466 6300 84476 6356
rect 84532 6300 86940 6356
rect 86996 6300 102508 6356
rect 114212 6356 114268 6412
rect 114212 6300 147756 6356
rect 147812 6300 147822 6356
rect 38022 6244 38032 6300
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38296 6244 38306 6300
rect 74842 6244 74852 6300
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 75116 6244 75126 6300
rect 111662 6244 111672 6300
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111936 6244 111946 6300
rect 148482 6244 148492 6300
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148756 6244 148766 6300
rect 76066 6188 76076 6244
rect 76132 6188 102508 6244
rect 102452 6132 102508 6188
rect 114212 6188 136556 6244
rect 136612 6188 136622 6244
rect 114212 6132 114268 6188
rect 102452 6076 114268 6132
rect 85362 5964 85372 6020
rect 85428 5964 147756 6020
rect 147812 5964 147822 6020
rect 11778 5852 11788 5908
rect 11844 5852 79660 5908
rect 79716 5852 79726 5908
rect 103058 5852 103068 5908
rect 103124 5852 103964 5908
rect 104020 5852 104412 5908
rect 104468 5852 111244 5908
rect 111300 5852 111468 5908
rect 111524 5852 117852 5908
rect 117908 5852 117918 5908
rect 140130 5852 140140 5908
rect 140196 5852 141372 5908
rect 141428 5852 141438 5908
rect 10098 5740 10108 5796
rect 10164 5740 77868 5796
rect 77924 5740 77934 5796
rect 123890 5740 123900 5796
rect 123956 5740 124348 5796
rect 124404 5740 124414 5796
rect 139906 5740 139916 5796
rect 139972 5740 140924 5796
rect 140980 5740 140990 5796
rect 149200 5684 150000 5712
rect 30706 5628 30716 5684
rect 30772 5628 97132 5684
rect 97188 5628 97198 5684
rect 147298 5628 147308 5684
rect 147364 5628 148092 5684
rect 148148 5628 150000 5684
rect 149200 5600 150000 5628
rect 19612 5460 19622 5516
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19886 5460 19896 5516
rect 56432 5460 56442 5516
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56706 5460 56716 5516
rect 93252 5460 93262 5516
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93526 5460 93536 5516
rect 130072 5460 130082 5516
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130346 5460 130356 5516
rect 55906 5292 55916 5348
rect 55972 5292 125916 5348
rect 125972 5292 125982 5348
rect 61282 5180 61292 5236
rect 61348 5180 85596 5236
rect 85652 5180 85662 5236
rect 87602 5180 87612 5236
rect 87668 5180 88060 5236
rect 88116 5180 89404 5236
rect 89460 5180 90188 5236
rect 90244 5180 90748 5236
rect 90804 5180 90814 5236
rect 109554 5180 109564 5236
rect 109620 5180 111020 5236
rect 111076 5180 111086 5236
rect 114034 5180 114044 5236
rect 114100 5180 115388 5236
rect 115444 5180 133084 5236
rect 133140 5180 133150 5236
rect 133298 5180 133308 5236
rect 133364 5180 136892 5236
rect 136948 5180 136958 5236
rect 133084 5124 133140 5180
rect 9650 5068 9660 5124
rect 9716 5068 75180 5124
rect 75236 5068 75246 5124
rect 75842 5068 75852 5124
rect 75908 5068 76972 5124
rect 77028 5068 77644 5124
rect 77700 5068 77710 5124
rect 78194 5068 78204 5124
rect 78260 5068 78540 5124
rect 78596 5068 78876 5124
rect 78932 5068 79436 5124
rect 79492 5068 79502 5124
rect 83234 5068 83244 5124
rect 83300 5068 83580 5124
rect 83636 5068 84588 5124
rect 84644 5068 85372 5124
rect 85428 5068 85438 5124
rect 99250 5068 99260 5124
rect 99316 5068 99484 5124
rect 99540 5068 99550 5124
rect 102610 5068 102620 5124
rect 102676 5068 103068 5124
rect 103124 5068 103134 5124
rect 104290 5068 104300 5124
rect 104356 5068 108332 5124
rect 108388 5068 108398 5124
rect 111794 5068 111804 5124
rect 111860 5068 112252 5124
rect 112308 5068 112318 5124
rect 117618 5068 117628 5124
rect 117684 5068 117852 5124
rect 117908 5068 127036 5124
rect 127092 5068 127102 5124
rect 133084 5068 140924 5124
rect 140980 5068 141596 5124
rect 141652 5068 143500 5124
rect 143556 5068 143566 5124
rect 75852 5012 75908 5068
rect 75506 4956 75516 5012
rect 75572 4956 75908 5012
rect 78932 4956 100380 5012
rect 100436 4956 100446 5012
rect 100594 4956 100604 5012
rect 100660 4956 102060 5012
rect 102116 4956 102126 5012
rect 102834 4956 102844 5012
rect 102900 4956 103740 5012
rect 103796 4956 103806 5012
rect 112130 4956 112140 5012
rect 112196 4956 112812 5012
rect 112868 4956 112878 5012
rect 113138 4956 113148 5012
rect 113204 4956 115164 5012
rect 115220 4956 115230 5012
rect 115602 4956 115612 5012
rect 115668 4956 115948 5012
rect 116004 4956 116014 5012
rect 116274 4956 116284 5012
rect 116340 4956 121884 5012
rect 121940 4956 121950 5012
rect 126690 4956 126700 5012
rect 126756 4956 129052 5012
rect 129108 4956 129118 5012
rect 132402 4956 132412 5012
rect 132468 4956 132972 5012
rect 133028 4956 133038 5012
rect 134082 4956 134092 5012
rect 134148 4956 134652 5012
rect 134708 4956 135548 5012
rect 135604 4956 135614 5012
rect 78932 4900 78988 4956
rect 134092 4900 134148 4956
rect 60386 4844 60396 4900
rect 60452 4844 78988 4900
rect 85922 4844 85932 4900
rect 85988 4844 86380 4900
rect 86436 4844 87948 4900
rect 88004 4844 88014 4900
rect 89282 4844 89292 4900
rect 89348 4844 89740 4900
rect 89796 4844 90524 4900
rect 90580 4844 90590 4900
rect 97570 4844 97580 4900
rect 97636 4844 98364 4900
rect 98420 4844 98430 4900
rect 102452 4844 112084 4900
rect 114146 4844 114156 4900
rect 114212 4844 114604 4900
rect 114660 4844 114670 4900
rect 129602 4844 129612 4900
rect 129668 4844 130620 4900
rect 130676 4844 131628 4900
rect 131684 4844 132076 4900
rect 132132 4844 134148 4900
rect 139682 4844 139692 4900
rect 139748 4844 140252 4900
rect 140308 4844 141148 4900
rect 141204 4844 141214 4900
rect 147298 4844 147308 4900
rect 147364 4844 148092 4900
rect 148148 4844 148932 4900
rect 102452 4788 102508 4844
rect 80882 4732 80892 4788
rect 80948 4732 81340 4788
rect 81396 4732 82124 4788
rect 82180 4732 82684 4788
rect 82740 4732 102508 4788
rect 112028 4788 112084 4844
rect 148876 4788 148932 4844
rect 149200 4788 150000 4816
rect 112028 4732 147756 4788
rect 147812 4732 147822 4788
rect 148876 4732 150000 4788
rect 38022 4676 38032 4732
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38296 4676 38306 4732
rect 74842 4676 74852 4732
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 75116 4676 75126 4732
rect 111662 4676 111672 4732
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111936 4676 111946 4732
rect 148482 4676 148492 4732
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148756 4676 148766 4732
rect 149200 4704 150000 4732
rect 102452 4620 109900 4676
rect 109956 4620 109966 4676
rect 130498 4620 130508 4676
rect 130564 4620 137844 4676
rect 138226 4620 138236 4676
rect 138292 4620 139132 4676
rect 139188 4620 139198 4676
rect 141810 4620 141820 4676
rect 141876 4620 143724 4676
rect 143780 4620 143790 4676
rect 143948 4620 147980 4676
rect 148036 4620 148046 4676
rect 102452 4564 102508 4620
rect 137788 4564 137844 4620
rect 10994 4508 11004 4564
rect 11060 4508 11340 4564
rect 11396 4508 11788 4564
rect 11844 4508 11854 4564
rect 13010 4508 13020 4564
rect 13076 4508 13468 4564
rect 13524 4508 13534 4564
rect 42466 4508 42476 4564
rect 42532 4508 102508 4564
rect 103506 4508 103516 4564
rect 103572 4508 103582 4564
rect 105634 4508 105644 4564
rect 105700 4508 106988 4564
rect 107044 4508 107054 4564
rect 110562 4508 110572 4564
rect 110628 4508 112140 4564
rect 112196 4508 112206 4564
rect 117058 4508 117068 4564
rect 117124 4508 118188 4564
rect 118244 4508 118254 4564
rect 127250 4508 127260 4564
rect 127316 4508 127932 4564
rect 127988 4508 127998 4564
rect 132850 4508 132860 4564
rect 132916 4508 133868 4564
rect 133924 4508 133934 4564
rect 137788 4508 139860 4564
rect 142146 4508 142156 4564
rect 142212 4508 142828 4564
rect 142884 4508 142894 4564
rect 18946 4396 18956 4452
rect 19012 4396 19404 4452
rect 19460 4396 61292 4452
rect 61348 4396 61358 4452
rect 73938 4396 73948 4452
rect 74004 4396 75292 4452
rect 75348 4396 76076 4452
rect 76132 4396 76142 4452
rect 79986 4396 79996 4452
rect 80052 4396 80444 4452
rect 80500 4396 81340 4452
rect 81396 4396 82124 4452
rect 82180 4396 82190 4452
rect 90514 4396 90524 4452
rect 90580 4396 91308 4452
rect 91364 4396 91374 4452
rect 97682 4396 97692 4452
rect 97748 4396 100716 4452
rect 100772 4396 100782 4452
rect 103516 4340 103572 4508
rect 139804 4452 139860 4508
rect 143948 4452 144004 4620
rect 146066 4508 146076 4564
rect 146132 4508 147756 4564
rect 147812 4508 147822 4564
rect 109778 4396 109788 4452
rect 109844 4396 112476 4452
rect 112532 4396 112542 4452
rect 122658 4396 122668 4452
rect 122724 4396 124012 4452
rect 124068 4396 124796 4452
rect 124852 4396 126700 4452
rect 126756 4396 126766 4452
rect 135090 4396 135100 4452
rect 135156 4396 136332 4452
rect 136388 4396 136398 4452
rect 136770 4396 136780 4452
rect 136836 4396 137228 4452
rect 137284 4396 137294 4452
rect 137732 4396 139580 4452
rect 139636 4396 139646 4452
rect 139804 4396 144004 4452
rect 145170 4396 145180 4452
rect 145236 4396 146860 4452
rect 146916 4396 146926 4452
rect 137732 4340 137788 4396
rect 8306 4284 8316 4340
rect 8372 4284 8876 4340
rect 8932 4284 9660 4340
rect 9716 4284 9726 4340
rect 9996 4284 73388 4340
rect 73444 4284 73454 4340
rect 99810 4284 99820 4340
rect 99876 4284 101052 4340
rect 101108 4284 101118 4340
rect 102722 4284 102732 4340
rect 102788 4284 104188 4340
rect 104244 4284 105308 4340
rect 105364 4284 105374 4340
rect 110002 4284 110012 4340
rect 110068 4284 110460 4340
rect 110516 4284 110796 4340
rect 110852 4284 111468 4340
rect 111524 4284 111804 4340
rect 111860 4284 111870 4340
rect 119634 4284 119644 4340
rect 119700 4284 120988 4340
rect 121044 4284 121054 4340
rect 129378 4284 129388 4340
rect 129444 4284 129612 4340
rect 129668 4284 129678 4340
rect 136098 4284 136108 4340
rect 136164 4284 137116 4340
rect 137172 4284 137788 4340
rect 142930 4284 142940 4340
rect 142996 4284 144060 4340
rect 144116 4284 145292 4340
rect 145348 4284 145358 4340
rect 9996 4228 10052 4284
rect 6626 4172 6636 4228
rect 6692 4172 10052 4228
rect 16930 4172 16940 4228
rect 16996 4172 17948 4228
rect 18004 4172 18014 4228
rect 32050 4172 32060 4228
rect 32116 4172 32620 4228
rect 32676 4172 32686 4228
rect 43810 4172 43820 4228
rect 43876 4172 44380 4228
rect 44436 4172 44446 4228
rect 55570 4172 55580 4228
rect 55636 4172 56140 4228
rect 56196 4172 56206 4228
rect 67330 4172 67340 4228
rect 67396 4172 67900 4228
rect 67956 4172 67966 4228
rect 72482 4172 72492 4228
rect 72548 4172 73276 4228
rect 73332 4172 73342 4228
rect 85810 4172 85820 4228
rect 85876 4172 86716 4228
rect 86772 4172 86782 4228
rect 86940 4172 98196 4228
rect 98354 4172 98364 4228
rect 98420 4172 98700 4228
rect 98756 4172 100492 4228
rect 100548 4172 100558 4228
rect 108546 4172 108556 4228
rect 108612 4172 109340 4228
rect 109396 4172 109406 4228
rect 141362 4172 141372 4228
rect 141428 4172 142828 4228
rect 142884 4172 143052 4228
rect 143108 4172 143118 4228
rect 143266 4172 143276 4228
rect 143332 4172 144844 4228
rect 144900 4172 144910 4228
rect 146402 4172 146412 4228
rect 146468 4172 147084 4228
rect 147140 4172 147150 4228
rect 86940 4116 86996 4172
rect 98140 4116 98196 4172
rect 54226 4060 54236 4116
rect 54292 4060 86996 4116
rect 90692 4060 95844 4116
rect 98140 4060 99596 4116
rect 99652 4060 99932 4116
rect 99988 4060 99998 4116
rect 102050 4060 102060 4116
rect 102116 4060 102956 4116
rect 103012 4060 103022 4116
rect 121650 4060 121660 4116
rect 121716 4060 122892 4116
rect 122948 4060 122958 4116
rect 125972 4060 137228 4116
rect 137284 4060 137294 4116
rect 90692 4004 90748 4060
rect 66210 3948 66220 4004
rect 66276 3948 90748 4004
rect 95788 4004 95844 4060
rect 125972 4004 126028 4060
rect 95788 3948 126028 4004
rect 19612 3892 19622 3948
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19886 3892 19896 3948
rect 56432 3892 56442 3948
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56706 3892 56716 3948
rect 93252 3892 93262 3948
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93526 3892 93536 3948
rect 130072 3892 130082 3948
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130346 3892 130356 3948
rect 149200 3892 150000 3920
rect 112242 3836 112252 3892
rect 112308 3836 114044 3892
rect 114100 3836 114110 3892
rect 115042 3836 115052 3892
rect 115108 3836 115948 3892
rect 116004 3836 116014 3892
rect 123666 3836 123676 3892
rect 123732 3836 126028 3892
rect 126084 3836 126094 3892
rect 128258 3836 128268 3892
rect 128324 3836 129724 3892
rect 129780 3836 129790 3892
rect 137732 3836 139692 3892
rect 139748 3836 139758 3892
rect 145954 3836 145964 3892
rect 146020 3836 148092 3892
rect 148148 3836 150000 3892
rect 137732 3780 137788 3836
rect 149200 3808 150000 3836
rect 72818 3724 72828 3780
rect 72884 3724 137788 3780
rect 143154 3724 143164 3780
rect 143220 3724 143836 3780
rect 143892 3724 143902 3780
rect 22642 3612 22652 3668
rect 22708 3612 22988 3668
rect 23044 3612 57260 3668
rect 57316 3612 57326 3668
rect 62626 3612 62636 3668
rect 62692 3612 104076 3668
rect 104132 3612 104142 3668
rect 107874 3612 107884 3668
rect 107940 3612 107950 3668
rect 109890 3612 109900 3668
rect 109956 3612 111692 3668
rect 111748 3612 111758 3668
rect 113932 3612 116172 3668
rect 116228 3612 116508 3668
rect 116564 3612 116574 3668
rect 120978 3612 120988 3668
rect 121044 3612 131292 3668
rect 131348 3612 131358 3668
rect 136434 3612 136444 3668
rect 136500 3612 139356 3668
rect 139412 3612 139422 3668
rect 107884 3556 107940 3612
rect 113932 3556 113988 3612
rect 8866 3500 8876 3556
rect 8932 3500 9772 3556
rect 9828 3500 9838 3556
rect 16706 3500 16716 3556
rect 16772 3500 17500 3556
rect 17556 3500 17566 3556
rect 20066 3500 20076 3556
rect 20132 3500 20636 3556
rect 20692 3500 21644 3556
rect 21700 3500 21710 3556
rect 80770 3500 80780 3556
rect 80836 3500 82684 3556
rect 82740 3500 82750 3556
rect 92530 3500 92540 3556
rect 92596 3500 93772 3556
rect 93828 3500 93838 3556
rect 96450 3500 96460 3556
rect 96516 3500 98588 3556
rect 98644 3500 98654 3556
rect 102946 3500 102956 3556
rect 103012 3500 104636 3556
rect 104692 3500 104702 3556
rect 106082 3500 106092 3556
rect 106148 3500 106764 3556
rect 106820 3500 107940 3556
rect 108210 3500 108220 3556
rect 108276 3500 110236 3556
rect 110292 3500 110302 3556
rect 112802 3500 112812 3556
rect 112868 3500 113988 3556
rect 114146 3500 114156 3556
rect 114212 3500 114604 3556
rect 114660 3500 114670 3556
rect 116722 3500 116732 3556
rect 116788 3500 118412 3556
rect 118468 3500 119644 3556
rect 119700 3500 119710 3556
rect 122546 3500 122556 3556
rect 122612 3500 124236 3556
rect 124292 3500 124302 3556
rect 126130 3500 126140 3556
rect 126196 3500 127484 3556
rect 127540 3500 128828 3556
rect 128884 3500 128894 3556
rect 129378 3500 129388 3556
rect 129444 3500 131068 3556
rect 131124 3500 131404 3556
rect 131460 3500 131740 3556
rect 131796 3500 131806 3556
rect 137890 3500 137900 3556
rect 137956 3500 141148 3556
rect 141204 3500 141214 3556
rect 142156 3500 145628 3556
rect 145684 3500 145694 3556
rect 142156 3444 142212 3500
rect 5170 3388 5180 3444
rect 5236 3388 6076 3444
rect 6132 3388 6142 3444
rect 15250 3388 15260 3444
rect 15316 3388 15820 3444
rect 15876 3388 15886 3444
rect 18610 3388 18620 3444
rect 18676 3388 19180 3444
rect 19236 3388 19246 3444
rect 20290 3388 20300 3444
rect 20356 3388 21756 3444
rect 21812 3388 21822 3444
rect 28690 3388 28700 3444
rect 28756 3388 29260 3444
rect 29316 3388 29326 3444
rect 40450 3388 40460 3444
rect 40516 3388 41020 3444
rect 41076 3388 41086 3444
rect 52210 3388 52220 3444
rect 52276 3388 52780 3444
rect 52836 3388 52846 3444
rect 63970 3388 63980 3444
rect 64036 3388 64540 3444
rect 64596 3388 64606 3444
rect 75730 3388 75740 3444
rect 75796 3388 77196 3444
rect 77252 3388 77262 3444
rect 77420 3388 78764 3444
rect 78820 3388 78830 3444
rect 79090 3388 79100 3444
rect 79156 3388 81116 3444
rect 81172 3388 81182 3444
rect 82450 3388 82460 3444
rect 82516 3388 83356 3444
rect 83412 3388 83422 3444
rect 84130 3388 84140 3444
rect 84196 3388 84700 3444
rect 84756 3388 84766 3444
rect 87490 3388 87500 3444
rect 87556 3388 88956 3444
rect 89012 3388 89022 3444
rect 89170 3388 89180 3444
rect 89236 3388 90524 3444
rect 90580 3388 90590 3444
rect 90860 3388 92876 3444
rect 92932 3388 92942 3444
rect 97122 3388 97132 3444
rect 97188 3388 97804 3444
rect 97860 3388 97870 3444
rect 104402 3388 104412 3444
rect 104468 3388 105980 3444
rect 106036 3388 107436 3444
rect 107492 3388 107502 3444
rect 107874 3388 107884 3444
rect 107940 3388 108668 3444
rect 108724 3388 108734 3444
rect 108994 3388 109004 3444
rect 109060 3388 109452 3444
rect 109508 3388 109518 3444
rect 111010 3388 111020 3444
rect 111076 3388 113372 3444
rect 113428 3388 113820 3444
rect 113876 3388 113886 3444
rect 114034 3388 114044 3444
rect 114100 3388 114380 3444
rect 114436 3388 114446 3444
rect 116050 3388 116060 3444
rect 116116 3388 117180 3444
rect 117236 3388 117740 3444
rect 117796 3388 117806 3444
rect 119186 3388 119196 3444
rect 119252 3388 119532 3444
rect 119588 3388 119598 3444
rect 122210 3388 122220 3444
rect 122276 3388 122780 3444
rect 122836 3388 122846 3444
rect 124450 3388 124460 3444
rect 124516 3388 125580 3444
rect 125636 3388 128044 3444
rect 128100 3388 128110 3444
rect 131170 3388 131180 3444
rect 131236 3388 132748 3444
rect 132804 3388 133420 3444
rect 133476 3388 133486 3444
rect 136210 3388 136220 3444
rect 136276 3388 137340 3444
rect 137396 3388 138124 3444
rect 138180 3388 138190 3444
rect 139682 3388 139692 3444
rect 139748 3388 142156 3444
rect 142212 3388 142222 3444
rect 145058 3388 145068 3444
rect 145124 3388 146076 3444
rect 146132 3388 146142 3444
rect 146514 3388 146524 3444
rect 146580 3388 148092 3444
rect 148148 3388 148158 3444
rect 77420 3332 77476 3388
rect 90860 3332 90916 3388
rect 25890 3276 25900 3332
rect 25956 3276 30716 3332
rect 30772 3276 30782 3332
rect 37650 3276 37660 3332
rect 37716 3276 39116 3332
rect 39172 3276 39182 3332
rect 39330 3276 39340 3332
rect 39396 3276 42476 3332
rect 42532 3276 42542 3332
rect 54450 3276 54460 3332
rect 54516 3276 56924 3332
rect 56980 3276 56990 3332
rect 57810 3276 57820 3332
rect 57876 3276 64092 3332
rect 64148 3276 64158 3332
rect 77410 3276 77420 3332
rect 77476 3276 77486 3332
rect 90850 3276 90860 3332
rect 90916 3276 90926 3332
rect 94994 3276 95004 3332
rect 95060 3276 99148 3332
rect 99204 3276 99214 3332
rect 111234 3276 111244 3332
rect 111300 3276 113484 3332
rect 113540 3276 113550 3332
rect 113922 3276 113932 3332
rect 113988 3276 114156 3332
rect 114212 3276 114222 3332
rect 132066 3276 132076 3332
rect 132132 3276 133084 3332
rect 133140 3276 133150 3332
rect 134204 3276 139468 3332
rect 139524 3276 139534 3332
rect 140018 3276 140028 3332
rect 140084 3276 141820 3332
rect 141876 3276 141886 3332
rect 142034 3276 142044 3332
rect 142100 3276 144844 3332
rect 144900 3276 144910 3332
rect 132514 3164 132524 3220
rect 132580 3164 133980 3220
rect 134036 3164 134046 3220
rect 38022 3108 38032 3164
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38296 3108 38306 3164
rect 74842 3108 74852 3164
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 75116 3108 75126 3164
rect 111662 3108 111672 3164
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111936 3108 111946 3164
rect 27570 2940 27580 2996
rect 27636 2940 54236 2996
rect 54292 2940 54302 2996
rect 62850 2940 62860 2996
rect 62916 2940 131852 2996
rect 131908 2940 131918 2996
rect 134204 2884 134260 3276
rect 136546 3164 136556 3220
rect 136612 3164 146860 3220
rect 146916 3164 146926 3220
rect 148482 3108 148492 3164
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148756 3108 148766 3164
rect 139458 3052 139468 3108
rect 139524 3052 141036 3108
rect 141092 3052 141102 3108
rect 149200 2996 150000 3024
rect 147074 2940 147084 2996
rect 147140 2940 150000 2996
rect 149200 2912 150000 2940
rect 29586 2828 29596 2884
rect 29652 2828 60396 2884
rect 60452 2828 60462 2884
rect 74610 2828 74620 2884
rect 74676 2828 134260 2884
rect 30930 2716 30940 2772
rect 30996 2716 95676 2772
rect 95732 2716 95742 2772
rect 61170 2604 61180 2660
rect 61236 2604 120988 2660
rect 121044 2604 121054 2660
rect 32386 2492 32396 2548
rect 32452 2492 62636 2548
rect 62692 2492 62702 2548
rect 64866 2492 64876 2548
rect 64932 2492 112476 2548
rect 112532 2492 112542 2548
rect 34290 2380 34300 2436
rect 34356 2380 102844 2436
rect 102900 2380 102910 2436
rect 94098 2268 94108 2324
rect 94164 2268 113596 2324
rect 113652 2268 113662 2324
rect 69570 2156 69580 2212
rect 69636 2156 138684 2212
rect 138740 2156 138750 2212
rect 149200 2100 150000 2128
rect 67666 2044 67676 2100
rect 67732 2044 136444 2100
rect 136500 2044 136510 2100
rect 148082 2044 148092 2100
rect 148148 2044 150000 2100
rect 149200 2016 150000 2044
rect 95666 1596 95676 1652
rect 95732 1596 101612 1652
rect 101668 1596 101678 1652
rect 24210 1484 24220 1540
rect 24276 1484 98476 1540
rect 98532 1484 98542 1540
rect 112466 1484 112476 1540
rect 112532 1484 135548 1540
rect 135604 1484 135614 1540
rect 49410 1372 49420 1428
rect 49476 1372 119532 1428
rect 119588 1372 119598 1428
rect 46050 1260 46060 1316
rect 46116 1260 115948 1316
rect 116004 1260 116014 1316
rect 149200 1204 150000 1232
rect 44146 1148 44156 1204
rect 44212 1148 112812 1204
rect 112868 1148 112878 1204
rect 117814 1148 117852 1204
rect 117908 1148 117918 1204
rect 120932 1148 124348 1204
rect 124404 1148 124414 1204
rect 147186 1148 147196 1204
rect 147252 1148 150000 1204
rect 120932 1092 120988 1148
rect 149200 1120 150000 1148
rect 56914 1036 56924 1092
rect 56980 1036 120988 1092
rect 64082 924 64092 980
rect 64148 924 128940 980
rect 128996 924 129006 980
rect 47730 812 47740 868
rect 47796 812 55468 868
rect 78866 812 78876 868
rect 78932 812 145180 868
rect 145236 812 145246 868
rect 55412 756 55468 812
rect 55412 700 117852 756
rect 117908 700 117918 756
<< via3 >>
rect 19622 36820 19678 36876
rect 19726 36820 19782 36876
rect 19830 36820 19886 36876
rect 56442 36820 56498 36876
rect 56546 36820 56602 36876
rect 56650 36820 56706 36876
rect 93262 36820 93318 36876
rect 93366 36820 93422 36876
rect 93470 36820 93526 36876
rect 130082 36820 130138 36876
rect 130186 36820 130242 36876
rect 130290 36820 130346 36876
rect 38032 36036 38088 36092
rect 38136 36036 38192 36092
rect 38240 36036 38296 36092
rect 74852 36036 74908 36092
rect 74956 36036 75012 36092
rect 75060 36036 75116 36092
rect 111672 36036 111728 36092
rect 111776 36036 111832 36092
rect 111880 36036 111936 36092
rect 148492 36036 148548 36092
rect 148596 36036 148652 36092
rect 148700 36036 148756 36092
rect 19622 35252 19678 35308
rect 19726 35252 19782 35308
rect 19830 35252 19886 35308
rect 56442 35252 56498 35308
rect 56546 35252 56602 35308
rect 56650 35252 56706 35308
rect 93262 35252 93318 35308
rect 93366 35252 93422 35308
rect 93470 35252 93526 35308
rect 130082 35252 130138 35308
rect 130186 35252 130242 35308
rect 130290 35252 130346 35308
rect 38032 34468 38088 34524
rect 38136 34468 38192 34524
rect 38240 34468 38296 34524
rect 74852 34468 74908 34524
rect 74956 34468 75012 34524
rect 75060 34468 75116 34524
rect 111672 34468 111728 34524
rect 111776 34468 111832 34524
rect 111880 34468 111936 34524
rect 148492 34468 148548 34524
rect 148596 34468 148652 34524
rect 148700 34468 148756 34524
rect 19622 33684 19678 33740
rect 19726 33684 19782 33740
rect 19830 33684 19886 33740
rect 56442 33684 56498 33740
rect 56546 33684 56602 33740
rect 56650 33684 56706 33740
rect 93262 33684 93318 33740
rect 93366 33684 93422 33740
rect 93470 33684 93526 33740
rect 130082 33684 130138 33740
rect 130186 33684 130242 33740
rect 130290 33684 130346 33740
rect 38032 32900 38088 32956
rect 38136 32900 38192 32956
rect 38240 32900 38296 32956
rect 74852 32900 74908 32956
rect 74956 32900 75012 32956
rect 75060 32900 75116 32956
rect 111672 32900 111728 32956
rect 111776 32900 111832 32956
rect 111880 32900 111936 32956
rect 148492 32900 148548 32956
rect 148596 32900 148652 32956
rect 148700 32900 148756 32956
rect 19622 32116 19678 32172
rect 19726 32116 19782 32172
rect 19830 32116 19886 32172
rect 56442 32116 56498 32172
rect 56546 32116 56602 32172
rect 56650 32116 56706 32172
rect 93262 32116 93318 32172
rect 93366 32116 93422 32172
rect 93470 32116 93526 32172
rect 130082 32116 130138 32172
rect 130186 32116 130242 32172
rect 130290 32116 130346 32172
rect 38032 31332 38088 31388
rect 38136 31332 38192 31388
rect 38240 31332 38296 31388
rect 74852 31332 74908 31388
rect 74956 31332 75012 31388
rect 75060 31332 75116 31388
rect 111672 31332 111728 31388
rect 111776 31332 111832 31388
rect 111880 31332 111936 31388
rect 148492 31332 148548 31388
rect 148596 31332 148652 31388
rect 148700 31332 148756 31388
rect 19622 30548 19678 30604
rect 19726 30548 19782 30604
rect 19830 30548 19886 30604
rect 56442 30548 56498 30604
rect 56546 30548 56602 30604
rect 56650 30548 56706 30604
rect 93262 30548 93318 30604
rect 93366 30548 93422 30604
rect 93470 30548 93526 30604
rect 130082 30548 130138 30604
rect 130186 30548 130242 30604
rect 130290 30548 130346 30604
rect 38032 29764 38088 29820
rect 38136 29764 38192 29820
rect 38240 29764 38296 29820
rect 74852 29764 74908 29820
rect 74956 29764 75012 29820
rect 75060 29764 75116 29820
rect 111672 29764 111728 29820
rect 111776 29764 111832 29820
rect 111880 29764 111936 29820
rect 148492 29764 148548 29820
rect 148596 29764 148652 29820
rect 148700 29764 148756 29820
rect 19622 28980 19678 29036
rect 19726 28980 19782 29036
rect 19830 28980 19886 29036
rect 56442 28980 56498 29036
rect 56546 28980 56602 29036
rect 56650 28980 56706 29036
rect 93262 28980 93318 29036
rect 93366 28980 93422 29036
rect 93470 28980 93526 29036
rect 130082 28980 130138 29036
rect 130186 28980 130242 29036
rect 130290 28980 130346 29036
rect 38032 28196 38088 28252
rect 38136 28196 38192 28252
rect 38240 28196 38296 28252
rect 74852 28196 74908 28252
rect 74956 28196 75012 28252
rect 75060 28196 75116 28252
rect 111672 28196 111728 28252
rect 111776 28196 111832 28252
rect 111880 28196 111936 28252
rect 148492 28196 148548 28252
rect 148596 28196 148652 28252
rect 148700 28196 148756 28252
rect 19622 27412 19678 27468
rect 19726 27412 19782 27468
rect 19830 27412 19886 27468
rect 56442 27412 56498 27468
rect 56546 27412 56602 27468
rect 56650 27412 56706 27468
rect 93262 27412 93318 27468
rect 93366 27412 93422 27468
rect 93470 27412 93526 27468
rect 130082 27412 130138 27468
rect 130186 27412 130242 27468
rect 130290 27412 130346 27468
rect 38032 26628 38088 26684
rect 38136 26628 38192 26684
rect 38240 26628 38296 26684
rect 74852 26628 74908 26684
rect 74956 26628 75012 26684
rect 75060 26628 75116 26684
rect 111672 26628 111728 26684
rect 111776 26628 111832 26684
rect 111880 26628 111936 26684
rect 148492 26628 148548 26684
rect 148596 26628 148652 26684
rect 148700 26628 148756 26684
rect 19622 25844 19678 25900
rect 19726 25844 19782 25900
rect 19830 25844 19886 25900
rect 56442 25844 56498 25900
rect 56546 25844 56602 25900
rect 56650 25844 56706 25900
rect 93262 25844 93318 25900
rect 93366 25844 93422 25900
rect 93470 25844 93526 25900
rect 130082 25844 130138 25900
rect 130186 25844 130242 25900
rect 130290 25844 130346 25900
rect 38032 25060 38088 25116
rect 38136 25060 38192 25116
rect 38240 25060 38296 25116
rect 74852 25060 74908 25116
rect 74956 25060 75012 25116
rect 75060 25060 75116 25116
rect 111672 25060 111728 25116
rect 111776 25060 111832 25116
rect 111880 25060 111936 25116
rect 148492 25060 148548 25116
rect 148596 25060 148652 25116
rect 148700 25060 148756 25116
rect 19622 24276 19678 24332
rect 19726 24276 19782 24332
rect 19830 24276 19886 24332
rect 56442 24276 56498 24332
rect 56546 24276 56602 24332
rect 56650 24276 56706 24332
rect 93262 24276 93318 24332
rect 93366 24276 93422 24332
rect 93470 24276 93526 24332
rect 130082 24276 130138 24332
rect 130186 24276 130242 24332
rect 130290 24276 130346 24332
rect 38032 23492 38088 23548
rect 38136 23492 38192 23548
rect 38240 23492 38296 23548
rect 74852 23492 74908 23548
rect 74956 23492 75012 23548
rect 75060 23492 75116 23548
rect 111672 23492 111728 23548
rect 111776 23492 111832 23548
rect 111880 23492 111936 23548
rect 148492 23492 148548 23548
rect 148596 23492 148652 23548
rect 148700 23492 148756 23548
rect 19622 22708 19678 22764
rect 19726 22708 19782 22764
rect 19830 22708 19886 22764
rect 56442 22708 56498 22764
rect 56546 22708 56602 22764
rect 56650 22708 56706 22764
rect 93262 22708 93318 22764
rect 93366 22708 93422 22764
rect 93470 22708 93526 22764
rect 130082 22708 130138 22764
rect 130186 22708 130242 22764
rect 130290 22708 130346 22764
rect 38032 21924 38088 21980
rect 38136 21924 38192 21980
rect 38240 21924 38296 21980
rect 74852 21924 74908 21980
rect 74956 21924 75012 21980
rect 75060 21924 75116 21980
rect 111672 21924 111728 21980
rect 111776 21924 111832 21980
rect 111880 21924 111936 21980
rect 148492 21924 148548 21980
rect 148596 21924 148652 21980
rect 148700 21924 148756 21980
rect 19622 21140 19678 21196
rect 19726 21140 19782 21196
rect 19830 21140 19886 21196
rect 56442 21140 56498 21196
rect 56546 21140 56602 21196
rect 56650 21140 56706 21196
rect 93262 21140 93318 21196
rect 93366 21140 93422 21196
rect 93470 21140 93526 21196
rect 130082 21140 130138 21196
rect 130186 21140 130242 21196
rect 130290 21140 130346 21196
rect 38032 20356 38088 20412
rect 38136 20356 38192 20412
rect 38240 20356 38296 20412
rect 74852 20356 74908 20412
rect 74956 20356 75012 20412
rect 75060 20356 75116 20412
rect 111672 20356 111728 20412
rect 111776 20356 111832 20412
rect 111880 20356 111936 20412
rect 148492 20356 148548 20412
rect 148596 20356 148652 20412
rect 148700 20356 148756 20412
rect 19622 19572 19678 19628
rect 19726 19572 19782 19628
rect 19830 19572 19886 19628
rect 56442 19572 56498 19628
rect 56546 19572 56602 19628
rect 56650 19572 56706 19628
rect 93262 19572 93318 19628
rect 93366 19572 93422 19628
rect 93470 19572 93526 19628
rect 130082 19572 130138 19628
rect 130186 19572 130242 19628
rect 130290 19572 130346 19628
rect 38032 18788 38088 18844
rect 38136 18788 38192 18844
rect 38240 18788 38296 18844
rect 74852 18788 74908 18844
rect 74956 18788 75012 18844
rect 75060 18788 75116 18844
rect 111672 18788 111728 18844
rect 111776 18788 111832 18844
rect 111880 18788 111936 18844
rect 148492 18788 148548 18844
rect 148596 18788 148652 18844
rect 148700 18788 148756 18844
rect 19622 18004 19678 18060
rect 19726 18004 19782 18060
rect 19830 18004 19886 18060
rect 56442 18004 56498 18060
rect 56546 18004 56602 18060
rect 56650 18004 56706 18060
rect 93262 18004 93318 18060
rect 93366 18004 93422 18060
rect 93470 18004 93526 18060
rect 130082 18004 130138 18060
rect 130186 18004 130242 18060
rect 130290 18004 130346 18060
rect 38032 17220 38088 17276
rect 38136 17220 38192 17276
rect 38240 17220 38296 17276
rect 74852 17220 74908 17276
rect 74956 17220 75012 17276
rect 75060 17220 75116 17276
rect 111672 17220 111728 17276
rect 111776 17220 111832 17276
rect 111880 17220 111936 17276
rect 148492 17220 148548 17276
rect 148596 17220 148652 17276
rect 148700 17220 148756 17276
rect 19622 16436 19678 16492
rect 19726 16436 19782 16492
rect 19830 16436 19886 16492
rect 56442 16436 56498 16492
rect 56546 16436 56602 16492
rect 56650 16436 56706 16492
rect 93262 16436 93318 16492
rect 93366 16436 93422 16492
rect 93470 16436 93526 16492
rect 130082 16436 130138 16492
rect 130186 16436 130242 16492
rect 130290 16436 130346 16492
rect 38032 15652 38088 15708
rect 38136 15652 38192 15708
rect 38240 15652 38296 15708
rect 74852 15652 74908 15708
rect 74956 15652 75012 15708
rect 75060 15652 75116 15708
rect 111672 15652 111728 15708
rect 111776 15652 111832 15708
rect 111880 15652 111936 15708
rect 148492 15652 148548 15708
rect 148596 15652 148652 15708
rect 148700 15652 148756 15708
rect 19622 14868 19678 14924
rect 19726 14868 19782 14924
rect 19830 14868 19886 14924
rect 56442 14868 56498 14924
rect 56546 14868 56602 14924
rect 56650 14868 56706 14924
rect 93262 14868 93318 14924
rect 93366 14868 93422 14924
rect 93470 14868 93526 14924
rect 130082 14868 130138 14924
rect 130186 14868 130242 14924
rect 130290 14868 130346 14924
rect 38032 14084 38088 14140
rect 38136 14084 38192 14140
rect 38240 14084 38296 14140
rect 74852 14084 74908 14140
rect 74956 14084 75012 14140
rect 75060 14084 75116 14140
rect 111672 14084 111728 14140
rect 111776 14084 111832 14140
rect 111880 14084 111936 14140
rect 148492 14084 148548 14140
rect 148596 14084 148652 14140
rect 148700 14084 148756 14140
rect 19622 13300 19678 13356
rect 19726 13300 19782 13356
rect 19830 13300 19886 13356
rect 56442 13300 56498 13356
rect 56546 13300 56602 13356
rect 56650 13300 56706 13356
rect 93262 13300 93318 13356
rect 93366 13300 93422 13356
rect 93470 13300 93526 13356
rect 130082 13300 130138 13356
rect 130186 13300 130242 13356
rect 130290 13300 130346 13356
rect 38032 12516 38088 12572
rect 38136 12516 38192 12572
rect 38240 12516 38296 12572
rect 74852 12516 74908 12572
rect 74956 12516 75012 12572
rect 75060 12516 75116 12572
rect 111672 12516 111728 12572
rect 111776 12516 111832 12572
rect 111880 12516 111936 12572
rect 148492 12516 148548 12572
rect 148596 12516 148652 12572
rect 148700 12516 148756 12572
rect 19622 11732 19678 11788
rect 19726 11732 19782 11788
rect 19830 11732 19886 11788
rect 56442 11732 56498 11788
rect 56546 11732 56602 11788
rect 56650 11732 56706 11788
rect 93262 11732 93318 11788
rect 93366 11732 93422 11788
rect 93470 11732 93526 11788
rect 130082 11732 130138 11788
rect 130186 11732 130242 11788
rect 130290 11732 130346 11788
rect 38032 10948 38088 11004
rect 38136 10948 38192 11004
rect 38240 10948 38296 11004
rect 74852 10948 74908 11004
rect 74956 10948 75012 11004
rect 75060 10948 75116 11004
rect 111672 10948 111728 11004
rect 111776 10948 111832 11004
rect 111880 10948 111936 11004
rect 148492 10948 148548 11004
rect 148596 10948 148652 11004
rect 148700 10948 148756 11004
rect 19622 10164 19678 10220
rect 19726 10164 19782 10220
rect 19830 10164 19886 10220
rect 56442 10164 56498 10220
rect 56546 10164 56602 10220
rect 56650 10164 56706 10220
rect 93262 10164 93318 10220
rect 93366 10164 93422 10220
rect 93470 10164 93526 10220
rect 130082 10164 130138 10220
rect 130186 10164 130242 10220
rect 130290 10164 130346 10220
rect 38032 9380 38088 9436
rect 38136 9380 38192 9436
rect 38240 9380 38296 9436
rect 74852 9380 74908 9436
rect 74956 9380 75012 9436
rect 75060 9380 75116 9436
rect 111672 9380 111728 9436
rect 111776 9380 111832 9436
rect 111880 9380 111936 9436
rect 148492 9380 148548 9436
rect 148596 9380 148652 9436
rect 148700 9380 148756 9436
rect 19622 8596 19678 8652
rect 19726 8596 19782 8652
rect 19830 8596 19886 8652
rect 56442 8596 56498 8652
rect 56546 8596 56602 8652
rect 56650 8596 56706 8652
rect 93262 8596 93318 8652
rect 93366 8596 93422 8652
rect 93470 8596 93526 8652
rect 130082 8596 130138 8652
rect 130186 8596 130242 8652
rect 130290 8596 130346 8652
rect 38032 7812 38088 7868
rect 38136 7812 38192 7868
rect 38240 7812 38296 7868
rect 74852 7812 74908 7868
rect 74956 7812 75012 7868
rect 75060 7812 75116 7868
rect 111672 7812 111728 7868
rect 111776 7812 111832 7868
rect 111880 7812 111936 7868
rect 148492 7812 148548 7868
rect 148596 7812 148652 7868
rect 148700 7812 148756 7868
rect 19622 7028 19678 7084
rect 19726 7028 19782 7084
rect 19830 7028 19886 7084
rect 56442 7028 56498 7084
rect 56546 7028 56602 7084
rect 56650 7028 56706 7084
rect 93262 7028 93318 7084
rect 93366 7028 93422 7084
rect 93470 7028 93526 7084
rect 130082 7028 130138 7084
rect 130186 7028 130242 7084
rect 130290 7028 130346 7084
rect 38032 6244 38088 6300
rect 38136 6244 38192 6300
rect 38240 6244 38296 6300
rect 74852 6244 74908 6300
rect 74956 6244 75012 6300
rect 75060 6244 75116 6300
rect 111672 6244 111728 6300
rect 111776 6244 111832 6300
rect 111880 6244 111936 6300
rect 148492 6244 148548 6300
rect 148596 6244 148652 6300
rect 148700 6244 148756 6300
rect 19622 5460 19678 5516
rect 19726 5460 19782 5516
rect 19830 5460 19886 5516
rect 56442 5460 56498 5516
rect 56546 5460 56602 5516
rect 56650 5460 56706 5516
rect 93262 5460 93318 5516
rect 93366 5460 93422 5516
rect 93470 5460 93526 5516
rect 130082 5460 130138 5516
rect 130186 5460 130242 5516
rect 130290 5460 130346 5516
rect 38032 4676 38088 4732
rect 38136 4676 38192 4732
rect 38240 4676 38296 4732
rect 74852 4676 74908 4732
rect 74956 4676 75012 4732
rect 75060 4676 75116 4732
rect 111672 4676 111728 4732
rect 111776 4676 111832 4732
rect 111880 4676 111936 4732
rect 148492 4676 148548 4732
rect 148596 4676 148652 4732
rect 148700 4676 148756 4732
rect 19622 3892 19678 3948
rect 19726 3892 19782 3948
rect 19830 3892 19886 3948
rect 56442 3892 56498 3948
rect 56546 3892 56602 3948
rect 56650 3892 56706 3948
rect 93262 3892 93318 3948
rect 93366 3892 93422 3948
rect 93470 3892 93526 3948
rect 130082 3892 130138 3948
rect 130186 3892 130242 3948
rect 130290 3892 130346 3948
rect 114156 3500 114212 3556
rect 114156 3276 114212 3332
rect 38032 3108 38088 3164
rect 38136 3108 38192 3164
rect 38240 3108 38296 3164
rect 74852 3108 74908 3164
rect 74956 3108 75012 3164
rect 75060 3108 75116 3164
rect 111672 3108 111728 3164
rect 111776 3108 111832 3164
rect 111880 3108 111936 3164
rect 148492 3108 148548 3164
rect 148596 3108 148652 3164
rect 148700 3108 148756 3164
rect 117852 1148 117908 1204
rect 117852 700 117908 756
<< metal4 >>
rect 19594 36876 19914 36908
rect 19594 36820 19622 36876
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19886 36820 19914 36876
rect 19594 35308 19914 36820
rect 19594 35252 19622 35308
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19886 35252 19914 35308
rect 19594 33740 19914 35252
rect 19594 33684 19622 33740
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19886 33684 19914 33740
rect 19594 32172 19914 33684
rect 19594 32116 19622 32172
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19886 32116 19914 32172
rect 19594 30604 19914 32116
rect 19594 30548 19622 30604
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19886 30548 19914 30604
rect 19594 29036 19914 30548
rect 19594 28980 19622 29036
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19886 28980 19914 29036
rect 19594 27468 19914 28980
rect 19594 27412 19622 27468
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19886 27412 19914 27468
rect 19594 25900 19914 27412
rect 19594 25844 19622 25900
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19886 25844 19914 25900
rect 19594 24332 19914 25844
rect 19594 24276 19622 24332
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19886 24276 19914 24332
rect 19594 22764 19914 24276
rect 19594 22708 19622 22764
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19886 22708 19914 22764
rect 19594 21196 19914 22708
rect 19594 21140 19622 21196
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19886 21140 19914 21196
rect 19594 19628 19914 21140
rect 19594 19572 19622 19628
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19886 19572 19914 19628
rect 19594 18060 19914 19572
rect 19594 18004 19622 18060
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19886 18004 19914 18060
rect 19594 16492 19914 18004
rect 19594 16436 19622 16492
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19886 16436 19914 16492
rect 19594 14924 19914 16436
rect 19594 14868 19622 14924
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19886 14868 19914 14924
rect 19594 13356 19914 14868
rect 19594 13300 19622 13356
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19886 13300 19914 13356
rect 19594 11788 19914 13300
rect 19594 11732 19622 11788
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19886 11732 19914 11788
rect 19594 10220 19914 11732
rect 19594 10164 19622 10220
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19886 10164 19914 10220
rect 19594 8652 19914 10164
rect 19594 8596 19622 8652
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19886 8596 19914 8652
rect 19594 7084 19914 8596
rect 19594 7028 19622 7084
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19886 7028 19914 7084
rect 19594 5516 19914 7028
rect 19594 5460 19622 5516
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19886 5460 19914 5516
rect 19594 3948 19914 5460
rect 19594 3892 19622 3948
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19886 3892 19914 3948
rect 19594 3076 19914 3892
rect 38004 36092 38324 36908
rect 38004 36036 38032 36092
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38296 36036 38324 36092
rect 38004 34524 38324 36036
rect 38004 34468 38032 34524
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38296 34468 38324 34524
rect 38004 32956 38324 34468
rect 38004 32900 38032 32956
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38296 32900 38324 32956
rect 38004 31388 38324 32900
rect 38004 31332 38032 31388
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38296 31332 38324 31388
rect 38004 29820 38324 31332
rect 38004 29764 38032 29820
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38296 29764 38324 29820
rect 38004 28252 38324 29764
rect 38004 28196 38032 28252
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38296 28196 38324 28252
rect 38004 26684 38324 28196
rect 38004 26628 38032 26684
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38296 26628 38324 26684
rect 38004 25116 38324 26628
rect 38004 25060 38032 25116
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38296 25060 38324 25116
rect 38004 23548 38324 25060
rect 38004 23492 38032 23548
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38296 23492 38324 23548
rect 38004 21980 38324 23492
rect 38004 21924 38032 21980
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38296 21924 38324 21980
rect 38004 20412 38324 21924
rect 38004 20356 38032 20412
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38296 20356 38324 20412
rect 38004 18844 38324 20356
rect 38004 18788 38032 18844
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38296 18788 38324 18844
rect 38004 17276 38324 18788
rect 38004 17220 38032 17276
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38296 17220 38324 17276
rect 38004 15708 38324 17220
rect 38004 15652 38032 15708
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38296 15652 38324 15708
rect 38004 14140 38324 15652
rect 38004 14084 38032 14140
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38296 14084 38324 14140
rect 38004 12572 38324 14084
rect 38004 12516 38032 12572
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38296 12516 38324 12572
rect 38004 11004 38324 12516
rect 38004 10948 38032 11004
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38296 10948 38324 11004
rect 38004 9436 38324 10948
rect 38004 9380 38032 9436
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38296 9380 38324 9436
rect 38004 7868 38324 9380
rect 38004 7812 38032 7868
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38296 7812 38324 7868
rect 38004 6300 38324 7812
rect 38004 6244 38032 6300
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38296 6244 38324 6300
rect 38004 4732 38324 6244
rect 38004 4676 38032 4732
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38296 4676 38324 4732
rect 38004 3164 38324 4676
rect 38004 3108 38032 3164
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38296 3108 38324 3164
rect 38004 3076 38324 3108
rect 56414 36876 56734 36908
rect 56414 36820 56442 36876
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56706 36820 56734 36876
rect 56414 35308 56734 36820
rect 56414 35252 56442 35308
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56706 35252 56734 35308
rect 56414 33740 56734 35252
rect 56414 33684 56442 33740
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56706 33684 56734 33740
rect 56414 32172 56734 33684
rect 56414 32116 56442 32172
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56706 32116 56734 32172
rect 56414 30604 56734 32116
rect 56414 30548 56442 30604
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56706 30548 56734 30604
rect 56414 29036 56734 30548
rect 56414 28980 56442 29036
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56706 28980 56734 29036
rect 56414 27468 56734 28980
rect 56414 27412 56442 27468
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56706 27412 56734 27468
rect 56414 25900 56734 27412
rect 56414 25844 56442 25900
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56706 25844 56734 25900
rect 56414 24332 56734 25844
rect 56414 24276 56442 24332
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56706 24276 56734 24332
rect 56414 22764 56734 24276
rect 56414 22708 56442 22764
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56706 22708 56734 22764
rect 56414 21196 56734 22708
rect 56414 21140 56442 21196
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56706 21140 56734 21196
rect 56414 19628 56734 21140
rect 56414 19572 56442 19628
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56706 19572 56734 19628
rect 56414 18060 56734 19572
rect 56414 18004 56442 18060
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56706 18004 56734 18060
rect 56414 16492 56734 18004
rect 56414 16436 56442 16492
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56706 16436 56734 16492
rect 56414 14924 56734 16436
rect 56414 14868 56442 14924
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56706 14868 56734 14924
rect 56414 13356 56734 14868
rect 56414 13300 56442 13356
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56706 13300 56734 13356
rect 56414 11788 56734 13300
rect 56414 11732 56442 11788
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56706 11732 56734 11788
rect 56414 10220 56734 11732
rect 56414 10164 56442 10220
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56706 10164 56734 10220
rect 56414 8652 56734 10164
rect 56414 8596 56442 8652
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56706 8596 56734 8652
rect 56414 7084 56734 8596
rect 56414 7028 56442 7084
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56706 7028 56734 7084
rect 56414 5516 56734 7028
rect 56414 5460 56442 5516
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56706 5460 56734 5516
rect 56414 3948 56734 5460
rect 56414 3892 56442 3948
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56706 3892 56734 3948
rect 56414 3076 56734 3892
rect 74824 36092 75144 36908
rect 74824 36036 74852 36092
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 75116 36036 75144 36092
rect 74824 34524 75144 36036
rect 74824 34468 74852 34524
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 75116 34468 75144 34524
rect 74824 32956 75144 34468
rect 74824 32900 74852 32956
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 75116 32900 75144 32956
rect 74824 31388 75144 32900
rect 74824 31332 74852 31388
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 75116 31332 75144 31388
rect 74824 29820 75144 31332
rect 74824 29764 74852 29820
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 75116 29764 75144 29820
rect 74824 28252 75144 29764
rect 74824 28196 74852 28252
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 75116 28196 75144 28252
rect 74824 26684 75144 28196
rect 74824 26628 74852 26684
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 75116 26628 75144 26684
rect 74824 25116 75144 26628
rect 74824 25060 74852 25116
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 75116 25060 75144 25116
rect 74824 23548 75144 25060
rect 74824 23492 74852 23548
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 75116 23492 75144 23548
rect 74824 21980 75144 23492
rect 74824 21924 74852 21980
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 75116 21924 75144 21980
rect 74824 20412 75144 21924
rect 74824 20356 74852 20412
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 75116 20356 75144 20412
rect 74824 18844 75144 20356
rect 74824 18788 74852 18844
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 75116 18788 75144 18844
rect 74824 17276 75144 18788
rect 74824 17220 74852 17276
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 75116 17220 75144 17276
rect 74824 15708 75144 17220
rect 74824 15652 74852 15708
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 75116 15652 75144 15708
rect 74824 14140 75144 15652
rect 74824 14084 74852 14140
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 75116 14084 75144 14140
rect 74824 12572 75144 14084
rect 74824 12516 74852 12572
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 75116 12516 75144 12572
rect 74824 11004 75144 12516
rect 74824 10948 74852 11004
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 75116 10948 75144 11004
rect 74824 9436 75144 10948
rect 74824 9380 74852 9436
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 75116 9380 75144 9436
rect 74824 7868 75144 9380
rect 74824 7812 74852 7868
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 75116 7812 75144 7868
rect 74824 6300 75144 7812
rect 74824 6244 74852 6300
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 75116 6244 75144 6300
rect 74824 4732 75144 6244
rect 74824 4676 74852 4732
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 75116 4676 75144 4732
rect 74824 3164 75144 4676
rect 74824 3108 74852 3164
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 75116 3108 75144 3164
rect 74824 3076 75144 3108
rect 93234 36876 93554 36908
rect 93234 36820 93262 36876
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93526 36820 93554 36876
rect 93234 35308 93554 36820
rect 93234 35252 93262 35308
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93526 35252 93554 35308
rect 93234 33740 93554 35252
rect 93234 33684 93262 33740
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93526 33684 93554 33740
rect 93234 32172 93554 33684
rect 93234 32116 93262 32172
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93526 32116 93554 32172
rect 93234 30604 93554 32116
rect 93234 30548 93262 30604
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93526 30548 93554 30604
rect 93234 29036 93554 30548
rect 93234 28980 93262 29036
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93526 28980 93554 29036
rect 93234 27468 93554 28980
rect 93234 27412 93262 27468
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93526 27412 93554 27468
rect 93234 25900 93554 27412
rect 93234 25844 93262 25900
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93526 25844 93554 25900
rect 93234 24332 93554 25844
rect 93234 24276 93262 24332
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93526 24276 93554 24332
rect 93234 22764 93554 24276
rect 93234 22708 93262 22764
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93526 22708 93554 22764
rect 93234 21196 93554 22708
rect 93234 21140 93262 21196
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93526 21140 93554 21196
rect 93234 19628 93554 21140
rect 93234 19572 93262 19628
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93526 19572 93554 19628
rect 93234 18060 93554 19572
rect 93234 18004 93262 18060
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93526 18004 93554 18060
rect 93234 16492 93554 18004
rect 93234 16436 93262 16492
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93526 16436 93554 16492
rect 93234 14924 93554 16436
rect 93234 14868 93262 14924
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93526 14868 93554 14924
rect 93234 13356 93554 14868
rect 93234 13300 93262 13356
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93526 13300 93554 13356
rect 93234 11788 93554 13300
rect 93234 11732 93262 11788
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93526 11732 93554 11788
rect 93234 10220 93554 11732
rect 93234 10164 93262 10220
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93526 10164 93554 10220
rect 93234 8652 93554 10164
rect 93234 8596 93262 8652
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93526 8596 93554 8652
rect 93234 7084 93554 8596
rect 93234 7028 93262 7084
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93526 7028 93554 7084
rect 93234 5516 93554 7028
rect 93234 5460 93262 5516
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93526 5460 93554 5516
rect 93234 3948 93554 5460
rect 93234 3892 93262 3948
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93526 3892 93554 3948
rect 93234 3076 93554 3892
rect 111644 36092 111964 36908
rect 111644 36036 111672 36092
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111936 36036 111964 36092
rect 111644 34524 111964 36036
rect 111644 34468 111672 34524
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111936 34468 111964 34524
rect 111644 32956 111964 34468
rect 111644 32900 111672 32956
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111936 32900 111964 32956
rect 111644 31388 111964 32900
rect 111644 31332 111672 31388
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111936 31332 111964 31388
rect 111644 29820 111964 31332
rect 111644 29764 111672 29820
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111936 29764 111964 29820
rect 111644 28252 111964 29764
rect 111644 28196 111672 28252
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111936 28196 111964 28252
rect 111644 26684 111964 28196
rect 111644 26628 111672 26684
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111936 26628 111964 26684
rect 111644 25116 111964 26628
rect 111644 25060 111672 25116
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111936 25060 111964 25116
rect 111644 23548 111964 25060
rect 111644 23492 111672 23548
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111936 23492 111964 23548
rect 111644 21980 111964 23492
rect 111644 21924 111672 21980
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111936 21924 111964 21980
rect 111644 20412 111964 21924
rect 111644 20356 111672 20412
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111936 20356 111964 20412
rect 111644 18844 111964 20356
rect 111644 18788 111672 18844
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111936 18788 111964 18844
rect 111644 17276 111964 18788
rect 111644 17220 111672 17276
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111936 17220 111964 17276
rect 111644 15708 111964 17220
rect 111644 15652 111672 15708
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111936 15652 111964 15708
rect 111644 14140 111964 15652
rect 111644 14084 111672 14140
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111936 14084 111964 14140
rect 111644 12572 111964 14084
rect 111644 12516 111672 12572
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111936 12516 111964 12572
rect 111644 11004 111964 12516
rect 111644 10948 111672 11004
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111936 10948 111964 11004
rect 111644 9436 111964 10948
rect 111644 9380 111672 9436
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111936 9380 111964 9436
rect 111644 7868 111964 9380
rect 111644 7812 111672 7868
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111936 7812 111964 7868
rect 111644 6300 111964 7812
rect 111644 6244 111672 6300
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111936 6244 111964 6300
rect 111644 4732 111964 6244
rect 111644 4676 111672 4732
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111936 4676 111964 4732
rect 111644 3164 111964 4676
rect 130054 36876 130374 36908
rect 130054 36820 130082 36876
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130346 36820 130374 36876
rect 130054 35308 130374 36820
rect 130054 35252 130082 35308
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130346 35252 130374 35308
rect 130054 33740 130374 35252
rect 130054 33684 130082 33740
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130346 33684 130374 33740
rect 130054 32172 130374 33684
rect 130054 32116 130082 32172
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130346 32116 130374 32172
rect 130054 30604 130374 32116
rect 130054 30548 130082 30604
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130346 30548 130374 30604
rect 130054 29036 130374 30548
rect 130054 28980 130082 29036
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130346 28980 130374 29036
rect 130054 27468 130374 28980
rect 130054 27412 130082 27468
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130346 27412 130374 27468
rect 130054 25900 130374 27412
rect 130054 25844 130082 25900
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130346 25844 130374 25900
rect 130054 24332 130374 25844
rect 130054 24276 130082 24332
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130346 24276 130374 24332
rect 130054 22764 130374 24276
rect 130054 22708 130082 22764
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130346 22708 130374 22764
rect 130054 21196 130374 22708
rect 130054 21140 130082 21196
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130346 21140 130374 21196
rect 130054 19628 130374 21140
rect 130054 19572 130082 19628
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130346 19572 130374 19628
rect 130054 18060 130374 19572
rect 130054 18004 130082 18060
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130346 18004 130374 18060
rect 130054 16492 130374 18004
rect 130054 16436 130082 16492
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130346 16436 130374 16492
rect 130054 14924 130374 16436
rect 130054 14868 130082 14924
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130346 14868 130374 14924
rect 130054 13356 130374 14868
rect 130054 13300 130082 13356
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130346 13300 130374 13356
rect 130054 11788 130374 13300
rect 130054 11732 130082 11788
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130346 11732 130374 11788
rect 130054 10220 130374 11732
rect 130054 10164 130082 10220
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130346 10164 130374 10220
rect 130054 8652 130374 10164
rect 130054 8596 130082 8652
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130346 8596 130374 8652
rect 130054 7084 130374 8596
rect 130054 7028 130082 7084
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130346 7028 130374 7084
rect 130054 5516 130374 7028
rect 130054 5460 130082 5516
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130346 5460 130374 5516
rect 130054 3948 130374 5460
rect 130054 3892 130082 3948
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130346 3892 130374 3948
rect 114156 3556 114212 3566
rect 114156 3332 114212 3500
rect 114156 3266 114212 3276
rect 111644 3108 111672 3164
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111936 3108 111964 3164
rect 111644 3076 111964 3108
rect 130054 3076 130374 3892
rect 148464 36092 148784 36908
rect 148464 36036 148492 36092
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148756 36036 148784 36092
rect 148464 34524 148784 36036
rect 148464 34468 148492 34524
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148756 34468 148784 34524
rect 148464 32956 148784 34468
rect 148464 32900 148492 32956
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148756 32900 148784 32956
rect 148464 31388 148784 32900
rect 148464 31332 148492 31388
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148756 31332 148784 31388
rect 148464 29820 148784 31332
rect 148464 29764 148492 29820
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148756 29764 148784 29820
rect 148464 28252 148784 29764
rect 148464 28196 148492 28252
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148756 28196 148784 28252
rect 148464 26684 148784 28196
rect 148464 26628 148492 26684
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148756 26628 148784 26684
rect 148464 25116 148784 26628
rect 148464 25060 148492 25116
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148756 25060 148784 25116
rect 148464 23548 148784 25060
rect 148464 23492 148492 23548
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148756 23492 148784 23548
rect 148464 21980 148784 23492
rect 148464 21924 148492 21980
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148756 21924 148784 21980
rect 148464 20412 148784 21924
rect 148464 20356 148492 20412
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148756 20356 148784 20412
rect 148464 18844 148784 20356
rect 148464 18788 148492 18844
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148756 18788 148784 18844
rect 148464 17276 148784 18788
rect 148464 17220 148492 17276
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148756 17220 148784 17276
rect 148464 15708 148784 17220
rect 148464 15652 148492 15708
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148756 15652 148784 15708
rect 148464 14140 148784 15652
rect 148464 14084 148492 14140
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148756 14084 148784 14140
rect 148464 12572 148784 14084
rect 148464 12516 148492 12572
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148756 12516 148784 12572
rect 148464 11004 148784 12516
rect 148464 10948 148492 11004
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148756 10948 148784 11004
rect 148464 9436 148784 10948
rect 148464 9380 148492 9436
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148756 9380 148784 9436
rect 148464 7868 148784 9380
rect 148464 7812 148492 7868
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148756 7812 148784 7868
rect 148464 6300 148784 7812
rect 148464 6244 148492 6300
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148756 6244 148784 6300
rect 148464 4732 148784 6244
rect 148464 4676 148492 4732
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148756 4676 148784 4732
rect 148464 3164 148784 4676
rect 148464 3108 148492 3164
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148756 3108 148784 3164
rect 148464 3076 148784 3108
rect 117852 1204 117908 1214
rect 117852 756 117908 1148
rect 117852 690 117908 700
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__042__I dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 135296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__043__I
timestamp 1666464484
transform 1 0 130480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__044__I0
timestamp 1666464484
transform 1 0 121408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__046__I0
timestamp 1666464484
transform 1 0 126000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__048__I0
timestamp 1666464484
transform -1 0 123984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__050__I0
timestamp 1666464484
transform -1 0 126672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__052__I
timestamp 1666464484
transform 1 0 132048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__053__I0
timestamp 1666464484
transform -1 0 128688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__055__I0
timestamp 1666464484
transform -1 0 129360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__057__I0
timestamp 1666464484
transform -1 0 131040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I0
timestamp 1666464484
transform -1 0 132048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__061__I
timestamp 1666464484
transform 1 0 135520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__062__I0
timestamp 1666464484
transform -1 0 136192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I0
timestamp 1666464484
transform -1 0 136864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__066__I0
timestamp 1666464484
transform -1 0 138880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__I0
timestamp 1666464484
transform -1 0 138768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__I
timestamp 1666464484
transform 1 0 134624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I0
timestamp 1666464484
transform 1 0 144816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__S
timestamp 1666464484
transform 1 0 143472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__I0
timestamp 1666464484
transform -1 0 140336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__S
timestamp 1666464484
transform 1 0 139888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__I0
timestamp 1666464484
transform -1 0 139664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__S
timestamp 1666464484
transform -1 0 141008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I0
timestamp 1666464484
transform 1 0 114912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I1
timestamp 1666464484
transform 1 0 113568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__S
timestamp 1666464484
transform 1 0 115360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__I
timestamp 1666464484
transform 1 0 127568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__I
timestamp 1666464484
transform 1 0 103040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I0
timestamp 1666464484
transform -1 0 98112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__083__I0
timestamp 1666464484
transform 1 0 97104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__I0
timestamp 1666464484
transform -1 0 99680 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__I
timestamp 1666464484
transform 1 0 101136 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__I0
timestamp 1666464484
transform -1 0 100464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__I
timestamp 1666464484
transform 1 0 104384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I0
timestamp 1666464484
transform -1 0 101696 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__I0
timestamp 1666464484
transform -1 0 103600 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__I0
timestamp 1666464484
transform -1 0 103040 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__I0
timestamp 1666464484
transform 1 0 106960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__I
timestamp 1666464484
transform -1 0 111664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__I0
timestamp 1666464484
transform -1 0 109088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__I0
timestamp 1666464484
transform -1 0 110320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__I
timestamp 1666464484
transform 1 0 113120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__I0
timestamp 1666464484
transform 1 0 112112 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__I0
timestamp 1666464484
transform -1 0 109648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__I
timestamp 1666464484
transform 1 0 117824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__I0
timestamp 1666464484
transform -1 0 116144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__I0
timestamp 1666464484
transform -1 0 115696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__I0
timestamp 1666464484
transform -1 0 117600 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__I0
timestamp 1666464484
transform -1 0 119280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__I
timestamp 1666464484
transform -1 0 75936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__I
timestamp 1666464484
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__I
timestamp 1666464484
transform 1 0 80416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I
timestamp 1666464484
transform 1 0 81312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__I
timestamp 1666464484
transform -1 0 83664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__I
timestamp 1666464484
transform 1 0 84448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__I
timestamp 1666464484
transform 1 0 86352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I
timestamp 1666464484
transform 1 0 88032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__I
timestamp 1666464484
transform 1 0 89712 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__I
timestamp 1666464484
transform -1 0 77728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__I
timestamp 1666464484
transform -1 0 79520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1666464484
transform 1 0 82096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__I
timestamp 1666464484
transform -1 0 82768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__I
timestamp 1666464484
transform -1 0 85456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__I
timestamp 1666464484
transform 1 0 86912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__I
timestamp 1666464484
transform 1 0 88368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I
timestamp 1666464484
transform 1 0 90160 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__I
timestamp 1666464484
transform -1 0 91392 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__I
timestamp 1666464484
transform 1 0 73920 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__I
timestamp 1666464484
transform 1 0 76048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1666464484
transform -1 0 146496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1666464484
transform -1 0 146496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1666464484
transform -1 0 146048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1666464484
transform -1 0 147392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1666464484
transform -1 0 147392 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1666464484
transform -1 0 147392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1666464484
transform -1 0 147392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1666464484
transform -1 0 147392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1666464484
transform -1 0 147392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1666464484
transform -1 0 147392 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1666464484
transform -1 0 146944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1666464484
transform -1 0 21840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1666464484
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1666464484
transform -1 0 40432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1666464484
transform -1 0 42000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1666464484
transform 1 0 44352 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1666464484
transform -1 0 45360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1666464484
transform -1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1666464484
transform -1 0 48944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1666464484
transform -1 0 50400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1666464484
transform -1 0 52192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1666464484
transform -1 0 53760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1666464484
transform -1 0 23520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1666464484
transform 1 0 56112 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1666464484
transform -1 0 57120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1666464484
transform -1 0 58800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1666464484
transform -1 0 60704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1666464484
transform -1 0 62160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1666464484
transform -1 0 63952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1666464484
transform -1 0 65520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1666464484
transform 1 0 67872 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1666464484
transform -1 0 68880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1666464484
transform -1 0 70560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1666464484
transform 1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1666464484
transform 1 0 73248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1666464484
transform 1 0 74368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1666464484
transform -1 0 26880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1666464484
transform -1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1666464484
transform -1 0 30240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1666464484
transform 1 0 32592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1666464484
transform -1 0 33600 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1666464484
transform -1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1666464484
transform -1 0 37184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1666464484
transform -1 0 93632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1666464484
transform -1 0 108640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1666464484
transform -1 0 113344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1666464484
transform -1 0 114240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1666464484
transform -1 0 114240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1666464484
transform -1 0 117152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1666464484
transform 1 0 118272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1666464484
transform 1 0 120960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1666464484
transform -1 0 121184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1666464484
transform 1 0 122752 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1666464484
transform 1 0 128016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1666464484
transform -1 0 94528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1666464484
transform 1 0 128912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1666464484
transform 1 0 128240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1666464484
transform -1 0 129360 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1666464484
transform -1 0 132944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1666464484
transform -1 0 133840 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1666464484
transform 1 0 135072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1666464484
transform 1 0 138096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1666464484
transform 1 0 141232 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1666464484
transform 1 0 145600 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1666464484
transform 1 0 143024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1666464484
transform -1 0 95984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1666464484
transform 1 0 145264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1666464484
transform 1 0 146048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1666464484
transform 1 0 98336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1666464484
transform -1 0 99120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1666464484
transform -1 0 101248 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1666464484
transform -1 0 102592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1666464484
transform 1 0 107408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1666464484
transform 1 0 107856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1666464484
transform 1 0 108640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output76_I
timestamp 1666464484
transform -1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output77_I
timestamp 1666464484
transform -1 0 9856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output78_I
timestamp 1666464484
transform -1 0 11424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output79_I
timestamp 1666464484
transform 1 0 12992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output80_I
timestamp 1666464484
transform 1 0 15120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output81_I
timestamp 1666464484
transform -1 0 17584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output82_I
timestamp 1666464484
transform 1 0 19376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output83_I
timestamp 1666464484
transform -1 0 20720 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output84_I
timestamp 1666464484
transform 1 0 22960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output94_I
timestamp 1666464484
transform -1 0 6720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output96_I
timestamp 1666464484
transform 1 0 146272 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output97_I
timestamp 1666464484
transform 1 0 146272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output98_I
timestamp 1666464484
transform -1 0 146496 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output99_I
timestamp 1666464484
transform 1 0 146272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output100_I
timestamp 1666464484
transform -1 0 146496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output101_I
timestamp 1666464484
transform 1 0 146272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output102_I
timestamp 1666464484
transform -1 0 146496 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output103_I
timestamp 1666464484
transform 1 0 146272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output104_I
timestamp 1666464484
transform 1 0 146272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output105_I
timestamp 1666464484
transform -1 0 146496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output106_I
timestamp 1666464484
transform 1 0 146272 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output107_I
timestamp 1666464484
transform -1 0 146496 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output108_I
timestamp 1666464484
transform -1 0 146496 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output109_I
timestamp 1666464484
transform 1 0 146272 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output110_I
timestamp 1666464484
transform -1 0 146496 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output111_I
timestamp 1666464484
transform 1 0 146272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output112_I
timestamp 1666464484
transform 1 0 146272 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output113_I
timestamp 1666464484
transform -1 0 146496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output114_I
timestamp 1666464484
transform 1 0 145824 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output115_I
timestamp 1666464484
transform 1 0 145376 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output116_I
timestamp 1666464484
transform 1 0 143808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output117_I
timestamp 1666464484
transform 1 0 144256 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output118_I
timestamp 1666464484
transform 1 0 146272 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output119_I
timestamp 1666464484
transform -1 0 144368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output120_I
timestamp 1666464484
transform 1 0 144480 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output121_I
timestamp 1666464484
transform 1 0 146272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output122_I
timestamp 1666464484
transform -1 0 146496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output123_I
timestamp 1666464484
transform 1 0 146272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output124_I
timestamp 1666464484
transform -1 0 146496 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output125_I
timestamp 1666464484
transform 1 0 146272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output126_I
timestamp 1666464484
transform -1 0 146496 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output127_I
timestamp 1666464484
transform 1 0 146272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1666464484
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 7168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54
timestamp 1666464484
transform 1 0 7392 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1666464484
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72
timestamp 1666464484
transform 1 0 9408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88
timestamp 1666464484
transform 1 0 11200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1666464484
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107
timestamp 1666464484
transform 1 0 13328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123
timestamp 1666464484
transform 1 0 15120 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1666464484
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1666464484
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_145 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 17584 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_153
timestamp 1666464484
transform 1 0 18480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_169
timestamp 1666464484
transform 1 0 20272 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_173
timestamp 1666464484
transform 1 0 20720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1666464484
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 22848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_198
timestamp 1666464484
transform 1 0 23520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_206
timestamp 1666464484
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_212
timestamp 1666464484
transform 1 0 25088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_214
timestamp 1666464484
transform 1 0 25312 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_221
timestamp 1666464484
transform 1 0 26096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_225
timestamp 1666464484
transform 1 0 26544 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_228
timestamp 1666464484
transform 1 0 26880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_236
timestamp 1666464484
transform 1 0 27776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_240
timestamp 1666464484
transform 1 0 28224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1666464484
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1666464484
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_254
timestamp 1666464484
transform 1 0 29792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_258
timestamp 1666464484
transform 1 0 30240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_266
timestamp 1666464484
transform 1 0 31136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_270
timestamp 1666464484
transform 1 0 31584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_272
timestamp 1666464484
transform 1 0 31808 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1666464484
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_282
timestamp 1666464484
transform 1 0 32928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_288
timestamp 1666464484
transform 1 0 33600 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_296
timestamp 1666464484
transform 1 0 34496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_300
timestamp 1666464484
transform 1 0 34944 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_303
timestamp 1666464484
transform 1 0 35280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_311
timestamp 1666464484
transform 1 0 36176 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_317
timestamp 1666464484
transform 1 0 36848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_319
timestamp 1666464484
transform 1 0 37072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_326
timestamp 1666464484
transform 1 0 37856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_330
timestamp 1666464484
transform 1 0 38304 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_333
timestamp 1666464484
transform 1 0 38640 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_341
timestamp 1666464484
transform 1 0 39536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_345
timestamp 1666464484
transform 1 0 39984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1666464484
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1666464484
transform 1 0 40768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_359
timestamp 1666464484
transform 1 0 41552 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_363
timestamp 1666464484
transform 1 0 42000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_371
timestamp 1666464484
transform 1 0 42896 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_375
timestamp 1666464484
transform 1 0 43344 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_377
timestamp 1666464484
transform 1 0 43568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1666464484
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_387
timestamp 1666464484
transform 1 0 44688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_393
timestamp 1666464484
transform 1 0 45360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_401
timestamp 1666464484
transform 1 0 46256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_405
timestamp 1666464484
transform 1 0 46704 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_408
timestamp 1666464484
transform 1 0 47040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_416
timestamp 1666464484
transform 1 0 47936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_422
timestamp 1666464484
transform 1 0 48608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_424
timestamp 1666464484
transform 1 0 48832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_431
timestamp 1666464484
transform 1 0 49616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_435
timestamp 1666464484
transform 1 0 50064 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_438
timestamp 1666464484
transform 1 0 50400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_446
timestamp 1666464484
transform 1 0 51296 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_450
timestamp 1666464484
transform 1 0 51744 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1666464484
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1666464484
transform 1 0 52528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_464
timestamp 1666464484
transform 1 0 53312 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_468
timestamp 1666464484
transform 1 0 53760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_476
timestamp 1666464484
transform 1 0 54656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_480
timestamp 1666464484
transform 1 0 55104 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_482
timestamp 1666464484
transform 1 0 55328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1666464484
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_492
timestamp 1666464484
transform 1 0 56448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_498
timestamp 1666464484
transform 1 0 57120 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_506
timestamp 1666464484
transform 1 0 58016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_510
timestamp 1666464484
transform 1 0 58464 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_513
timestamp 1666464484
transform 1 0 58800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_521
timestamp 1666464484
transform 1 0 59696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_527
timestamp 1666464484
transform 1 0 60368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_529
timestamp 1666464484
transform 1 0 60592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_536
timestamp 1666464484
transform 1 0 61376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_540
timestamp 1666464484
transform 1 0 61824 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_543
timestamp 1666464484
transform 1 0 62160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_551
timestamp 1666464484
transform 1 0 63056 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_555
timestamp 1666464484
transform 1 0 63504 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_559
timestamp 1666464484
transform 1 0 63952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_562
timestamp 1666464484
transform 1 0 64288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_569
timestamp 1666464484
transform 1 0 65072 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_573
timestamp 1666464484
transform 1 0 65520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_581
timestamp 1666464484
transform 1 0 66416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_585
timestamp 1666464484
transform 1 0 66864 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_587
timestamp 1666464484
transform 1 0 67088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_594
timestamp 1666464484
transform 1 0 67872 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_597
timestamp 1666464484
transform 1 0 68208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_603
timestamp 1666464484
transform 1 0 68880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_611
timestamp 1666464484
transform 1 0 69776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_615
timestamp 1666464484
transform 1 0 70224 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_618
timestamp 1666464484
transform 1 0 70560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_626
timestamp 1666464484
transform 1 0 71456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_632
timestamp 1666464484
transform 1 0 72128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_640
timestamp 1666464484
transform 1 0 73024 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_648
timestamp 1666464484
transform 1 0 73920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_656
timestamp 1666464484
transform 1 0 74816 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1666464484
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1666464484
transform 1 0 76048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_682
timestamp 1666464484
transform 1 0 77728 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_698
timestamp 1666464484
transform 1 0 79520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_702
timestamp 1666464484
transform 1 0 79968 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_717
timestamp 1666464484
transform 1 0 81648 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_733
timestamp 1666464484
transform 1 0 83440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_737
timestamp 1666464484
transform 1 0 83888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_739
timestamp 1666464484
transform 1 0 84112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_754
timestamp 1666464484
transform 1 0 85792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_762
timestamp 1666464484
transform 1 0 86688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_766
timestamp 1666464484
transform 1 0 87136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_772
timestamp 1666464484
transform 1 0 87808 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_787
timestamp 1666464484
transform 1 0 89488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_803
timestamp 1666464484
transform 1 0 91280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_807
timestamp 1666464484
transform 1 0 91728 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_822
timestamp 1666464484
transform 1 0 93408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_830
timestamp 1666464484
transform 1 0 94304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_838
timestamp 1666464484
transform 1 0 95200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_842
timestamp 1666464484
transform 1 0 95648 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_844
timestamp 1666464484
transform 1 0 95872 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_851
timestamp 1666464484
transform 1 0 96656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_857
timestamp 1666464484
transform 1 0 97328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_874
timestamp 1666464484
transform 1 0 99232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_877
timestamp 1666464484
transform 1 0 99568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_893
timestamp 1666464484
transform 1 0 101360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_901
timestamp 1666464484
transform 1 0 102256 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_909
timestamp 1666464484
transform 1 0 103152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_912
timestamp 1666464484
transform 1 0 103488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_928
timestamp 1666464484
transform 1 0 105280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_936
timestamp 1666464484
transform 1 0 106176 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_944
timestamp 1666464484
transform 1 0 107072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_947
timestamp 1666464484
transform 1 0 107408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_949
timestamp 1666464484
transform 1 0 107632 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_956
timestamp 1666464484
transform 1 0 108416 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_960
timestamp 1666464484
transform 1 0 108864 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_962
timestamp 1666464484
transform 1 0 109088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_978
timestamp 1666464484
transform 1 0 110880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_982
timestamp 1666464484
transform 1 0 111328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_998
timestamp 1666464484
transform 1 0 113120 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1006
timestamp 1666464484
transform 1 0 114016 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1014
timestamp 1666464484
transform 1 0 114912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1017
timestamp 1666464484
transform 1 0 115248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1033
timestamp 1666464484
transform 1 0 117040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1041
timestamp 1666464484
transform 1 0 117936 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1049
timestamp 1666464484
transform 1 0 118832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1052
timestamp 1666464484
transform 1 0 119168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1068
timestamp 1666464484
transform 1 0 120960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1076
timestamp 1666464484
transform 1 0 121856 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1084
timestamp 1666464484
transform 1 0 122752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1087
timestamp 1666464484
transform 1 0 123088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1103
timestamp 1666464484
transform 1 0 124880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1111
timestamp 1666464484
transform 1 0 125776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1115
timestamp 1666464484
transform 1 0 126224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1119
timestamp 1666464484
transform 1 0 126672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1122
timestamp 1666464484
transform 1 0 127008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1129
timestamp 1666464484
transform 1 0 127792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1133
timestamp 1666464484
transform 1 0 128240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1152
timestamp 1666464484
transform 1 0 130368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1154
timestamp 1666464484
transform 1 0 130592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1157
timestamp 1666464484
transform 1 0 130928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1173
timestamp 1666464484
transform 1 0 132720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1181
timestamp 1666464484
transform 1 0 133616 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1189
timestamp 1666464484
transform 1 0 134512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1192
timestamp 1666464484
transform 1 0 134848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1211
timestamp 1666464484
transform 1 0 136976 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1219
timestamp 1666464484
transform 1 0 137872 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1223
timestamp 1666464484
transform 1 0 138320 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1227
timestamp 1666464484
transform 1 0 138768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1243
timestamp 1666464484
transform 1 0 140560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1251
timestamp 1666464484
transform 1 0 141456 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1259
timestamp 1666464484
transform 1 0 142352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1262
timestamp 1666464484
transform 1 0 142688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1278
timestamp 1666464484
transform 1 0 144480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1286
timestamp 1666464484
transform 1 0 145376 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1290
timestamp 1666464484
transform 1 0 145824 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1294
timestamp 1666464484
transform 1 0 146272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1297
timestamp 1666464484
transform 1 0 146608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1304
timestamp 1666464484
transform 1 0 147392 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1312
timestamp 1666464484
transform 1 0 148288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_2
timestamp 1666464484
transform 1 0 1568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_34
timestamp 1666464484
transform 1 0 5152 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_42
timestamp 1666464484
transform 1 0 6048 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_48
timestamp 1666464484
transform 1 0 6720 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_64
timestamp 1666464484
transform 1 0 8512 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_68
timestamp 1666464484
transform 1 0 8960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1666464484
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1666464484
transform 1 0 9520 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_76
timestamp 1666464484
transform 1 0 9856 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_84
timestamp 1666464484
transform 1 0 10752 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_90
timestamp 1666464484
transform 1 0 11424 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_98
timestamp 1666464484
transform 1 0 12320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_102
timestamp 1666464484
transform 1 0 12768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_106 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 13216 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_122
timestamp 1666464484
transform 1 0 15008 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_125
timestamp 1666464484
transform 1 0 15344 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1666464484
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1666464484
transform 1 0 17472 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_159
timestamp 1666464484
transform 1 0 19152 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_163
timestamp 1666464484
transform 1 0 19600 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_179
timestamp 1666464484
transform 1 0 21392 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_183
timestamp 1666464484
transform 1 0 21840 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_191
timestamp 1666464484
transform 1 0 22736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_195
timestamp 1666464484
transform 1 0 23184 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_211
timestamp 1666464484
transform 1 0 24976 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1666464484
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_218
timestamp 1666464484
transform 1 0 25760 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_250
timestamp 1666464484
transform 1 0 29344 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_266
timestamp 1666464484
transform 1 0 31136 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_274
timestamp 1666464484
transform 1 0 32032 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_278
timestamp 1666464484
transform 1 0 32480 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_281
timestamp 1666464484
transform 1 0 32816 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1666464484
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_286
timestamp 1666464484
transform 1 0 33376 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_320
timestamp 1666464484
transform 1 0 37184 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_352
timestamp 1666464484
transform 1 0 40768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1666464484
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_357
timestamp 1666464484
transform 1 0 41328 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_373
timestamp 1666464484
transform 1 0 43120 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_381
timestamp 1666464484
transform 1 0 44016 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_383
timestamp 1666464484
transform 1 0 44240 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_386
timestamp 1666464484
transform 1 0 44576 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_418
timestamp 1666464484
transform 1 0 48160 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_422
timestamp 1666464484
transform 1 0 48608 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1666464484
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_428
timestamp 1666464484
transform 1 0 49280 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_460
timestamp 1666464484
transform 1 0 52864 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_476
timestamp 1666464484
transform 1 0 54656 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_484
timestamp 1666464484
transform 1 0 55552 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_488
timestamp 1666464484
transform 1 0 56000 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_491
timestamp 1666464484
transform 1 0 56336 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_495
timestamp 1666464484
transform 1 0 56784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_499
timestamp 1666464484
transform 1 0 57232 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_515
timestamp 1666464484
transform 1 0 59024 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_523
timestamp 1666464484
transform 1 0 59920 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_527
timestamp 1666464484
transform 1 0 60368 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_530
timestamp 1666464484
transform 1 0 60704 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_562
timestamp 1666464484
transform 1 0 64288 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_566
timestamp 1666464484
transform 1 0 64736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_570
timestamp 1666464484
transform 1 0 65184 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_586
timestamp 1666464484
transform 1 0 66976 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_596
timestamp 1666464484
transform 1 0 68096 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_628
timestamp 1666464484
transform 1 0 71680 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_636
timestamp 1666464484
transform 1 0 72576 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_638
timestamp 1666464484
transform 1 0 72800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1666464484
transform 1 0 73136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_644
timestamp 1666464484
transform 1 0 73472 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_650
timestamp 1666464484
transform 1 0 74144 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_654
timestamp 1666464484
transform 1 0 74592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_658
timestamp 1666464484
transform 1 0 75040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_665
timestamp 1666464484
transform 1 0 75824 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_669
timestamp 1666464484
transform 1 0 76272 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_673
timestamp 1666464484
transform 1 0 76720 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_680
timestamp 1666464484
transform 1 0 77504 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_688
timestamp 1666464484
transform 1 0 78400 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_696
timestamp 1666464484
transform 1 0 79296 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_704
timestamp 1666464484
transform 1 0 80192 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_708
timestamp 1666464484
transform 1 0 80640 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_712
timestamp 1666464484
transform 1 0 81088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_719
timestamp 1666464484
transform 1 0 81872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_723
timestamp 1666464484
transform 1 0 82320 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_739
timestamp 1666464484
transform 1 0 84112 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_747
timestamp 1666464484
transform 1 0 85008 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_751
timestamp 1666464484
transform 1 0 85456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_769
timestamp 1666464484
transform 1 0 87472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_777
timestamp 1666464484
transform 1 0 88368 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_783
timestamp 1666464484
transform 1 0 89040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_790
timestamp 1666464484
transform 1 0 89824 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_800
timestamp 1666464484
transform 1 0 90944 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_804
timestamp 1666464484
transform 1 0 91392 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_820
timestamp 1666464484
transform 1 0 93184 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_824
timestamp 1666464484
transform 1 0 93632 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_828
timestamp 1666464484
transform 1 0 94080 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_832
timestamp 1666464484
transform 1 0 94528 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_840
timestamp 1666464484
transform 1 0 95424 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_842
timestamp 1666464484
transform 1 0 95648 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_845
timestamp 1666464484
transform 1 0 95984 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_849
timestamp 1666464484
transform 1 0 96432 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_851
timestamp 1666464484
transform 1 0 96656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_854
timestamp 1666464484
transform 1 0 96992 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_862
timestamp 1666464484
transform 1 0 97888 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_879
timestamp 1666464484
transform 1 0 99792 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_896
timestamp 1666464484
transform 1 0 101696 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_913
timestamp 1666464484
transform 1 0 103600 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_921
timestamp 1666464484
transform 1 0 104496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_925
timestamp 1666464484
transform 1 0 104944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_941
timestamp 1666464484
transform 1 0 106736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_945
timestamp 1666464484
transform 1 0 107184 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_949
timestamp 1666464484
transform 1 0 107632 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_953
timestamp 1666464484
transform 1 0 108080 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_955
timestamp 1666464484
transform 1 0 108304 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_958
timestamp 1666464484
transform 1 0 108640 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_962
timestamp 1666464484
transform 1 0 109088 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_970
timestamp 1666464484
transform 1 0 109984 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_987
timestamp 1666464484
transform 1 0 111888 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_991
timestamp 1666464484
transform 1 0 112336 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_993
timestamp 1666464484
transform 1 0 112560 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_996
timestamp 1666464484
transform 1 0 112896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1012
timestamp 1666464484
transform 1 0 114688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1016
timestamp 1666464484
transform 1 0 115136 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1020
timestamp 1666464484
transform 1 0 115584 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1036
timestamp 1666464484
transform 1 0 117376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1053
timestamp 1666464484
transform 1 0 119280 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1061
timestamp 1666464484
transform 1 0 120176 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1067
timestamp 1666464484
transform 1 0 120848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1070
timestamp 1666464484
transform 1 0 121184 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1074
timestamp 1666464484
transform 1 0 121632 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1091
timestamp 1666464484
transform 1 0 123536 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1110
timestamp 1666464484
transform 1 0 125664 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1127
timestamp 1666464484
transform 1 0 127568 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1135
timestamp 1666464484
transform 1 0 128464 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1138
timestamp 1666464484
transform 1 0 128800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1141
timestamp 1666464484
transform 1 0 129136 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1158
timestamp 1666464484
transform 1 0 131040 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1177
timestamp 1666464484
transform 1 0 133168 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1187
timestamp 1666464484
transform 1 0 134288 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1189
timestamp 1666464484
transform 1 0 134512 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1196
timestamp 1666464484
transform 1 0 135296 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1206
timestamp 1666464484
transform 1 0 136416 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1209
timestamp 1666464484
transform 1 0 136752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1225
timestamp 1666464484
transform 1 0 138544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1227
timestamp 1666464484
transform 1 0 138768 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1243
timestamp 1666464484
transform 1 0 140560 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1260
timestamp 1666464484
transform 1 0 142464 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1268
timestamp 1666464484
transform 1 0 143360 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1276
timestamp 1666464484
transform 1 0 144256 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1280
timestamp 1666464484
transform 1 0 144704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1283
timestamp 1666464484
transform 1 0 145040 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1287
timestamp 1666464484
transform 1 0 145488 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1289
timestamp 1666464484
transform 1 0 145712 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1292
timestamp 1666464484
transform 1 0 146048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1296
timestamp 1666464484
transform 1 0 146496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1304
timestamp 1666464484
transform 1 0 147392 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1312
timestamp 1666464484
transform 1 0 148288 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1666464484
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1666464484
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1666464484
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1666464484
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1666464484
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1666464484
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1666464484
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1666464484
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1666464484
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1666464484
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1666464484
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1666464484
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1666464484
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1666464484
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1666464484
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1666464484
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_392
timestamp 1666464484
transform 1 0 45248 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_456
timestamp 1666464484
transform 1 0 52416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1666464484
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_463
timestamp 1666464484
transform 1 0 53200 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_527
timestamp 1666464484
transform 1 0 60368 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1666464484
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_534
timestamp 1666464484
transform 1 0 61152 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_598
timestamp 1666464484
transform 1 0 68320 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_602
timestamp 1666464484
transform 1 0 68768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_605
timestamp 1666464484
transform 1 0 69104 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_637
timestamp 1666464484
transform 1 0 72688 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_653
timestamp 1666464484
transform 1 0 74480 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_661
timestamp 1666464484
transform 1 0 75376 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_663
timestamp 1666464484
transform 1 0 75600 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_666
timestamp 1666464484
transform 1 0 75936 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_676
timestamp 1666464484
transform 1 0 77056 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_682
timestamp 1666464484
transform 1 0 77728 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_686
timestamp 1666464484
transform 1 0 78176 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_690
timestamp 1666464484
transform 1 0 78624 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_694
timestamp 1666464484
transform 1 0 79072 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_698
timestamp 1666464484
transform 1 0 79520 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_712
timestamp 1666464484
transform 1 0 81088 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_716
timestamp 1666464484
transform 1 0 81536 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_718
timestamp 1666464484
transform 1 0 81760 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_725
timestamp 1666464484
transform 1 0 82544 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_733
timestamp 1666464484
transform 1 0 83440 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_735
timestamp 1666464484
transform 1 0 83664 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_742
timestamp 1666464484
transform 1 0 84448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_744
timestamp 1666464484
transform 1 0 84672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_747
timestamp 1666464484
transform 1 0 85008 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_757
timestamp 1666464484
transform 1 0 86128 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_761
timestamp 1666464484
transform 1 0 86576 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_765
timestamp 1666464484
transform 1 0 87024 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_772
timestamp 1666464484
transform 1 0 87808 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_776
timestamp 1666464484
transform 1 0 88256 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_780
timestamp 1666464484
transform 1 0 88704 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_787
timestamp 1666464484
transform 1 0 89488 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_791
timestamp 1666464484
transform 1 0 89936 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_795
timestamp 1666464484
transform 1 0 90384 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_811
timestamp 1666464484
transform 1 0 92176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_815
timestamp 1666464484
transform 1 0 92624 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_818
timestamp 1666464484
transform 1 0 92960 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_850
timestamp 1666464484
transform 1 0 96544 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_858
timestamp 1666464484
transform 1 0 97440 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_864
timestamp 1666464484
transform 1 0 98112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_868
timestamp 1666464484
transform 1 0 98560 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_870
timestamp 1666464484
transform 1 0 98784 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_873
timestamp 1666464484
transform 1 0 99120 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_881
timestamp 1666464484
transform 1 0 100016 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_885
timestamp 1666464484
transform 1 0 100464 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_889
timestamp 1666464484
transform 1 0 100912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_892
timestamp 1666464484
transform 1 0 101248 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_896
timestamp 1666464484
transform 1 0 101696 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_906
timestamp 1666464484
transform 1 0 102816 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_910
timestamp 1666464484
transform 1 0 103264 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_927
timestamp 1666464484
transform 1 0 105168 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_935
timestamp 1666464484
transform 1 0 106064 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_943
timestamp 1666464484
transform 1 0 106960 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_951
timestamp 1666464484
transform 1 0 107856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_955
timestamp 1666464484
transform 1 0 108304 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_957
timestamp 1666464484
transform 1 0 108528 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_960
timestamp 1666464484
transform 1 0 108864 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_964
timestamp 1666464484
transform 1 0 109312 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_967
timestamp 1666464484
transform 1 0 109648 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_975
timestamp 1666464484
transform 1 0 110544 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_992
timestamp 1666464484
transform 1 0 112448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1000
timestamp 1666464484
transform 1 0 113344 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1004
timestamp 1666464484
transform 1 0 113792 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1008
timestamp 1666464484
transform 1 0 114240 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1016
timestamp 1666464484
transform 1 0 115136 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1020
timestamp 1666464484
transform 1 0 115584 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1028
timestamp 1666464484
transform 1 0 116480 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1031
timestamp 1666464484
transform 1 0 116816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1040
timestamp 1666464484
transform 1 0 117824 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1048
timestamp 1666464484
transform 1 0 118720 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1056
timestamp 1666464484
transform 1 0 119616 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1064
timestamp 1666464484
transform 1 0 120512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1070
timestamp 1666464484
transform 1 0 121184 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1078
timestamp 1666464484
transform 1 0 122080 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1082
timestamp 1666464484
transform 1 0 122528 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1086
timestamp 1666464484
transform 1 0 122976 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1096
timestamp 1666464484
transform 1 0 124096 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1102
timestamp 1666464484
transform 1 0 124768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1109
timestamp 1666464484
transform 1 0 125552 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1117
timestamp 1666464484
transform 1 0 126448 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1127
timestamp 1666464484
transform 1 0 127568 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1135
timestamp 1666464484
transform 1 0 128464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1147
timestamp 1666464484
transform 1 0 129808 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1155
timestamp 1666464484
transform 1 0 130704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1165
timestamp 1666464484
transform 1 0 131824 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1169
timestamp 1666464484
transform 1 0 132272 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1173
timestamp 1666464484
transform 1 0 132720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1180
timestamp 1666464484
transform 1 0 133504 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1188
timestamp 1666464484
transform 1 0 134400 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1192
timestamp 1666464484
transform 1 0 134848 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1196
timestamp 1666464484
transform 1 0 135296 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1200
timestamp 1666464484
transform 1 0 135744 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1204
timestamp 1666464484
transform 1 0 136192 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1210
timestamp 1666464484
transform 1 0 136864 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1220
timestamp 1666464484
transform 1 0 137984 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1224
timestamp 1666464484
transform 1 0 138432 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1227
timestamp 1666464484
transform 1 0 138768 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1235
timestamp 1666464484
transform 1 0 139664 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1241
timestamp 1666464484
transform 1 0 140336 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1244
timestamp 1666464484
transform 1 0 140672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1260
timestamp 1666464484
transform 1 0 142464 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1268
timestamp 1666464484
transform 1 0 143360 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1276
timestamp 1666464484
transform 1 0 144256 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1292
timestamp 1666464484
transform 1 0 146048 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1296
timestamp 1666464484
transform 1 0 146496 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1300
timestamp 1666464484
transform 1 0 146944 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1304
timestamp 1666464484
transform 1 0 147392 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1312
timestamp 1666464484
transform 1 0 148288 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1666464484
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1666464484
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1666464484
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1666464484
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1666464484
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1666464484
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1666464484
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1666464484
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1666464484
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1666464484
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1666464484
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1666464484
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1666464484
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1666464484
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1666464484
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1666464484
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1666464484
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1666464484
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_428
timestamp 1666464484
transform 1 0 49280 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1666464484
transform 1 0 56448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1666464484
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_499
timestamp 1666464484
transform 1 0 57232 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_563
timestamp 1666464484
transform 1 0 64400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1666464484
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_570
timestamp 1666464484
transform 1 0 65184 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_634
timestamp 1666464484
transform 1 0 72352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1666464484
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_641
timestamp 1666464484
transform 1 0 73136 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_705
timestamp 1666464484
transform 1 0 80304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_709
timestamp 1666464484
transform 1 0 80752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_712
timestamp 1666464484
transform 1 0 81088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_720
timestamp 1666464484
transform 1 0 81984 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_724
timestamp 1666464484
transform 1 0 82432 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_727
timestamp 1666464484
transform 1 0 82768 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_731
timestamp 1666464484
transform 1 0 83216 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_735
timestamp 1666464484
transform 1 0 83664 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_739
timestamp 1666464484
transform 1 0 84112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_741
timestamp 1666464484
transform 1 0 84336 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_744
timestamp 1666464484
transform 1 0 84672 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_776
timestamp 1666464484
transform 1 0 88256 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_779
timestamp 1666464484
transform 1 0 88592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_783
timestamp 1666464484
transform 1 0 89040 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_847
timestamp 1666464484
transform 1 0 96208 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_851
timestamp 1666464484
transform 1 0 96656 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_854
timestamp 1666464484
transform 1 0 96992 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_870
timestamp 1666464484
transform 1 0 98784 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_874
timestamp 1666464484
transform 1 0 99232 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_878
timestamp 1666464484
transform 1 0 99680 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_894
timestamp 1666464484
transform 1 0 101472 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_904
timestamp 1666464484
transform 1 0 102592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_908
timestamp 1666464484
transform 1 0 103040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_918
timestamp 1666464484
transform 1 0 104160 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_922
timestamp 1666464484
transform 1 0 104608 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_925
timestamp 1666464484
transform 1 0 104944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_932
timestamp 1666464484
transform 1 0 105728 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_964
timestamp 1666464484
transform 1 0 109312 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_968
timestamp 1666464484
transform 1 0 109760 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_970
timestamp 1666464484
transform 1 0 109984 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_973
timestamp 1666464484
transform 1 0 110320 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_983
timestamp 1666464484
transform 1 0 111440 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_991
timestamp 1666464484
transform 1 0 112336 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_993
timestamp 1666464484
transform 1 0 112560 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_996
timestamp 1666464484
transform 1 0 112896 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1000
timestamp 1666464484
transform 1 0 113344 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1004
timestamp 1666464484
transform 1 0 113792 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1008
timestamp 1666464484
transform 1 0 114240 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1016
timestamp 1666464484
transform 1 0 115136 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1018
timestamp 1666464484
transform 1 0 115360 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1021
timestamp 1666464484
transform 1 0 115696 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1025
timestamp 1666464484
transform 1 0 116144 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1029
timestamp 1666464484
transform 1 0 116592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1031
timestamp 1666464484
transform 1 0 116816 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1034
timestamp 1666464484
transform 1 0 117152 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1038
timestamp 1666464484
transform 1 0 117600 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1042
timestamp 1666464484
transform 1 0 118048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1046
timestamp 1666464484
transform 1 0 118496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1050
timestamp 1666464484
transform 1 0 118944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1053
timestamp 1666464484
transform 1 0 119280 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1061
timestamp 1666464484
transform 1 0 120176 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1067
timestamp 1666464484
transform 1 0 120848 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1083
timestamp 1666464484
transform 1 0 122640 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1091
timestamp 1666464484
transform 1 0 123536 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_1095
timestamp 1666464484
transform 1 0 123984 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1129
timestamp 1666464484
transform 1 0 127792 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1135
timestamp 1666464484
transform 1 0 128464 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1138
timestamp 1666464484
transform 1 0 128800 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1140
timestamp 1666464484
transform 1 0 129024 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1143
timestamp 1666464484
transform 1 0 129360 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1151
timestamp 1666464484
transform 1 0 130256 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1155
timestamp 1666464484
transform 1 0 130704 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1163
timestamp 1666464484
transform 1 0 131600 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1167
timestamp 1666464484
transform 1 0 132048 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1171
timestamp 1666464484
transform 1 0 132496 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1175
timestamp 1666464484
transform 1 0 132944 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1179
timestamp 1666464484
transform 1 0 133392 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1183
timestamp 1666464484
transform 1 0 133840 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1199
timestamp 1666464484
transform 1 0 135632 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1209
timestamp 1666464484
transform 1 0 136752 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1225
timestamp 1666464484
transform 1 0 138544 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1228
timestamp 1666464484
transform 1 0 138880 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1232
timestamp 1666464484
transform 1 0 139328 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1235
timestamp 1666464484
transform 1 0 139664 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1239
timestamp 1666464484
transform 1 0 140112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1247
timestamp 1666464484
transform 1 0 141008 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1255
timestamp 1666464484
transform 1 0 141904 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1263
timestamp 1666464484
transform 1 0 142800 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1267
timestamp 1666464484
transform 1 0 143248 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1271
timestamp 1666464484
transform 1 0 143696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1275
timestamp 1666464484
transform 1 0 144144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1277
timestamp 1666464484
transform 1 0 144368 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1280
timestamp 1666464484
transform 1 0 144704 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1296
timestamp 1666464484
transform 1 0 146496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1300
timestamp 1666464484
transform 1 0 146944 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1304
timestamp 1666464484
transform 1 0 147392 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1312
timestamp 1666464484
transform 1 0 148288 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1666464484
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1666464484
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1666464484
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1666464484
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1666464484
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1666464484
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1666464484
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1666464484
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1666464484
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1666464484
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1666464484
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1666464484
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1666464484
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1666464484
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1666464484
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1666464484
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1666464484
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1666464484
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1666464484
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1666464484
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_463
timestamp 1666464484
transform 1 0 53200 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1666464484
transform 1 0 60368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1666464484
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_534
timestamp 1666464484
transform 1 0 61152 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_598
timestamp 1666464484
transform 1 0 68320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1666464484
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_605
timestamp 1666464484
transform 1 0 69104 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_669
timestamp 1666464484
transform 1 0 76272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1666464484
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_676
timestamp 1666464484
transform 1 0 77056 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_740
timestamp 1666464484
transform 1 0 84224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_744
timestamp 1666464484
transform 1 0 84672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_747
timestamp 1666464484
transform 1 0 85008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_811
timestamp 1666464484
transform 1 0 92176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_815
timestamp 1666464484
transform 1 0 92624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_818
timestamp 1666464484
transform 1 0 92960 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_882
timestamp 1666464484
transform 1 0 100128 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_886
timestamp 1666464484
transform 1 0 100576 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_889
timestamp 1666464484
transform 1 0 100912 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_905
timestamp 1666464484
transform 1 0 102704 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_909
timestamp 1666464484
transform 1 0 103152 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_913
timestamp 1666464484
transform 1 0 103600 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_945
timestamp 1666464484
transform 1 0 107184 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_953
timestamp 1666464484
transform 1 0 108080 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_957
timestamp 1666464484
transform 1 0 108528 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_960
timestamp 1666464484
transform 1 0 108864 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_976
timestamp 1666464484
transform 1 0 110656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_980
timestamp 1666464484
transform 1 0 111104 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_982
timestamp 1666464484
transform 1 0 111328 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_985
timestamp 1666464484
transform 1 0 111664 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1017
timestamp 1666464484
transform 1 0 115248 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1025
timestamp 1666464484
transform 1 0 116144 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1031
timestamp 1666464484
transform 1 0 116816 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1095
timestamp 1666464484
transform 1 0 123984 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1099
timestamp 1666464484
transform 1 0 124432 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_1102
timestamp 1666464484
transform 1 0 124768 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1134
timestamp 1666464484
transform 1 0 128352 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1137
timestamp 1666464484
transform 1 0 128688 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1143
timestamp 1666464484
transform 1 0 129360 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1151
timestamp 1666464484
transform 1 0 130256 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1155
timestamp 1666464484
transform 1 0 130704 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1158
timestamp 1666464484
transform 1 0 131040 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1166
timestamp 1666464484
transform 1 0 131936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1170
timestamp 1666464484
transform 1 0 132384 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1173
timestamp 1666464484
transform 1 0 132720 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1237
timestamp 1666464484
transform 1 0 139888 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1241
timestamp 1666464484
transform 1 0 140336 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1244
timestamp 1666464484
transform 1 0 140672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1247
timestamp 1666464484
transform 1 0 141008 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_1251
timestamp 1666464484
transform 1 0 141456 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1283
timestamp 1666464484
transform 1 0 145040 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1299
timestamp 1666464484
transform 1 0 146832 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1301
timestamp 1666464484
transform 1 0 147056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1304
timestamp 1666464484
transform 1 0 147392 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1312
timestamp 1666464484
transform 1 0 148288 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1666464484
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1666464484
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1666464484
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1666464484
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1666464484
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1666464484
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1666464484
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1666464484
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1666464484
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1666464484
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1666464484
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1666464484
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1666464484
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1666464484
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1666464484
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1666464484
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1666464484
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1666464484
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1666464484
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1666464484
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1666464484
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_499
timestamp 1666464484
transform 1 0 57232 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_563
timestamp 1666464484
transform 1 0 64400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1666464484
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_570
timestamp 1666464484
transform 1 0 65184 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_634
timestamp 1666464484
transform 1 0 72352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1666464484
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_641
timestamp 1666464484
transform 1 0 73136 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_705
timestamp 1666464484
transform 1 0 80304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_709
timestamp 1666464484
transform 1 0 80752 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_712
timestamp 1666464484
transform 1 0 81088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_776
timestamp 1666464484
transform 1 0 88256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_780
timestamp 1666464484
transform 1 0 88704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_783
timestamp 1666464484
transform 1 0 89040 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_847
timestamp 1666464484
transform 1 0 96208 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_851
timestamp 1666464484
transform 1 0 96656 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_854
timestamp 1666464484
transform 1 0 96992 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_870
timestamp 1666464484
transform 1 0 98784 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_872
timestamp 1666464484
transform 1 0 99008 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_879
timestamp 1666464484
transform 1 0 99792 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_911
timestamp 1666464484
transform 1 0 103376 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_919
timestamp 1666464484
transform 1 0 104272 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_925
timestamp 1666464484
transform 1 0 104944 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_989
timestamp 1666464484
transform 1 0 112112 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_993
timestamp 1666464484
transform 1 0 112560 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_996
timestamp 1666464484
transform 1 0 112896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_1003
timestamp 1666464484
transform 1 0 113680 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_1035
timestamp 1666464484
transform 1 0 117264 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1051
timestamp 1666464484
transform 1 0 119056 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1059
timestamp 1666464484
transform 1 0 119952 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1063
timestamp 1666464484
transform 1 0 120400 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1067
timestamp 1666464484
transform 1 0 120848 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1131
timestamp 1666464484
transform 1 0 128016 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1135
timestamp 1666464484
transform 1 0 128464 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1138
timestamp 1666464484
transform 1 0 128800 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1202
timestamp 1666464484
transform 1 0 135968 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1206
timestamp 1666464484
transform 1 0 136416 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1209
timestamp 1666464484
transform 1 0 136752 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1273
timestamp 1666464484
transform 1 0 143920 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1277
timestamp 1666464484
transform 1 0 144368 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_1280
timestamp 1666464484
transform 1 0 144704 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1312
timestamp 1666464484
transform 1 0 148288 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1666464484
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1666464484
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1666464484
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1666464484
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1666464484
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1666464484
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1666464484
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1666464484
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1666464484
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1666464484
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1666464484
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1666464484
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1666464484
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1666464484
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1666464484
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1666464484
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1666464484
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1666464484
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1666464484
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1666464484
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1666464484
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1666464484
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_534
timestamp 1666464484
transform 1 0 61152 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_598
timestamp 1666464484
transform 1 0 68320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1666464484
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1666464484
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_669
timestamp 1666464484
transform 1 0 76272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1666464484
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_676
timestamp 1666464484
transform 1 0 77056 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_740
timestamp 1666464484
transform 1 0 84224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_744
timestamp 1666464484
transform 1 0 84672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_747
timestamp 1666464484
transform 1 0 85008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_811
timestamp 1666464484
transform 1 0 92176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_815
timestamp 1666464484
transform 1 0 92624 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_818
timestamp 1666464484
transform 1 0 92960 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_882
timestamp 1666464484
transform 1 0 100128 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_886
timestamp 1666464484
transform 1 0 100576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_889
timestamp 1666464484
transform 1 0 100912 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_953
timestamp 1666464484
transform 1 0 108080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_957
timestamp 1666464484
transform 1 0 108528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_960
timestamp 1666464484
transform 1 0 108864 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1024
timestamp 1666464484
transform 1 0 116032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1028
timestamp 1666464484
transform 1 0 116480 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1031
timestamp 1666464484
transform 1 0 116816 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1095
timestamp 1666464484
transform 1 0 123984 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1099
timestamp 1666464484
transform 1 0 124432 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1102
timestamp 1666464484
transform 1 0 124768 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1166
timestamp 1666464484
transform 1 0 131936 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1170
timestamp 1666464484
transform 1 0 132384 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1173
timestamp 1666464484
transform 1 0 132720 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1181
timestamp 1666464484
transform 1 0 133616 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1185
timestamp 1666464484
transform 1 0 134064 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1187
timestamp 1666464484
transform 1 0 134288 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1194
timestamp 1666464484
transform 1 0 135072 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_1198
timestamp 1666464484
transform 1 0 135520 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1230
timestamp 1666464484
transform 1 0 139104 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1238
timestamp 1666464484
transform 1 0 140000 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_1244
timestamp 1666464484
transform 1 0 140672 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_1276
timestamp 1666464484
transform 1 0 144256 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1292
timestamp 1666464484
transform 1 0 146048 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1300
timestamp 1666464484
transform 1 0 146944 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1304
timestamp 1666464484
transform 1 0 147392 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1312
timestamp 1666464484
transform 1 0 148288 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1666464484
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1666464484
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1666464484
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1666464484
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1666464484
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1666464484
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1666464484
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1666464484
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1666464484
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1666464484
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1666464484
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1666464484
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1666464484
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1666464484
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1666464484
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1666464484
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1666464484
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1666464484
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1666464484
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1666464484
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1666464484
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_499
timestamp 1666464484
transform 1 0 57232 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_563
timestamp 1666464484
transform 1 0 64400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1666464484
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_570
timestamp 1666464484
transform 1 0 65184 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_634
timestamp 1666464484
transform 1 0 72352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1666464484
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_641
timestamp 1666464484
transform 1 0 73136 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_705
timestamp 1666464484
transform 1 0 80304 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_709
timestamp 1666464484
transform 1 0 80752 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_712
timestamp 1666464484
transform 1 0 81088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_776
timestamp 1666464484
transform 1 0 88256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_780
timestamp 1666464484
transform 1 0 88704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_783
timestamp 1666464484
transform 1 0 89040 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_847
timestamp 1666464484
transform 1 0 96208 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_851
timestamp 1666464484
transform 1 0 96656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_854
timestamp 1666464484
transform 1 0 96992 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_918
timestamp 1666464484
transform 1 0 104160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_922
timestamp 1666464484
transform 1 0 104608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_925
timestamp 1666464484
transform 1 0 104944 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_989
timestamp 1666464484
transform 1 0 112112 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_993
timestamp 1666464484
transform 1 0 112560 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_996
timestamp 1666464484
transform 1 0 112896 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1060
timestamp 1666464484
transform 1 0 120064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1064
timestamp 1666464484
transform 1 0 120512 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1067
timestamp 1666464484
transform 1 0 120848 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1131
timestamp 1666464484
transform 1 0 128016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1135
timestamp 1666464484
transform 1 0 128464 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1138
timestamp 1666464484
transform 1 0 128800 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1202
timestamp 1666464484
transform 1 0 135968 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1206
timestamp 1666464484
transform 1 0 136416 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1209
timestamp 1666464484
transform 1 0 136752 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1273
timestamp 1666464484
transform 1 0 143920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1277
timestamp 1666464484
transform 1 0 144368 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_1280
timestamp 1666464484
transform 1 0 144704 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1296
timestamp 1666464484
transform 1 0 146496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1300
timestamp 1666464484
transform 1 0 146944 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1304
timestamp 1666464484
transform 1 0 147392 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1312
timestamp 1666464484
transform 1 0 148288 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1666464484
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1666464484
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1666464484
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1666464484
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1666464484
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1666464484
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1666464484
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1666464484
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1666464484
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1666464484
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1666464484
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1666464484
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1666464484
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1666464484
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1666464484
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1666464484
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1666464484
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1666464484
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1666464484
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1666464484
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1666464484
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1666464484
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1666464484
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1666464484
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_598
timestamp 1666464484
transform 1 0 68320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1666464484
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1666464484
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_669
timestamp 1666464484
transform 1 0 76272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1666464484
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_676
timestamp 1666464484
transform 1 0 77056 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_740
timestamp 1666464484
transform 1 0 84224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_744
timestamp 1666464484
transform 1 0 84672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_747
timestamp 1666464484
transform 1 0 85008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_811
timestamp 1666464484
transform 1 0 92176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_815
timestamp 1666464484
transform 1 0 92624 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_818
timestamp 1666464484
transform 1 0 92960 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_882
timestamp 1666464484
transform 1 0 100128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_886
timestamp 1666464484
transform 1 0 100576 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_889
timestamp 1666464484
transform 1 0 100912 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_953
timestamp 1666464484
transform 1 0 108080 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_957
timestamp 1666464484
transform 1 0 108528 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_960
timestamp 1666464484
transform 1 0 108864 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1024
timestamp 1666464484
transform 1 0 116032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1028
timestamp 1666464484
transform 1 0 116480 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1031
timestamp 1666464484
transform 1 0 116816 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1095
timestamp 1666464484
transform 1 0 123984 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1099
timestamp 1666464484
transform 1 0 124432 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1102
timestamp 1666464484
transform 1 0 124768 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1166
timestamp 1666464484
transform 1 0 131936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1170
timestamp 1666464484
transform 1 0 132384 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1173
timestamp 1666464484
transform 1 0 132720 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1237
timestamp 1666464484
transform 1 0 139888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1241
timestamp 1666464484
transform 1 0 140336 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_1244
timestamp 1666464484
transform 1 0 140672 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_1276
timestamp 1666464484
transform 1 0 144256 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_1292
timestamp 1666464484
transform 1 0 146048 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1300
timestamp 1666464484
transform 1 0 146944 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1304
timestamp 1666464484
transform 1 0 147392 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1312
timestamp 1666464484
transform 1 0 148288 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1666464484
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1666464484
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1666464484
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1666464484
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1666464484
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1666464484
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1666464484
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1666464484
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1666464484
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1666464484
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1666464484
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1666464484
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1666464484
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1666464484
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1666464484
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1666464484
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1666464484
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1666464484
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1666464484
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1666464484
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1666464484
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1666464484
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_563
timestamp 1666464484
transform 1 0 64400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1666464484
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1666464484
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1666464484
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1666464484
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_641
timestamp 1666464484
transform 1 0 73136 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_705
timestamp 1666464484
transform 1 0 80304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_709
timestamp 1666464484
transform 1 0 80752 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_712
timestamp 1666464484
transform 1 0 81088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_776
timestamp 1666464484
transform 1 0 88256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_780
timestamp 1666464484
transform 1 0 88704 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_783
timestamp 1666464484
transform 1 0 89040 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_847
timestamp 1666464484
transform 1 0 96208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_851
timestamp 1666464484
transform 1 0 96656 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_854
timestamp 1666464484
transform 1 0 96992 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_918
timestamp 1666464484
transform 1 0 104160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_922
timestamp 1666464484
transform 1 0 104608 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_925
timestamp 1666464484
transform 1 0 104944 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_989
timestamp 1666464484
transform 1 0 112112 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_993
timestamp 1666464484
transform 1 0 112560 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_996
timestamp 1666464484
transform 1 0 112896 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1060
timestamp 1666464484
transform 1 0 120064 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1064
timestamp 1666464484
transform 1 0 120512 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1067
timestamp 1666464484
transform 1 0 120848 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1131
timestamp 1666464484
transform 1 0 128016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1135
timestamp 1666464484
transform 1 0 128464 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1138
timestamp 1666464484
transform 1 0 128800 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1202
timestamp 1666464484
transform 1 0 135968 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1206
timestamp 1666464484
transform 1 0 136416 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1209
timestamp 1666464484
transform 1 0 136752 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1273
timestamp 1666464484
transform 1 0 143920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1277
timestamp 1666464484
transform 1 0 144368 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_1280
timestamp 1666464484
transform 1 0 144704 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1296
timestamp 1666464484
transform 1 0 146496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1300
timestamp 1666464484
transform 1 0 146944 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1304
timestamp 1666464484
transform 1 0 147392 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1312
timestamp 1666464484
transform 1 0 148288 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1666464484
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1666464484
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1666464484
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1666464484
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1666464484
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1666464484
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1666464484
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1666464484
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1666464484
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1666464484
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1666464484
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1666464484
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1666464484
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1666464484
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1666464484
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1666464484
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1666464484
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1666464484
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1666464484
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1666464484
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1666464484
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1666464484
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1666464484
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1666464484
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_598
timestamp 1666464484
transform 1 0 68320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1666464484
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_605
timestamp 1666464484
transform 1 0 69104 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_669
timestamp 1666464484
transform 1 0 76272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1666464484
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_676
timestamp 1666464484
transform 1 0 77056 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_740
timestamp 1666464484
transform 1 0 84224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_744
timestamp 1666464484
transform 1 0 84672 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_747
timestamp 1666464484
transform 1 0 85008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_811
timestamp 1666464484
transform 1 0 92176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_815
timestamp 1666464484
transform 1 0 92624 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_818
timestamp 1666464484
transform 1 0 92960 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_850
timestamp 1666464484
transform 1 0 96544 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_866
timestamp 1666464484
transform 1 0 98336 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_874
timestamp 1666464484
transform 1 0 99232 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_881
timestamp 1666464484
transform 1 0 100016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_885
timestamp 1666464484
transform 1 0 100464 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_889
timestamp 1666464484
transform 1 0 100912 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_953
timestamp 1666464484
transform 1 0 108080 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_957
timestamp 1666464484
transform 1 0 108528 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_960
timestamp 1666464484
transform 1 0 108864 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1024
timestamp 1666464484
transform 1 0 116032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1028
timestamp 1666464484
transform 1 0 116480 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1031
timestamp 1666464484
transform 1 0 116816 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1095
timestamp 1666464484
transform 1 0 123984 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1099
timestamp 1666464484
transform 1 0 124432 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1102
timestamp 1666464484
transform 1 0 124768 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1166
timestamp 1666464484
transform 1 0 131936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1170
timestamp 1666464484
transform 1 0 132384 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1173
timestamp 1666464484
transform 1 0 132720 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1237
timestamp 1666464484
transform 1 0 139888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1241
timestamp 1666464484
transform 1 0 140336 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_1244
timestamp 1666464484
transform 1 0 140672 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_1276
timestamp 1666464484
transform 1 0 144256 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_1292
timestamp 1666464484
transform 1 0 146048 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_1296
timestamp 1666464484
transform 1 0 146496 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1312
timestamp 1666464484
transform 1 0 148288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1666464484
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1666464484
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1666464484
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1666464484
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1666464484
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1666464484
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1666464484
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1666464484
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1666464484
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1666464484
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1666464484
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1666464484
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1666464484
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1666464484
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1666464484
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1666464484
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1666464484
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1666464484
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1666464484
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1666464484
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1666464484
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1666464484
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_563
timestamp 1666464484
transform 1 0 64400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1666464484
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1666464484
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1666464484
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1666464484
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_641
timestamp 1666464484
transform 1 0 73136 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_705
timestamp 1666464484
transform 1 0 80304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_709
timestamp 1666464484
transform 1 0 80752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_712
timestamp 1666464484
transform 1 0 81088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_776
timestamp 1666464484
transform 1 0 88256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_780
timestamp 1666464484
transform 1 0 88704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_783
timestamp 1666464484
transform 1 0 89040 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_847
timestamp 1666464484
transform 1 0 96208 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_851
timestamp 1666464484
transform 1 0 96656 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_854
timestamp 1666464484
transform 1 0 96992 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_870
timestamp 1666464484
transform 1 0 98784 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_878
timestamp 1666464484
transform 1 0 99680 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_882
timestamp 1666464484
transform 1 0 100128 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_889
timestamp 1666464484
transform 1 0 100912 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_893
timestamp 1666464484
transform 1 0 101360 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_909
timestamp 1666464484
transform 1 0 103152 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_917
timestamp 1666464484
transform 1 0 104048 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_921
timestamp 1666464484
transform 1 0 104496 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_925
timestamp 1666464484
transform 1 0 104944 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_989
timestamp 1666464484
transform 1 0 112112 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_993
timestamp 1666464484
transform 1 0 112560 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_996
timestamp 1666464484
transform 1 0 112896 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1060
timestamp 1666464484
transform 1 0 120064 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1064
timestamp 1666464484
transform 1 0 120512 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1067
timestamp 1666464484
transform 1 0 120848 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1131
timestamp 1666464484
transform 1 0 128016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1135
timestamp 1666464484
transform 1 0 128464 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1138
timestamp 1666464484
transform 1 0 128800 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1202
timestamp 1666464484
transform 1 0 135968 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1206
timestamp 1666464484
transform 1 0 136416 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1209
timestamp 1666464484
transform 1 0 136752 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1273
timestamp 1666464484
transform 1 0 143920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1277
timestamp 1666464484
transform 1 0 144368 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_1280
timestamp 1666464484
transform 1 0 144704 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1288
timestamp 1666464484
transform 1 0 145600 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_1292
timestamp 1666464484
transform 1 0 146048 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_1296
timestamp 1666464484
transform 1 0 146496 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1312
timestamp 1666464484
transform 1 0 148288 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1666464484
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1666464484
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1666464484
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1666464484
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1666464484
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1666464484
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1666464484
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1666464484
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1666464484
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1666464484
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1666464484
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1666464484
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1666464484
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1666464484
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1666464484
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1666464484
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1666464484
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1666464484
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1666464484
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1666464484
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1666464484
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1666464484
transform 1 0 60368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1666464484
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1666464484
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_598
timestamp 1666464484
transform 1 0 68320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1666464484
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1666464484
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_669
timestamp 1666464484
transform 1 0 76272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1666464484
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_676
timestamp 1666464484
transform 1 0 77056 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_740
timestamp 1666464484
transform 1 0 84224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_744
timestamp 1666464484
transform 1 0 84672 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_747
timestamp 1666464484
transform 1 0 85008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_811
timestamp 1666464484
transform 1 0 92176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_815
timestamp 1666464484
transform 1 0 92624 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_818
timestamp 1666464484
transform 1 0 92960 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_882
timestamp 1666464484
transform 1 0 100128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_886
timestamp 1666464484
transform 1 0 100576 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_889
timestamp 1666464484
transform 1 0 100912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_899
timestamp 1666464484
transform 1 0 102032 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_931
timestamp 1666464484
transform 1 0 105616 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_947
timestamp 1666464484
transform 1 0 107408 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_955
timestamp 1666464484
transform 1 0 108304 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_957
timestamp 1666464484
transform 1 0 108528 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_960
timestamp 1666464484
transform 1 0 108864 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1024
timestamp 1666464484
transform 1 0 116032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1028
timestamp 1666464484
transform 1 0 116480 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1031
timestamp 1666464484
transform 1 0 116816 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1095
timestamp 1666464484
transform 1 0 123984 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1099
timestamp 1666464484
transform 1 0 124432 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1102
timestamp 1666464484
transform 1 0 124768 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1166
timestamp 1666464484
transform 1 0 131936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1170
timestamp 1666464484
transform 1 0 132384 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1173
timestamp 1666464484
transform 1 0 132720 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1237
timestamp 1666464484
transform 1 0 139888 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1241
timestamp 1666464484
transform 1 0 140336 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_1244
timestamp 1666464484
transform 1 0 140672 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_1276
timestamp 1666464484
transform 1 0 144256 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_1292
timestamp 1666464484
transform 1 0 146048 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_1296
timestamp 1666464484
transform 1 0 146496 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1312
timestamp 1666464484
transform 1 0 148288 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1666464484
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1666464484
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1666464484
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1666464484
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1666464484
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1666464484
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1666464484
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1666464484
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1666464484
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1666464484
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1666464484
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1666464484
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1666464484
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1666464484
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1666464484
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1666464484
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1666464484
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1666464484
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1666464484
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1666464484
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1666464484
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_499
timestamp 1666464484
transform 1 0 57232 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_563
timestamp 1666464484
transform 1 0 64400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1666464484
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1666464484
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1666464484
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1666464484
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_641
timestamp 1666464484
transform 1 0 73136 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_705
timestamp 1666464484
transform 1 0 80304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_709
timestamp 1666464484
transform 1 0 80752 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_712
timestamp 1666464484
transform 1 0 81088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_776
timestamp 1666464484
transform 1 0 88256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_780
timestamp 1666464484
transform 1 0 88704 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_783
timestamp 1666464484
transform 1 0 89040 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_847
timestamp 1666464484
transform 1 0 96208 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_851
timestamp 1666464484
transform 1 0 96656 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_854
timestamp 1666464484
transform 1 0 96992 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_918
timestamp 1666464484
transform 1 0 104160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_922
timestamp 1666464484
transform 1 0 104608 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_925
timestamp 1666464484
transform 1 0 104944 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_989
timestamp 1666464484
transform 1 0 112112 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_993
timestamp 1666464484
transform 1 0 112560 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_996
timestamp 1666464484
transform 1 0 112896 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1060
timestamp 1666464484
transform 1 0 120064 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1064
timestamp 1666464484
transform 1 0 120512 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1067
timestamp 1666464484
transform 1 0 120848 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1131
timestamp 1666464484
transform 1 0 128016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1135
timestamp 1666464484
transform 1 0 128464 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1138
timestamp 1666464484
transform 1 0 128800 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1202
timestamp 1666464484
transform 1 0 135968 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1206
timestamp 1666464484
transform 1 0 136416 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1209
timestamp 1666464484
transform 1 0 136752 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1273
timestamp 1666464484
transform 1 0 143920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1277
timestamp 1666464484
transform 1 0 144368 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_1280
timestamp 1666464484
transform 1 0 144704 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1312
timestamp 1666464484
transform 1 0 148288 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1666464484
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1666464484
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1666464484
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1666464484
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1666464484
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1666464484
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1666464484
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1666464484
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1666464484
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1666464484
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1666464484
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1666464484
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1666464484
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1666464484
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1666464484
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1666464484
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1666464484
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1666464484
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1666464484
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1666464484
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_463
timestamp 1666464484
transform 1 0 53200 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1666464484
transform 1 0 60368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1666464484
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1666464484
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1666464484
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1666464484
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1666464484
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_669
timestamp 1666464484
transform 1 0 76272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1666464484
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_676
timestamp 1666464484
transform 1 0 77056 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_740
timestamp 1666464484
transform 1 0 84224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_744
timestamp 1666464484
transform 1 0 84672 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_747
timestamp 1666464484
transform 1 0 85008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_811
timestamp 1666464484
transform 1 0 92176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_815
timestamp 1666464484
transform 1 0 92624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_818
timestamp 1666464484
transform 1 0 92960 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_882
timestamp 1666464484
transform 1 0 100128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_886
timestamp 1666464484
transform 1 0 100576 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_889
timestamp 1666464484
transform 1 0 100912 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_953
timestamp 1666464484
transform 1 0 108080 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_957
timestamp 1666464484
transform 1 0 108528 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_960
timestamp 1666464484
transform 1 0 108864 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1024
timestamp 1666464484
transform 1 0 116032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1028
timestamp 1666464484
transform 1 0 116480 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1031
timestamp 1666464484
transform 1 0 116816 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1095
timestamp 1666464484
transform 1 0 123984 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1099
timestamp 1666464484
transform 1 0 124432 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1102
timestamp 1666464484
transform 1 0 124768 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1166
timestamp 1666464484
transform 1 0 131936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1170
timestamp 1666464484
transform 1 0 132384 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1173
timestamp 1666464484
transform 1 0 132720 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1237
timestamp 1666464484
transform 1 0 139888 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1241
timestamp 1666464484
transform 1 0 140336 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_1244
timestamp 1666464484
transform 1 0 140672 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_1276
timestamp 1666464484
transform 1 0 144256 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_1292
timestamp 1666464484
transform 1 0 146048 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_1296
timestamp 1666464484
transform 1 0 146496 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1312
timestamp 1666464484
transform 1 0 148288 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1666464484
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1666464484
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1666464484
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1666464484
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1666464484
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1666464484
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1666464484
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1666464484
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1666464484
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1666464484
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1666464484
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1666464484
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1666464484
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1666464484
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1666464484
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1666464484
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1666464484
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1666464484
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1666464484
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1666464484
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1666464484
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1666464484
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1666464484
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1666464484
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1666464484
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1666464484
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1666464484
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_641
timestamp 1666464484
transform 1 0 73136 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_705
timestamp 1666464484
transform 1 0 80304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_709
timestamp 1666464484
transform 1 0 80752 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_712
timestamp 1666464484
transform 1 0 81088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_776
timestamp 1666464484
transform 1 0 88256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_780
timestamp 1666464484
transform 1 0 88704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_783
timestamp 1666464484
transform 1 0 89040 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_847
timestamp 1666464484
transform 1 0 96208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_851
timestamp 1666464484
transform 1 0 96656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_854
timestamp 1666464484
transform 1 0 96992 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_918
timestamp 1666464484
transform 1 0 104160 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_922
timestamp 1666464484
transform 1 0 104608 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_925
timestamp 1666464484
transform 1 0 104944 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_989
timestamp 1666464484
transform 1 0 112112 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_993
timestamp 1666464484
transform 1 0 112560 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_996
timestamp 1666464484
transform 1 0 112896 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1060
timestamp 1666464484
transform 1 0 120064 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1064
timestamp 1666464484
transform 1 0 120512 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1067
timestamp 1666464484
transform 1 0 120848 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1131
timestamp 1666464484
transform 1 0 128016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1135
timestamp 1666464484
transform 1 0 128464 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1138
timestamp 1666464484
transform 1 0 128800 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1202
timestamp 1666464484
transform 1 0 135968 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1206
timestamp 1666464484
transform 1 0 136416 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1209
timestamp 1666464484
transform 1 0 136752 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1273
timestamp 1666464484
transform 1 0 143920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1277
timestamp 1666464484
transform 1 0 144368 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_1280
timestamp 1666464484
transform 1 0 144704 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1288
timestamp 1666464484
transform 1 0 145600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_1292
timestamp 1666464484
transform 1 0 146048 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_1296
timestamp 1666464484
transform 1 0 146496 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1312
timestamp 1666464484
transform 1 0 148288 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1666464484
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1666464484
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1666464484
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1666464484
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1666464484
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1666464484
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1666464484
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1666464484
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1666464484
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1666464484
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1666464484
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1666464484
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1666464484
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1666464484
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1666464484
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1666464484
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1666464484
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1666464484
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1666464484
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1666464484
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1666464484
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1666464484
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1666464484
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1666464484
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_598
timestamp 1666464484
transform 1 0 68320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1666464484
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_605
timestamp 1666464484
transform 1 0 69104 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_669
timestamp 1666464484
transform 1 0 76272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_673
timestamp 1666464484
transform 1 0 76720 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_676
timestamp 1666464484
transform 1 0 77056 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_740
timestamp 1666464484
transform 1 0 84224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_744
timestamp 1666464484
transform 1 0 84672 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_747
timestamp 1666464484
transform 1 0 85008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_811
timestamp 1666464484
transform 1 0 92176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_815
timestamp 1666464484
transform 1 0 92624 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_818
timestamp 1666464484
transform 1 0 92960 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_882
timestamp 1666464484
transform 1 0 100128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_886
timestamp 1666464484
transform 1 0 100576 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_889
timestamp 1666464484
transform 1 0 100912 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_953
timestamp 1666464484
transform 1 0 108080 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_957
timestamp 1666464484
transform 1 0 108528 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_960
timestamp 1666464484
transform 1 0 108864 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1024
timestamp 1666464484
transform 1 0 116032 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1028
timestamp 1666464484
transform 1 0 116480 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1031
timestamp 1666464484
transform 1 0 116816 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1095
timestamp 1666464484
transform 1 0 123984 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1099
timestamp 1666464484
transform 1 0 124432 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1102
timestamp 1666464484
transform 1 0 124768 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1166
timestamp 1666464484
transform 1 0 131936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1170
timestamp 1666464484
transform 1 0 132384 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1173
timestamp 1666464484
transform 1 0 132720 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1237
timestamp 1666464484
transform 1 0 139888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1241
timestamp 1666464484
transform 1 0 140336 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_1244
timestamp 1666464484
transform 1 0 140672 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1276
timestamp 1666464484
transform 1 0 144256 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1292
timestamp 1666464484
transform 1 0 146048 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1296
timestamp 1666464484
transform 1 0 146496 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1312
timestamp 1666464484
transform 1 0 148288 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1666464484
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1666464484
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1666464484
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1666464484
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1666464484
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1666464484
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1666464484
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1666464484
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1666464484
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1666464484
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1666464484
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1666464484
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1666464484
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1666464484
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1666464484
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1666464484
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1666464484
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1666464484
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1666464484
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1666464484
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1666464484
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1666464484
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_563
timestamp 1666464484
transform 1 0 64400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1666464484
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1666464484
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_634
timestamp 1666464484
transform 1 0 72352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1666464484
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_641
timestamp 1666464484
transform 1 0 73136 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_705
timestamp 1666464484
transform 1 0 80304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_709
timestamp 1666464484
transform 1 0 80752 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_712
timestamp 1666464484
transform 1 0 81088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_776
timestamp 1666464484
transform 1 0 88256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_780
timestamp 1666464484
transform 1 0 88704 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_783
timestamp 1666464484
transform 1 0 89040 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_847
timestamp 1666464484
transform 1 0 96208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_851
timestamp 1666464484
transform 1 0 96656 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_854
timestamp 1666464484
transform 1 0 96992 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_918
timestamp 1666464484
transform 1 0 104160 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_922
timestamp 1666464484
transform 1 0 104608 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_925
timestamp 1666464484
transform 1 0 104944 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_989
timestamp 1666464484
transform 1 0 112112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_993
timestamp 1666464484
transform 1 0 112560 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_996
timestamp 1666464484
transform 1 0 112896 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1060
timestamp 1666464484
transform 1 0 120064 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1064
timestamp 1666464484
transform 1 0 120512 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1067
timestamp 1666464484
transform 1 0 120848 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1131
timestamp 1666464484
transform 1 0 128016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1135
timestamp 1666464484
transform 1 0 128464 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1138
timestamp 1666464484
transform 1 0 128800 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1202
timestamp 1666464484
transform 1 0 135968 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1206
timestamp 1666464484
transform 1 0 136416 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1209
timestamp 1666464484
transform 1 0 136752 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1273
timestamp 1666464484
transform 1 0 143920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1277
timestamp 1666464484
transform 1 0 144368 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_1280
timestamp 1666464484
transform 1 0 144704 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1288
timestamp 1666464484
transform 1 0 145600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_1292
timestamp 1666464484
transform 1 0 146048 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_1296
timestamp 1666464484
transform 1 0 146496 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1312
timestamp 1666464484
transform 1 0 148288 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1666464484
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1666464484
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1666464484
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1666464484
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1666464484
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1666464484
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1666464484
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1666464484
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1666464484
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1666464484
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1666464484
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1666464484
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1666464484
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1666464484
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1666464484
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1666464484
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1666464484
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1666464484
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1666464484
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1666464484
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_463
timestamp 1666464484
transform 1 0 53200 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_527
timestamp 1666464484
transform 1 0 60368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1666464484
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1666464484
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_598
timestamp 1666464484
transform 1 0 68320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1666464484
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_605
timestamp 1666464484
transform 1 0 69104 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_669
timestamp 1666464484
transform 1 0 76272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_673
timestamp 1666464484
transform 1 0 76720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_676
timestamp 1666464484
transform 1 0 77056 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_740
timestamp 1666464484
transform 1 0 84224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_744
timestamp 1666464484
transform 1 0 84672 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_747
timestamp 1666464484
transform 1 0 85008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_811
timestamp 1666464484
transform 1 0 92176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_815
timestamp 1666464484
transform 1 0 92624 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_818
timestamp 1666464484
transform 1 0 92960 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_882
timestamp 1666464484
transform 1 0 100128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_886
timestamp 1666464484
transform 1 0 100576 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_889
timestamp 1666464484
transform 1 0 100912 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_953
timestamp 1666464484
transform 1 0 108080 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_957
timestamp 1666464484
transform 1 0 108528 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_960
timestamp 1666464484
transform 1 0 108864 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1024
timestamp 1666464484
transform 1 0 116032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1028
timestamp 1666464484
transform 1 0 116480 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1031
timestamp 1666464484
transform 1 0 116816 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1095
timestamp 1666464484
transform 1 0 123984 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1099
timestamp 1666464484
transform 1 0 124432 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1102
timestamp 1666464484
transform 1 0 124768 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1166
timestamp 1666464484
transform 1 0 131936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1170
timestamp 1666464484
transform 1 0 132384 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1173
timestamp 1666464484
transform 1 0 132720 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1237
timestamp 1666464484
transform 1 0 139888 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1241
timestamp 1666464484
transform 1 0 140336 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_1244
timestamp 1666464484
transform 1 0 140672 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_1276
timestamp 1666464484
transform 1 0 144256 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_1292
timestamp 1666464484
transform 1 0 146048 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_1296
timestamp 1666464484
transform 1 0 146496 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1312
timestamp 1666464484
transform 1 0 148288 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1666464484
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1666464484
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1666464484
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1666464484
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1666464484
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1666464484
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1666464484
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1666464484
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1666464484
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1666464484
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1666464484
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1666464484
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1666464484
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1666464484
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1666464484
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1666464484
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1666464484
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1666464484
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1666464484
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1666464484
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1666464484
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1666464484
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_563
timestamp 1666464484
transform 1 0 64400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1666464484
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1666464484
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1666464484
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1666464484
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_641
timestamp 1666464484
transform 1 0 73136 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_705
timestamp 1666464484
transform 1 0 80304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_709
timestamp 1666464484
transform 1 0 80752 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_712
timestamp 1666464484
transform 1 0 81088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_776
timestamp 1666464484
transform 1 0 88256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_780
timestamp 1666464484
transform 1 0 88704 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_783
timestamp 1666464484
transform 1 0 89040 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_847
timestamp 1666464484
transform 1 0 96208 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_851
timestamp 1666464484
transform 1 0 96656 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_854
timestamp 1666464484
transform 1 0 96992 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_918
timestamp 1666464484
transform 1 0 104160 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_922
timestamp 1666464484
transform 1 0 104608 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_925
timestamp 1666464484
transform 1 0 104944 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_989
timestamp 1666464484
transform 1 0 112112 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_993
timestamp 1666464484
transform 1 0 112560 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_996
timestamp 1666464484
transform 1 0 112896 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_1000
timestamp 1666464484
transform 1 0 113344 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_1008
timestamp 1666464484
transform 1 0 114240 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_1040
timestamp 1666464484
transform 1 0 117824 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_1056
timestamp 1666464484
transform 1 0 119616 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1064
timestamp 1666464484
transform 1 0 120512 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1067
timestamp 1666464484
transform 1 0 120848 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1131
timestamp 1666464484
transform 1 0 128016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1135
timestamp 1666464484
transform 1 0 128464 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1138
timestamp 1666464484
transform 1 0 128800 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1202
timestamp 1666464484
transform 1 0 135968 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1206
timestamp 1666464484
transform 1 0 136416 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1209
timestamp 1666464484
transform 1 0 136752 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1273
timestamp 1666464484
transform 1 0 143920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1277
timestamp 1666464484
transform 1 0 144368 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_1280
timestamp 1666464484
transform 1 0 144704 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1288
timestamp 1666464484
transform 1 0 145600 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_1292
timestamp 1666464484
transform 1 0 146048 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_1296
timestamp 1666464484
transform 1 0 146496 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1312
timestamp 1666464484
transform 1 0 148288 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1666464484
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1666464484
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1666464484
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1666464484
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1666464484
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1666464484
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1666464484
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1666464484
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1666464484
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1666464484
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1666464484
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1666464484
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1666464484
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1666464484
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1666464484
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1666464484
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1666464484
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1666464484
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1666464484
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1666464484
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1666464484
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_527
timestamp 1666464484
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1666464484
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1666464484
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_598
timestamp 1666464484
transform 1 0 68320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1666464484
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_605
timestamp 1666464484
transform 1 0 69104 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_669
timestamp 1666464484
transform 1 0 76272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_673
timestamp 1666464484
transform 1 0 76720 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_676
timestamp 1666464484
transform 1 0 77056 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_740
timestamp 1666464484
transform 1 0 84224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_744
timestamp 1666464484
transform 1 0 84672 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_747
timestamp 1666464484
transform 1 0 85008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_811
timestamp 1666464484
transform 1 0 92176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_815
timestamp 1666464484
transform 1 0 92624 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_818
timestamp 1666464484
transform 1 0 92960 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_882
timestamp 1666464484
transform 1 0 100128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_886
timestamp 1666464484
transform 1 0 100576 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_889
timestamp 1666464484
transform 1 0 100912 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_953
timestamp 1666464484
transform 1 0 108080 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_957
timestamp 1666464484
transform 1 0 108528 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_960
timestamp 1666464484
transform 1 0 108864 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1024
timestamp 1666464484
transform 1 0 116032 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1028
timestamp 1666464484
transform 1 0 116480 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1031
timestamp 1666464484
transform 1 0 116816 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1095
timestamp 1666464484
transform 1 0 123984 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1099
timestamp 1666464484
transform 1 0 124432 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1102
timestamp 1666464484
transform 1 0 124768 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1166
timestamp 1666464484
transform 1 0 131936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1170
timestamp 1666464484
transform 1 0 132384 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1173
timestamp 1666464484
transform 1 0 132720 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1237
timestamp 1666464484
transform 1 0 139888 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1241
timestamp 1666464484
transform 1 0 140336 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_1244
timestamp 1666464484
transform 1 0 140672 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_1276
timestamp 1666464484
transform 1 0 144256 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_1292
timestamp 1666464484
transform 1 0 146048 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_1296
timestamp 1666464484
transform 1 0 146496 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1312
timestamp 1666464484
transform 1 0 148288 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1666464484
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1666464484
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1666464484
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1666464484
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1666464484
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1666464484
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1666464484
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1666464484
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1666464484
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1666464484
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1666464484
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1666464484
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1666464484
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1666464484
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1666464484
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1666464484
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1666464484
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1666464484
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1666464484
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1666464484
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1666464484
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1666464484
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_563
timestamp 1666464484
transform 1 0 64400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1666464484
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1666464484
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_634
timestamp 1666464484
transform 1 0 72352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1666464484
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_641
timestamp 1666464484
transform 1 0 73136 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_705
timestamp 1666464484
transform 1 0 80304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_709
timestamp 1666464484
transform 1 0 80752 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_712
timestamp 1666464484
transform 1 0 81088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_776
timestamp 1666464484
transform 1 0 88256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_780
timestamp 1666464484
transform 1 0 88704 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_783
timestamp 1666464484
transform 1 0 89040 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_847
timestamp 1666464484
transform 1 0 96208 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_851
timestamp 1666464484
transform 1 0 96656 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_854
timestamp 1666464484
transform 1 0 96992 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_918
timestamp 1666464484
transform 1 0 104160 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_922
timestamp 1666464484
transform 1 0 104608 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_925
timestamp 1666464484
transform 1 0 104944 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_989
timestamp 1666464484
transform 1 0 112112 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_993
timestamp 1666464484
transform 1 0 112560 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_996
timestamp 1666464484
transform 1 0 112896 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1060
timestamp 1666464484
transform 1 0 120064 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1064
timestamp 1666464484
transform 1 0 120512 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1067
timestamp 1666464484
transform 1 0 120848 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1131
timestamp 1666464484
transform 1 0 128016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1135
timestamp 1666464484
transform 1 0 128464 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1138
timestamp 1666464484
transform 1 0 128800 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1202
timestamp 1666464484
transform 1 0 135968 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1206
timestamp 1666464484
transform 1 0 136416 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1209
timestamp 1666464484
transform 1 0 136752 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1273
timestamp 1666464484
transform 1 0 143920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1277
timestamp 1666464484
transform 1 0 144368 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_1280
timestamp 1666464484
transform 1 0 144704 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1312
timestamp 1666464484
transform 1 0 148288 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1666464484
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1666464484
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1666464484
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1666464484
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1666464484
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1666464484
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1666464484
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1666464484
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1666464484
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1666464484
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1666464484
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1666464484
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1666464484
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1666464484
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1666464484
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1666464484
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1666464484
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1666464484
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1666464484
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1666464484
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1666464484
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_527
timestamp 1666464484
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1666464484
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1666464484
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_598
timestamp 1666464484
transform 1 0 68320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1666464484
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_605
timestamp 1666464484
transform 1 0 69104 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_669
timestamp 1666464484
transform 1 0 76272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_673
timestamp 1666464484
transform 1 0 76720 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_676
timestamp 1666464484
transform 1 0 77056 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_740
timestamp 1666464484
transform 1 0 84224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_744
timestamp 1666464484
transform 1 0 84672 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_747
timestamp 1666464484
transform 1 0 85008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_811
timestamp 1666464484
transform 1 0 92176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_815
timestamp 1666464484
transform 1 0 92624 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_818
timestamp 1666464484
transform 1 0 92960 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_882
timestamp 1666464484
transform 1 0 100128 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_886
timestamp 1666464484
transform 1 0 100576 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_889
timestamp 1666464484
transform 1 0 100912 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_953
timestamp 1666464484
transform 1 0 108080 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_957
timestamp 1666464484
transform 1 0 108528 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_960
timestamp 1666464484
transform 1 0 108864 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1024
timestamp 1666464484
transform 1 0 116032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1028
timestamp 1666464484
transform 1 0 116480 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1031
timestamp 1666464484
transform 1 0 116816 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1095
timestamp 1666464484
transform 1 0 123984 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1099
timestamp 1666464484
transform 1 0 124432 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1102
timestamp 1666464484
transform 1 0 124768 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1166
timestamp 1666464484
transform 1 0 131936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1170
timestamp 1666464484
transform 1 0 132384 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1173
timestamp 1666464484
transform 1 0 132720 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1237
timestamp 1666464484
transform 1 0 139888 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1241
timestamp 1666464484
transform 1 0 140336 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_1244
timestamp 1666464484
transform 1 0 140672 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_1276
timestamp 1666464484
transform 1 0 144256 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_1292
timestamp 1666464484
transform 1 0 146048 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_1296
timestamp 1666464484
transform 1 0 146496 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1312
timestamp 1666464484
transform 1 0 148288 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1666464484
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1666464484
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1666464484
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1666464484
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1666464484
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1666464484
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1666464484
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1666464484
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1666464484
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1666464484
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1666464484
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1666464484
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1666464484
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1666464484
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1666464484
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1666464484
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1666464484
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1666464484
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1666464484
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1666464484
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1666464484
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1666464484
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_563
timestamp 1666464484
transform 1 0 64400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1666464484
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1666464484
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_634
timestamp 1666464484
transform 1 0 72352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1666464484
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_641
timestamp 1666464484
transform 1 0 73136 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_705
timestamp 1666464484
transform 1 0 80304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_709
timestamp 1666464484
transform 1 0 80752 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_712
timestamp 1666464484
transform 1 0 81088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_776
timestamp 1666464484
transform 1 0 88256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_780
timestamp 1666464484
transform 1 0 88704 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_783
timestamp 1666464484
transform 1 0 89040 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_847
timestamp 1666464484
transform 1 0 96208 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_851
timestamp 1666464484
transform 1 0 96656 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_854
timestamp 1666464484
transform 1 0 96992 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_918
timestamp 1666464484
transform 1 0 104160 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_922
timestamp 1666464484
transform 1 0 104608 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_925
timestamp 1666464484
transform 1 0 104944 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_989
timestamp 1666464484
transform 1 0 112112 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_993
timestamp 1666464484
transform 1 0 112560 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_996
timestamp 1666464484
transform 1 0 112896 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1060
timestamp 1666464484
transform 1 0 120064 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1064
timestamp 1666464484
transform 1 0 120512 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1067
timestamp 1666464484
transform 1 0 120848 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1131
timestamp 1666464484
transform 1 0 128016 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1135
timestamp 1666464484
transform 1 0 128464 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1138
timestamp 1666464484
transform 1 0 128800 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1202
timestamp 1666464484
transform 1 0 135968 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1206
timestamp 1666464484
transform 1 0 136416 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1209
timestamp 1666464484
transform 1 0 136752 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1273
timestamp 1666464484
transform 1 0 143920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1277
timestamp 1666464484
transform 1 0 144368 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_1280
timestamp 1666464484
transform 1 0 144704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1288
timestamp 1666464484
transform 1 0 145600 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_1292
timestamp 1666464484
transform 1 0 146048 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_1296
timestamp 1666464484
transform 1 0 146496 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1312
timestamp 1666464484
transform 1 0 148288 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1666464484
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1666464484
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1666464484
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1666464484
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1666464484
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1666464484
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1666464484
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1666464484
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1666464484
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1666464484
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1666464484
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1666464484
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1666464484
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1666464484
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1666464484
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1666464484
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1666464484
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1666464484
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1666464484
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1666464484
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1666464484
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_527
timestamp 1666464484
transform 1 0 60368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1666464484
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1666464484
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_598
timestamp 1666464484
transform 1 0 68320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1666464484
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_605
timestamp 1666464484
transform 1 0 69104 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_669
timestamp 1666464484
transform 1 0 76272 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1666464484
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_676
timestamp 1666464484
transform 1 0 77056 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_740
timestamp 1666464484
transform 1 0 84224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_744
timestamp 1666464484
transform 1 0 84672 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_747
timestamp 1666464484
transform 1 0 85008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_811
timestamp 1666464484
transform 1 0 92176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_815
timestamp 1666464484
transform 1 0 92624 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_818
timestamp 1666464484
transform 1 0 92960 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_882
timestamp 1666464484
transform 1 0 100128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_886
timestamp 1666464484
transform 1 0 100576 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_889
timestamp 1666464484
transform 1 0 100912 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_953
timestamp 1666464484
transform 1 0 108080 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_957
timestamp 1666464484
transform 1 0 108528 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_960
timestamp 1666464484
transform 1 0 108864 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1024
timestamp 1666464484
transform 1 0 116032 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1028
timestamp 1666464484
transform 1 0 116480 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1031
timestamp 1666464484
transform 1 0 116816 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1095
timestamp 1666464484
transform 1 0 123984 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1099
timestamp 1666464484
transform 1 0 124432 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1102
timestamp 1666464484
transform 1 0 124768 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1166
timestamp 1666464484
transform 1 0 131936 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1170
timestamp 1666464484
transform 1 0 132384 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1173
timestamp 1666464484
transform 1 0 132720 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1237
timestamp 1666464484
transform 1 0 139888 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1241
timestamp 1666464484
transform 1 0 140336 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_1244
timestamp 1666464484
transform 1 0 140672 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_1276
timestamp 1666464484
transform 1 0 144256 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_1292
timestamp 1666464484
transform 1 0 146048 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_1296
timestamp 1666464484
transform 1 0 146496 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1312
timestamp 1666464484
transform 1 0 148288 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1666464484
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1666464484
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1666464484
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1666464484
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1666464484
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1666464484
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1666464484
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1666464484
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1666464484
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1666464484
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1666464484
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1666464484
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1666464484
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1666464484
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1666464484
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1666464484
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1666464484
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1666464484
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1666464484
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1666464484
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1666464484
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1666464484
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_563
timestamp 1666464484
transform 1 0 64400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1666464484
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1666464484
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1666464484
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1666464484
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_641
timestamp 1666464484
transform 1 0 73136 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_705
timestamp 1666464484
transform 1 0 80304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_709
timestamp 1666464484
transform 1 0 80752 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_712
timestamp 1666464484
transform 1 0 81088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_776
timestamp 1666464484
transform 1 0 88256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_780
timestamp 1666464484
transform 1 0 88704 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_783
timestamp 1666464484
transform 1 0 89040 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_847
timestamp 1666464484
transform 1 0 96208 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_851
timestamp 1666464484
transform 1 0 96656 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_854
timestamp 1666464484
transform 1 0 96992 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_918
timestamp 1666464484
transform 1 0 104160 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_922
timestamp 1666464484
transform 1 0 104608 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_925
timestamp 1666464484
transform 1 0 104944 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_989
timestamp 1666464484
transform 1 0 112112 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_993
timestamp 1666464484
transform 1 0 112560 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_996
timestamp 1666464484
transform 1 0 112896 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1060
timestamp 1666464484
transform 1 0 120064 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1064
timestamp 1666464484
transform 1 0 120512 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1067
timestamp 1666464484
transform 1 0 120848 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1131
timestamp 1666464484
transform 1 0 128016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1135
timestamp 1666464484
transform 1 0 128464 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1138
timestamp 1666464484
transform 1 0 128800 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1202
timestamp 1666464484
transform 1 0 135968 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1206
timestamp 1666464484
transform 1 0 136416 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1209
timestamp 1666464484
transform 1 0 136752 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1273
timestamp 1666464484
transform 1 0 143920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1277
timestamp 1666464484
transform 1 0 144368 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_1280
timestamp 1666464484
transform 1 0 144704 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1288
timestamp 1666464484
transform 1 0 145600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_1292
timestamp 1666464484
transform 1 0 146048 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_1296
timestamp 1666464484
transform 1 0 146496 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1312
timestamp 1666464484
transform 1 0 148288 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1666464484
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1666464484
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1666464484
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1666464484
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1666464484
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1666464484
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1666464484
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1666464484
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1666464484
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1666464484
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1666464484
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1666464484
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1666464484
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1666464484
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1666464484
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1666464484
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1666464484
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1666464484
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1666464484
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1666464484
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1666464484
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_527
timestamp 1666464484
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1666464484
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1666464484
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_598
timestamp 1666464484
transform 1 0 68320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1666464484
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605
timestamp 1666464484
transform 1 0 69104 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_669
timestamp 1666464484
transform 1 0 76272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1666464484
transform 1 0 76720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_676
timestamp 1666464484
transform 1 0 77056 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_740
timestamp 1666464484
transform 1 0 84224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_744
timestamp 1666464484
transform 1 0 84672 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_747
timestamp 1666464484
transform 1 0 85008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_811
timestamp 1666464484
transform 1 0 92176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_815
timestamp 1666464484
transform 1 0 92624 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_818
timestamp 1666464484
transform 1 0 92960 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_882
timestamp 1666464484
transform 1 0 100128 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_886
timestamp 1666464484
transform 1 0 100576 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_889
timestamp 1666464484
transform 1 0 100912 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_953
timestamp 1666464484
transform 1 0 108080 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_957
timestamp 1666464484
transform 1 0 108528 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_960
timestamp 1666464484
transform 1 0 108864 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1024
timestamp 1666464484
transform 1 0 116032 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1028
timestamp 1666464484
transform 1 0 116480 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1031
timestamp 1666464484
transform 1 0 116816 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1095
timestamp 1666464484
transform 1 0 123984 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1099
timestamp 1666464484
transform 1 0 124432 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1102
timestamp 1666464484
transform 1 0 124768 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1166
timestamp 1666464484
transform 1 0 131936 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1170
timestamp 1666464484
transform 1 0 132384 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1173
timestamp 1666464484
transform 1 0 132720 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1237
timestamp 1666464484
transform 1 0 139888 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1241
timestamp 1666464484
transform 1 0 140336 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_1244
timestamp 1666464484
transform 1 0 140672 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_1276
timestamp 1666464484
transform 1 0 144256 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_1292
timestamp 1666464484
transform 1 0 146048 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_1296
timestamp 1666464484
transform 1 0 146496 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1312
timestamp 1666464484
transform 1 0 148288 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1666464484
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1666464484
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1666464484
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1666464484
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1666464484
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1666464484
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1666464484
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1666464484
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1666464484
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1666464484
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1666464484
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1666464484
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1666464484
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1666464484
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1666464484
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1666464484
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1666464484
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1666464484
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1666464484
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1666464484
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1666464484
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1666464484
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_563
timestamp 1666464484
transform 1 0 64400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1666464484
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1666464484
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1666464484
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1666464484
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_641
timestamp 1666464484
transform 1 0 73136 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_705
timestamp 1666464484
transform 1 0 80304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_709
timestamp 1666464484
transform 1 0 80752 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_712
timestamp 1666464484
transform 1 0 81088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_776
timestamp 1666464484
transform 1 0 88256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_780
timestamp 1666464484
transform 1 0 88704 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_783
timestamp 1666464484
transform 1 0 89040 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_847
timestamp 1666464484
transform 1 0 96208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_851
timestamp 1666464484
transform 1 0 96656 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_854
timestamp 1666464484
transform 1 0 96992 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_918
timestamp 1666464484
transform 1 0 104160 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_922
timestamp 1666464484
transform 1 0 104608 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_925
timestamp 1666464484
transform 1 0 104944 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_989
timestamp 1666464484
transform 1 0 112112 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_993
timestamp 1666464484
transform 1 0 112560 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_996
timestamp 1666464484
transform 1 0 112896 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1060
timestamp 1666464484
transform 1 0 120064 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1064
timestamp 1666464484
transform 1 0 120512 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1067
timestamp 1666464484
transform 1 0 120848 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1131
timestamp 1666464484
transform 1 0 128016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1135
timestamp 1666464484
transform 1 0 128464 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1138
timestamp 1666464484
transform 1 0 128800 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1202
timestamp 1666464484
transform 1 0 135968 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1206
timestamp 1666464484
transform 1 0 136416 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1209
timestamp 1666464484
transform 1 0 136752 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1273
timestamp 1666464484
transform 1 0 143920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1277
timestamp 1666464484
transform 1 0 144368 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_1280
timestamp 1666464484
transform 1 0 144704 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1288
timestamp 1666464484
transform 1 0 145600 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_1292
timestamp 1666464484
transform 1 0 146048 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_1296
timestamp 1666464484
transform 1 0 146496 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1312
timestamp 1666464484
transform 1 0 148288 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1666464484
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1666464484
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1666464484
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1666464484
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1666464484
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1666464484
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1666464484
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1666464484
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1666464484
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1666464484
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1666464484
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1666464484
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1666464484
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1666464484
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1666464484
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1666464484
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1666464484
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1666464484
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1666464484
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1666464484
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1666464484
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_527
timestamp 1666464484
transform 1 0 60368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1666464484
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1666464484
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1666464484
transform 1 0 68320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1666464484
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1666464484
transform 1 0 69104 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_669
timestamp 1666464484
transform 1 0 76272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1666464484
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_676
timestamp 1666464484
transform 1 0 77056 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_740
timestamp 1666464484
transform 1 0 84224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_744
timestamp 1666464484
transform 1 0 84672 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_747
timestamp 1666464484
transform 1 0 85008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_811
timestamp 1666464484
transform 1 0 92176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_815
timestamp 1666464484
transform 1 0 92624 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_818
timestamp 1666464484
transform 1 0 92960 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_882
timestamp 1666464484
transform 1 0 100128 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_886
timestamp 1666464484
transform 1 0 100576 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_889
timestamp 1666464484
transform 1 0 100912 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_953
timestamp 1666464484
transform 1 0 108080 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_957
timestamp 1666464484
transform 1 0 108528 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_960
timestamp 1666464484
transform 1 0 108864 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1024
timestamp 1666464484
transform 1 0 116032 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1028
timestamp 1666464484
transform 1 0 116480 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1031
timestamp 1666464484
transform 1 0 116816 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1095
timestamp 1666464484
transform 1 0 123984 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1099
timestamp 1666464484
transform 1 0 124432 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1102
timestamp 1666464484
transform 1 0 124768 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1166
timestamp 1666464484
transform 1 0 131936 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1170
timestamp 1666464484
transform 1 0 132384 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1173
timestamp 1666464484
transform 1 0 132720 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1237
timestamp 1666464484
transform 1 0 139888 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1241
timestamp 1666464484
transform 1 0 140336 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_1244
timestamp 1666464484
transform 1 0 140672 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_1276
timestamp 1666464484
transform 1 0 144256 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_1292
timestamp 1666464484
transform 1 0 146048 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_1296
timestamp 1666464484
transform 1 0 146496 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1312
timestamp 1666464484
transform 1 0 148288 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1666464484
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1666464484
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1666464484
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1666464484
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1666464484
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1666464484
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1666464484
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1666464484
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1666464484
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1666464484
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1666464484
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1666464484
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1666464484
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1666464484
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1666464484
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1666464484
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1666464484
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1666464484
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1666464484
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1666464484
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1666464484
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1666464484
transform 1 0 57232 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_563
timestamp 1666464484
transform 1 0 64400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1666464484
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1666464484
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1666464484
transform 1 0 72352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1666464484
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_641
timestamp 1666464484
transform 1 0 73136 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_705
timestamp 1666464484
transform 1 0 80304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_709
timestamp 1666464484
transform 1 0 80752 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_712
timestamp 1666464484
transform 1 0 81088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_776
timestamp 1666464484
transform 1 0 88256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_780
timestamp 1666464484
transform 1 0 88704 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_783
timestamp 1666464484
transform 1 0 89040 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_847
timestamp 1666464484
transform 1 0 96208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_851
timestamp 1666464484
transform 1 0 96656 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_854
timestamp 1666464484
transform 1 0 96992 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_918
timestamp 1666464484
transform 1 0 104160 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_922
timestamp 1666464484
transform 1 0 104608 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_925
timestamp 1666464484
transform 1 0 104944 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_989
timestamp 1666464484
transform 1 0 112112 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_993
timestamp 1666464484
transform 1 0 112560 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_996
timestamp 1666464484
transform 1 0 112896 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1060
timestamp 1666464484
transform 1 0 120064 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1064
timestamp 1666464484
transform 1 0 120512 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1067
timestamp 1666464484
transform 1 0 120848 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1131
timestamp 1666464484
transform 1 0 128016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1135
timestamp 1666464484
transform 1 0 128464 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1138
timestamp 1666464484
transform 1 0 128800 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1202
timestamp 1666464484
transform 1 0 135968 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1206
timestamp 1666464484
transform 1 0 136416 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1209
timestamp 1666464484
transform 1 0 136752 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1273
timestamp 1666464484
transform 1 0 143920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1277
timestamp 1666464484
transform 1 0 144368 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_1280
timestamp 1666464484
transform 1 0 144704 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1312
timestamp 1666464484
transform 1 0 148288 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1666464484
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1666464484
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1666464484
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1666464484
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1666464484
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1666464484
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1666464484
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1666464484
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1666464484
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1666464484
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1666464484
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1666464484
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1666464484
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1666464484
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1666464484
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1666464484
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1666464484
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1666464484
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1666464484
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1666464484
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1666464484
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1666464484
transform 1 0 60368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1666464484
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1666464484
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1666464484
transform 1 0 68320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1666464484
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1666464484
transform 1 0 69104 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_669
timestamp 1666464484
transform 1 0 76272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1666464484
transform 1 0 76720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_676
timestamp 1666464484
transform 1 0 77056 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_740
timestamp 1666464484
transform 1 0 84224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_744
timestamp 1666464484
transform 1 0 84672 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_747
timestamp 1666464484
transform 1 0 85008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_811
timestamp 1666464484
transform 1 0 92176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_815
timestamp 1666464484
transform 1 0 92624 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_818
timestamp 1666464484
transform 1 0 92960 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_882
timestamp 1666464484
transform 1 0 100128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_886
timestamp 1666464484
transform 1 0 100576 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_889
timestamp 1666464484
transform 1 0 100912 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_953
timestamp 1666464484
transform 1 0 108080 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_957
timestamp 1666464484
transform 1 0 108528 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_960
timestamp 1666464484
transform 1 0 108864 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1024
timestamp 1666464484
transform 1 0 116032 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1028
timestamp 1666464484
transform 1 0 116480 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1031
timestamp 1666464484
transform 1 0 116816 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1095
timestamp 1666464484
transform 1 0 123984 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1099
timestamp 1666464484
transform 1 0 124432 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1102
timestamp 1666464484
transform 1 0 124768 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1166
timestamp 1666464484
transform 1 0 131936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1170
timestamp 1666464484
transform 1 0 132384 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1173
timestamp 1666464484
transform 1 0 132720 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1237
timestamp 1666464484
transform 1 0 139888 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1241
timestamp 1666464484
transform 1 0 140336 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_1244
timestamp 1666464484
transform 1 0 140672 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_1276
timestamp 1666464484
transform 1 0 144256 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_1292
timestamp 1666464484
transform 1 0 146048 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_1296
timestamp 1666464484
transform 1 0 146496 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1312
timestamp 1666464484
transform 1 0 148288 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1666464484
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1666464484
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1666464484
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1666464484
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1666464484
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1666464484
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1666464484
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1666464484
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1666464484
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1666464484
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1666464484
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1666464484
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1666464484
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1666464484
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1666464484
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1666464484
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1666464484
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1666464484
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1666464484
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1666464484
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1666464484
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1666464484
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1666464484
transform 1 0 64400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1666464484
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1666464484
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1666464484
transform 1 0 72352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1666464484
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_641
timestamp 1666464484
transform 1 0 73136 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_705
timestamp 1666464484
transform 1 0 80304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_709
timestamp 1666464484
transform 1 0 80752 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_712
timestamp 1666464484
transform 1 0 81088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_776
timestamp 1666464484
transform 1 0 88256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_780
timestamp 1666464484
transform 1 0 88704 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_783
timestamp 1666464484
transform 1 0 89040 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_847
timestamp 1666464484
transform 1 0 96208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_851
timestamp 1666464484
transform 1 0 96656 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_854
timestamp 1666464484
transform 1 0 96992 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_918
timestamp 1666464484
transform 1 0 104160 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_922
timestamp 1666464484
transform 1 0 104608 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_925
timestamp 1666464484
transform 1 0 104944 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_989
timestamp 1666464484
transform 1 0 112112 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_993
timestamp 1666464484
transform 1 0 112560 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_996
timestamp 1666464484
transform 1 0 112896 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1060
timestamp 1666464484
transform 1 0 120064 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1064
timestamp 1666464484
transform 1 0 120512 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1067
timestamp 1666464484
transform 1 0 120848 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1131
timestamp 1666464484
transform 1 0 128016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1135
timestamp 1666464484
transform 1 0 128464 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1138
timestamp 1666464484
transform 1 0 128800 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1202
timestamp 1666464484
transform 1 0 135968 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1206
timestamp 1666464484
transform 1 0 136416 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1209
timestamp 1666464484
transform 1 0 136752 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1273
timestamp 1666464484
transform 1 0 143920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1277
timestamp 1666464484
transform 1 0 144368 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_1280
timestamp 1666464484
transform 1 0 144704 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1288
timestamp 1666464484
transform 1 0 145600 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_1292
timestamp 1666464484
transform 1 0 146048 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_1296
timestamp 1666464484
transform 1 0 146496 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1312
timestamp 1666464484
transform 1 0 148288 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1666464484
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1666464484
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1666464484
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1666464484
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1666464484
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1666464484
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1666464484
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1666464484
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1666464484
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1666464484
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1666464484
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1666464484
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1666464484
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1666464484
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1666464484
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1666464484
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1666464484
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1666464484
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1666464484
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1666464484
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1666464484
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1666464484
transform 1 0 60368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1666464484
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1666464484
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1666464484
transform 1 0 68320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1666464484
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1666464484
transform 1 0 69104 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_669
timestamp 1666464484
transform 1 0 76272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1666464484
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_676
timestamp 1666464484
transform 1 0 77056 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_740
timestamp 1666464484
transform 1 0 84224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_744
timestamp 1666464484
transform 1 0 84672 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_747
timestamp 1666464484
transform 1 0 85008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_811
timestamp 1666464484
transform 1 0 92176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_815
timestamp 1666464484
transform 1 0 92624 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_818
timestamp 1666464484
transform 1 0 92960 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_882
timestamp 1666464484
transform 1 0 100128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_886
timestamp 1666464484
transform 1 0 100576 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_889
timestamp 1666464484
transform 1 0 100912 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_953
timestamp 1666464484
transform 1 0 108080 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_957
timestamp 1666464484
transform 1 0 108528 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_960
timestamp 1666464484
transform 1 0 108864 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1024
timestamp 1666464484
transform 1 0 116032 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1028
timestamp 1666464484
transform 1 0 116480 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1031
timestamp 1666464484
transform 1 0 116816 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1095
timestamp 1666464484
transform 1 0 123984 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1099
timestamp 1666464484
transform 1 0 124432 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1102
timestamp 1666464484
transform 1 0 124768 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1166
timestamp 1666464484
transform 1 0 131936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1170
timestamp 1666464484
transform 1 0 132384 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1173
timestamp 1666464484
transform 1 0 132720 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1237
timestamp 1666464484
transform 1 0 139888 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1241
timestamp 1666464484
transform 1 0 140336 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_1244
timestamp 1666464484
transform 1 0 140672 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_1276
timestamp 1666464484
transform 1 0 144256 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_1292
timestamp 1666464484
transform 1 0 146048 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_1296
timestamp 1666464484
transform 1 0 146496 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1312
timestamp 1666464484
transform 1 0 148288 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1666464484
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1666464484
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1666464484
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1666464484
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1666464484
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1666464484
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1666464484
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1666464484
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1666464484
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1666464484
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1666464484
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1666464484
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1666464484
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1666464484
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1666464484
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1666464484
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1666464484
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1666464484
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1666464484
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1666464484
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1666464484
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1666464484
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1666464484
transform 1 0 64400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1666464484
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1666464484
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1666464484
transform 1 0 72352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1666464484
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_641
timestamp 1666464484
transform 1 0 73136 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_705
timestamp 1666464484
transform 1 0 80304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_709
timestamp 1666464484
transform 1 0 80752 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_712
timestamp 1666464484
transform 1 0 81088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_776
timestamp 1666464484
transform 1 0 88256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_780
timestamp 1666464484
transform 1 0 88704 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_783
timestamp 1666464484
transform 1 0 89040 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_847
timestamp 1666464484
transform 1 0 96208 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_851
timestamp 1666464484
transform 1 0 96656 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_854
timestamp 1666464484
transform 1 0 96992 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_918
timestamp 1666464484
transform 1 0 104160 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_922
timestamp 1666464484
transform 1 0 104608 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_925
timestamp 1666464484
transform 1 0 104944 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_989
timestamp 1666464484
transform 1 0 112112 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_993
timestamp 1666464484
transform 1 0 112560 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_996
timestamp 1666464484
transform 1 0 112896 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1060
timestamp 1666464484
transform 1 0 120064 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1064
timestamp 1666464484
transform 1 0 120512 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1067
timestamp 1666464484
transform 1 0 120848 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1131
timestamp 1666464484
transform 1 0 128016 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1135
timestamp 1666464484
transform 1 0 128464 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1138
timestamp 1666464484
transform 1 0 128800 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1202
timestamp 1666464484
transform 1 0 135968 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1206
timestamp 1666464484
transform 1 0 136416 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1209
timestamp 1666464484
transform 1 0 136752 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1273
timestamp 1666464484
transform 1 0 143920 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1277
timestamp 1666464484
transform 1 0 144368 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_1280
timestamp 1666464484
transform 1 0 144704 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1288
timestamp 1666464484
transform 1 0 145600 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_1292
timestamp 1666464484
transform 1 0 146048 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_1296
timestamp 1666464484
transform 1 0 146496 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1312
timestamp 1666464484
transform 1 0 148288 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1666464484
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1666464484
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1666464484
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1666464484
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1666464484
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1666464484
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1666464484
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1666464484
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1666464484
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1666464484
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1666464484
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1666464484
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1666464484
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1666464484
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1666464484
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1666464484
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1666464484
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1666464484
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1666464484
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1666464484
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1666464484
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1666464484
transform 1 0 60368 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1666464484
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1666464484
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1666464484
transform 1 0 68320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1666464484
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_605
timestamp 1666464484
transform 1 0 69104 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_669
timestamp 1666464484
transform 1 0 76272 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1666464484
transform 1 0 76720 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_676
timestamp 1666464484
transform 1 0 77056 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_740
timestamp 1666464484
transform 1 0 84224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_744
timestamp 1666464484
transform 1 0 84672 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_747
timestamp 1666464484
transform 1 0 85008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_811
timestamp 1666464484
transform 1 0 92176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_815
timestamp 1666464484
transform 1 0 92624 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_818
timestamp 1666464484
transform 1 0 92960 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_882
timestamp 1666464484
transform 1 0 100128 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_886
timestamp 1666464484
transform 1 0 100576 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_889
timestamp 1666464484
transform 1 0 100912 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_953
timestamp 1666464484
transform 1 0 108080 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_957
timestamp 1666464484
transform 1 0 108528 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_960
timestamp 1666464484
transform 1 0 108864 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1024
timestamp 1666464484
transform 1 0 116032 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1028
timestamp 1666464484
transform 1 0 116480 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1031
timestamp 1666464484
transform 1 0 116816 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1095
timestamp 1666464484
transform 1 0 123984 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1099
timestamp 1666464484
transform 1 0 124432 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1102
timestamp 1666464484
transform 1 0 124768 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1166
timestamp 1666464484
transform 1 0 131936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1170
timestamp 1666464484
transform 1 0 132384 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1173
timestamp 1666464484
transform 1 0 132720 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1237
timestamp 1666464484
transform 1 0 139888 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1241
timestamp 1666464484
transform 1 0 140336 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_1244
timestamp 1666464484
transform 1 0 140672 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_1276
timestamp 1666464484
transform 1 0 144256 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_1292
timestamp 1666464484
transform 1 0 146048 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_1296
timestamp 1666464484
transform 1 0 146496 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1312
timestamp 1666464484
transform 1 0 148288 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1666464484
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1666464484
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1666464484
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1666464484
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1666464484
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1666464484
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1666464484
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1666464484
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1666464484
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1666464484
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1666464484
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1666464484
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1666464484
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1666464484
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1666464484
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1666464484
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1666464484
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1666464484
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1666464484
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1666464484
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1666464484
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1666464484
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1666464484
transform 1 0 64400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1666464484
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1666464484
transform 1 0 65184 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1666464484
transform 1 0 72352 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1666464484
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_641
timestamp 1666464484
transform 1 0 73136 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_705
timestamp 1666464484
transform 1 0 80304 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_709
timestamp 1666464484
transform 1 0 80752 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_712
timestamp 1666464484
transform 1 0 81088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_776
timestamp 1666464484
transform 1 0 88256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_780
timestamp 1666464484
transform 1 0 88704 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_783
timestamp 1666464484
transform 1 0 89040 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_847
timestamp 1666464484
transform 1 0 96208 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_851
timestamp 1666464484
transform 1 0 96656 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_854
timestamp 1666464484
transform 1 0 96992 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_918
timestamp 1666464484
transform 1 0 104160 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_922
timestamp 1666464484
transform 1 0 104608 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_925
timestamp 1666464484
transform 1 0 104944 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_989
timestamp 1666464484
transform 1 0 112112 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_993
timestamp 1666464484
transform 1 0 112560 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_996
timestamp 1666464484
transform 1 0 112896 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1060
timestamp 1666464484
transform 1 0 120064 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1064
timestamp 1666464484
transform 1 0 120512 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1067
timestamp 1666464484
transform 1 0 120848 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1131
timestamp 1666464484
transform 1 0 128016 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1135
timestamp 1666464484
transform 1 0 128464 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1138
timestamp 1666464484
transform 1 0 128800 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1202
timestamp 1666464484
transform 1 0 135968 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1206
timestamp 1666464484
transform 1 0 136416 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1209
timestamp 1666464484
transform 1 0 136752 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1273
timestamp 1666464484
transform 1 0 143920 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1277
timestamp 1666464484
transform 1 0 144368 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_1280
timestamp 1666464484
transform 1 0 144704 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1288
timestamp 1666464484
transform 1 0 145600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_1292
timestamp 1666464484
transform 1 0 146048 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_1296
timestamp 1666464484
transform 1 0 146496 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1312
timestamp 1666464484
transform 1 0 148288 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1666464484
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1666464484
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1666464484
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1666464484
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1666464484
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1666464484
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1666464484
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1666464484
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1666464484
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1666464484
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1666464484
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1666464484
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1666464484
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1666464484
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1666464484
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1666464484
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1666464484
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1666464484
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1666464484
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1666464484
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1666464484
transform 1 0 53200 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1666464484
transform 1 0 60368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1666464484
transform 1 0 60816 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1666464484
transform 1 0 61152 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_598
timestamp 1666464484
transform 1 0 68320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1666464484
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1666464484
transform 1 0 69104 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_669
timestamp 1666464484
transform 1 0 76272 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1666464484
transform 1 0 76720 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_676
timestamp 1666464484
transform 1 0 77056 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_740
timestamp 1666464484
transform 1 0 84224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_744
timestamp 1666464484
transform 1 0 84672 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_747
timestamp 1666464484
transform 1 0 85008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_811
timestamp 1666464484
transform 1 0 92176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_815
timestamp 1666464484
transform 1 0 92624 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_818
timestamp 1666464484
transform 1 0 92960 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_882
timestamp 1666464484
transform 1 0 100128 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_886
timestamp 1666464484
transform 1 0 100576 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_889
timestamp 1666464484
transform 1 0 100912 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_953
timestamp 1666464484
transform 1 0 108080 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_957
timestamp 1666464484
transform 1 0 108528 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_960
timestamp 1666464484
transform 1 0 108864 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1024
timestamp 1666464484
transform 1 0 116032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1028
timestamp 1666464484
transform 1 0 116480 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1031
timestamp 1666464484
transform 1 0 116816 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1095
timestamp 1666464484
transform 1 0 123984 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1099
timestamp 1666464484
transform 1 0 124432 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1102
timestamp 1666464484
transform 1 0 124768 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1166
timestamp 1666464484
transform 1 0 131936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1170
timestamp 1666464484
transform 1 0 132384 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1173
timestamp 1666464484
transform 1 0 132720 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1237
timestamp 1666464484
transform 1 0 139888 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1241
timestamp 1666464484
transform 1 0 140336 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_1244
timestamp 1666464484
transform 1 0 140672 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_1276
timestamp 1666464484
transform 1 0 144256 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_1292
timestamp 1666464484
transform 1 0 146048 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_1296
timestamp 1666464484
transform 1 0 146496 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1312
timestamp 1666464484
transform 1 0 148288 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1666464484
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1666464484
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1666464484
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1666464484
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1666464484
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1666464484
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1666464484
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1666464484
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1666464484
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1666464484
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1666464484
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1666464484
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1666464484
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1666464484
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1666464484
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1666464484
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1666464484
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1666464484
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1666464484
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1666464484
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1666464484
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_499
timestamp 1666464484
transform 1 0 57232 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_563
timestamp 1666464484
transform 1 0 64400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1666464484
transform 1 0 64848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1666464484
transform 1 0 65184 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_634
timestamp 1666464484
transform 1 0 72352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1666464484
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_641
timestamp 1666464484
transform 1 0 73136 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_705
timestamp 1666464484
transform 1 0 80304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_709
timestamp 1666464484
transform 1 0 80752 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_712
timestamp 1666464484
transform 1 0 81088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_776
timestamp 1666464484
transform 1 0 88256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_780
timestamp 1666464484
transform 1 0 88704 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_783
timestamp 1666464484
transform 1 0 89040 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_847
timestamp 1666464484
transform 1 0 96208 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_851
timestamp 1666464484
transform 1 0 96656 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_854
timestamp 1666464484
transform 1 0 96992 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_918
timestamp 1666464484
transform 1 0 104160 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_922
timestamp 1666464484
transform 1 0 104608 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_925
timestamp 1666464484
transform 1 0 104944 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_989
timestamp 1666464484
transform 1 0 112112 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_993
timestamp 1666464484
transform 1 0 112560 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_996
timestamp 1666464484
transform 1 0 112896 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1060
timestamp 1666464484
transform 1 0 120064 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1064
timestamp 1666464484
transform 1 0 120512 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1067
timestamp 1666464484
transform 1 0 120848 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1131
timestamp 1666464484
transform 1 0 128016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1135
timestamp 1666464484
transform 1 0 128464 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1138
timestamp 1666464484
transform 1 0 128800 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1202
timestamp 1666464484
transform 1 0 135968 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1206
timestamp 1666464484
transform 1 0 136416 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1209
timestamp 1666464484
transform 1 0 136752 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1273
timestamp 1666464484
transform 1 0 143920 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1277
timestamp 1666464484
transform 1 0 144368 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_1280
timestamp 1666464484
transform 1 0 144704 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1312
timestamp 1666464484
transform 1 0 148288 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1666464484
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1666464484
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1666464484
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1666464484
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1666464484
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1666464484
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1666464484
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1666464484
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1666464484
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1666464484
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1666464484
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1666464484
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1666464484
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1666464484
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1666464484
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1666464484
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1666464484
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1666464484
transform 1 0 45248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1666464484
transform 1 0 52416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1666464484
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_463
timestamp 1666464484
transform 1 0 53200 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_527
timestamp 1666464484
transform 1 0 60368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1666464484
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_534
timestamp 1666464484
transform 1 0 61152 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_598
timestamp 1666464484
transform 1 0 68320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1666464484
transform 1 0 68768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_605
timestamp 1666464484
transform 1 0 69104 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_669
timestamp 1666464484
transform 1 0 76272 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1666464484
transform 1 0 76720 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_676
timestamp 1666464484
transform 1 0 77056 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_740
timestamp 1666464484
transform 1 0 84224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_744
timestamp 1666464484
transform 1 0 84672 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_747
timestamp 1666464484
transform 1 0 85008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_811
timestamp 1666464484
transform 1 0 92176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_815
timestamp 1666464484
transform 1 0 92624 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_818
timestamp 1666464484
transform 1 0 92960 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_882
timestamp 1666464484
transform 1 0 100128 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_886
timestamp 1666464484
transform 1 0 100576 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_889
timestamp 1666464484
transform 1 0 100912 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_953
timestamp 1666464484
transform 1 0 108080 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_957
timestamp 1666464484
transform 1 0 108528 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_960
timestamp 1666464484
transform 1 0 108864 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1024
timestamp 1666464484
transform 1 0 116032 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1028
timestamp 1666464484
transform 1 0 116480 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1031
timestamp 1666464484
transform 1 0 116816 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1095
timestamp 1666464484
transform 1 0 123984 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1099
timestamp 1666464484
transform 1 0 124432 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1102
timestamp 1666464484
transform 1 0 124768 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1166
timestamp 1666464484
transform 1 0 131936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1170
timestamp 1666464484
transform 1 0 132384 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1173
timestamp 1666464484
transform 1 0 132720 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1237
timestamp 1666464484
transform 1 0 139888 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1241
timestamp 1666464484
transform 1 0 140336 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_1244
timestamp 1666464484
transform 1 0 140672 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_1276
timestamp 1666464484
transform 1 0 144256 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1292
timestamp 1666464484
transform 1 0 146048 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1296
timestamp 1666464484
transform 1 0 146496 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1312
timestamp 1666464484
transform 1 0 148288 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1666464484
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1666464484
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1666464484
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1666464484
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1666464484
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1666464484
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1666464484
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1666464484
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1666464484
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1666464484
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1666464484
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1666464484
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1666464484
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1666464484
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1666464484
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1666464484
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1666464484
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1666464484
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1666464484
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1666464484
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1666464484
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_499
timestamp 1666464484
transform 1 0 57232 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_563
timestamp 1666464484
transform 1 0 64400 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1666464484
transform 1 0 64848 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_570
timestamp 1666464484
transform 1 0 65184 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_634
timestamp 1666464484
transform 1 0 72352 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1666464484
transform 1 0 72800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_641
timestamp 1666464484
transform 1 0 73136 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_705
timestamp 1666464484
transform 1 0 80304 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_709
timestamp 1666464484
transform 1 0 80752 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_712
timestamp 1666464484
transform 1 0 81088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_776
timestamp 1666464484
transform 1 0 88256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_780
timestamp 1666464484
transform 1 0 88704 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_783
timestamp 1666464484
transform 1 0 89040 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_847
timestamp 1666464484
transform 1 0 96208 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_851
timestamp 1666464484
transform 1 0 96656 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_854
timestamp 1666464484
transform 1 0 96992 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_918
timestamp 1666464484
transform 1 0 104160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_922
timestamp 1666464484
transform 1 0 104608 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_925
timestamp 1666464484
transform 1 0 104944 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_989
timestamp 1666464484
transform 1 0 112112 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_993
timestamp 1666464484
transform 1 0 112560 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_996
timestamp 1666464484
transform 1 0 112896 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1060
timestamp 1666464484
transform 1 0 120064 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1064
timestamp 1666464484
transform 1 0 120512 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1067
timestamp 1666464484
transform 1 0 120848 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1131
timestamp 1666464484
transform 1 0 128016 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1135
timestamp 1666464484
transform 1 0 128464 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1138
timestamp 1666464484
transform 1 0 128800 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1202
timestamp 1666464484
transform 1 0 135968 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1206
timestamp 1666464484
transform 1 0 136416 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1209
timestamp 1666464484
transform 1 0 136752 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1273
timestamp 1666464484
transform 1 0 143920 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1277
timestamp 1666464484
transform 1 0 144368 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1280
timestamp 1666464484
transform 1 0 144704 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1284
timestamp 1666464484
transform 1 0 145152 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1288
timestamp 1666464484
transform 1 0 145600 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1292
timestamp 1666464484
transform 1 0 146048 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1296
timestamp 1666464484
transform 1 0 146496 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1312
timestamp 1666464484
transform 1 0 148288 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1666464484
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1666464484
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1666464484
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1666464484
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1666464484
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1666464484
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1666464484
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1666464484
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1666464484
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1666464484
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1666464484
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1666464484
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1666464484
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1666464484
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1666464484
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1666464484
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1666464484
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1666464484
transform 1 0 45248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1666464484
transform 1 0 52416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1666464484
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_463
timestamp 1666464484
transform 1 0 53200 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_527
timestamp 1666464484
transform 1 0 60368 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_534
timestamp 1666464484
transform 1 0 61152 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_598
timestamp 1666464484
transform 1 0 68320 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1666464484
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_605
timestamp 1666464484
transform 1 0 69104 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_669
timestamp 1666464484
transform 1 0 76272 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1666464484
transform 1 0 76720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_676
timestamp 1666464484
transform 1 0 77056 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_740
timestamp 1666464484
transform 1 0 84224 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_744
timestamp 1666464484
transform 1 0 84672 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_747
timestamp 1666464484
transform 1 0 85008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_811
timestamp 1666464484
transform 1 0 92176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_815
timestamp 1666464484
transform 1 0 92624 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_818
timestamp 1666464484
transform 1 0 92960 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_882
timestamp 1666464484
transform 1 0 100128 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_886
timestamp 1666464484
transform 1 0 100576 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_889
timestamp 1666464484
transform 1 0 100912 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_953
timestamp 1666464484
transform 1 0 108080 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_957
timestamp 1666464484
transform 1 0 108528 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_960
timestamp 1666464484
transform 1 0 108864 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1024
timestamp 1666464484
transform 1 0 116032 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1028
timestamp 1666464484
transform 1 0 116480 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1031
timestamp 1666464484
transform 1 0 116816 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1095
timestamp 1666464484
transform 1 0 123984 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1099
timestamp 1666464484
transform 1 0 124432 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1102
timestamp 1666464484
transform 1 0 124768 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1166
timestamp 1666464484
transform 1 0 131936 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1170
timestamp 1666464484
transform 1 0 132384 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1173
timestamp 1666464484
transform 1 0 132720 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1237
timestamp 1666464484
transform 1 0 139888 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1241
timestamp 1666464484
transform 1 0 140336 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_1244
timestamp 1666464484
transform 1 0 140672 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1276
timestamp 1666464484
transform 1 0 144256 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1280
timestamp 1666464484
transform 1 0 144704 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1296
timestamp 1666464484
transform 1 0 146496 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1312
timestamp 1666464484
transform 1 0 148288 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1666464484
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1666464484
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1666464484
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1666464484
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1666464484
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1666464484
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1666464484
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1666464484
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1666464484
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1666464484
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1666464484
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1666464484
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1666464484
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1666464484
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1666464484
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1666464484
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1666464484
transform 1 0 48496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1666464484
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1666464484
transform 1 0 49280 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1666464484
transform 1 0 56448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1666464484
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_499
timestamp 1666464484
transform 1 0 57232 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_563
timestamp 1666464484
transform 1 0 64400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1666464484
transform 1 0 64848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_570
timestamp 1666464484
transform 1 0 65184 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_634
timestamp 1666464484
transform 1 0 72352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1666464484
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_641
timestamp 1666464484
transform 1 0 73136 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_705
timestamp 1666464484
transform 1 0 80304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_709
timestamp 1666464484
transform 1 0 80752 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_712
timestamp 1666464484
transform 1 0 81088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_776
timestamp 1666464484
transform 1 0 88256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_780
timestamp 1666464484
transform 1 0 88704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_783
timestamp 1666464484
transform 1 0 89040 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_847
timestamp 1666464484
transform 1 0 96208 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_851
timestamp 1666464484
transform 1 0 96656 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_854
timestamp 1666464484
transform 1 0 96992 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_918
timestamp 1666464484
transform 1 0 104160 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_922
timestamp 1666464484
transform 1 0 104608 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_925
timestamp 1666464484
transform 1 0 104944 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_989
timestamp 1666464484
transform 1 0 112112 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_993
timestamp 1666464484
transform 1 0 112560 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_996
timestamp 1666464484
transform 1 0 112896 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1060
timestamp 1666464484
transform 1 0 120064 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1064
timestamp 1666464484
transform 1 0 120512 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1067
timestamp 1666464484
transform 1 0 120848 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1131
timestamp 1666464484
transform 1 0 128016 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1135
timestamp 1666464484
transform 1 0 128464 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1138
timestamp 1666464484
transform 1 0 128800 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1202
timestamp 1666464484
transform 1 0 135968 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1206
timestamp 1666464484
transform 1 0 136416 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1209
timestamp 1666464484
transform 1 0 136752 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1273
timestamp 1666464484
transform 1 0 143920 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1277
timestamp 1666464484
transform 1 0 144368 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1280
timestamp 1666464484
transform 1 0 144704 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1296
timestamp 1666464484
transform 1 0 146496 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1312
timestamp 1666464484
transform 1 0 148288 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1666464484
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1666464484
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_37
timestamp 1666464484
transform 1 0 5488 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_69
timestamp 1666464484
transform 1 0 9072 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_72
timestamp 1666464484
transform 1 0 9408 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_104
timestamp 1666464484
transform 1 0 12992 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_107
timestamp 1666464484
transform 1 0 13328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 16912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_142
timestamp 1666464484
transform 1 0 17248 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_174
timestamp 1666464484
transform 1 0 20832 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_177
timestamp 1666464484
transform 1 0 21168 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_209
timestamp 1666464484
transform 1 0 24752 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_212
timestamp 1666464484
transform 1 0 25088 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_244
timestamp 1666464484
transform 1 0 28672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_247
timestamp 1666464484
transform 1 0 29008 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_279
timestamp 1666464484
transform 1 0 32592 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_282
timestamp 1666464484
transform 1 0 32928 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_314
timestamp 1666464484
transform 1 0 36512 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_317
timestamp 1666464484
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_349
timestamp 1666464484
transform 1 0 40432 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_352
timestamp 1666464484
transform 1 0 40768 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_384
timestamp 1666464484
transform 1 0 44352 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_387
timestamp 1666464484
transform 1 0 44688 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_419
timestamp 1666464484
transform 1 0 48272 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_422
timestamp 1666464484
transform 1 0 48608 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_454
timestamp 1666464484
transform 1 0 52192 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_457
timestamp 1666464484
transform 1 0 52528 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_489
timestamp 1666464484
transform 1 0 56112 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_492
timestamp 1666464484
transform 1 0 56448 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_524
timestamp 1666464484
transform 1 0 60032 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_527
timestamp 1666464484
transform 1 0 60368 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_559
timestamp 1666464484
transform 1 0 63952 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_562
timestamp 1666464484
transform 1 0 64288 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_594
timestamp 1666464484
transform 1 0 67872 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_597
timestamp 1666464484
transform 1 0 68208 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_629
timestamp 1666464484
transform 1 0 71792 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_632
timestamp 1666464484
transform 1 0 72128 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_664
timestamp 1666464484
transform 1 0 75712 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_667
timestamp 1666464484
transform 1 0 76048 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_699
timestamp 1666464484
transform 1 0 79632 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_702
timestamp 1666464484
transform 1 0 79968 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_734
timestamp 1666464484
transform 1 0 83552 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_737
timestamp 1666464484
transform 1 0 83888 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_769
timestamp 1666464484
transform 1 0 87472 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_772
timestamp 1666464484
transform 1 0 87808 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_804
timestamp 1666464484
transform 1 0 91392 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_807
timestamp 1666464484
transform 1 0 91728 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_839
timestamp 1666464484
transform 1 0 95312 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_842
timestamp 1666464484
transform 1 0 95648 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_874
timestamp 1666464484
transform 1 0 99232 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_877
timestamp 1666464484
transform 1 0 99568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_909
timestamp 1666464484
transform 1 0 103152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_912
timestamp 1666464484
transform 1 0 103488 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_944
timestamp 1666464484
transform 1 0 107072 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_947
timestamp 1666464484
transform 1 0 107408 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_979
timestamp 1666464484
transform 1 0 110992 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_982
timestamp 1666464484
transform 1 0 111328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1014
timestamp 1666464484
transform 1 0 114912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1017
timestamp 1666464484
transform 1 0 115248 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1049
timestamp 1666464484
transform 1 0 118832 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1052
timestamp 1666464484
transform 1 0 119168 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1084
timestamp 1666464484
transform 1 0 122752 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1087
timestamp 1666464484
transform 1 0 123088 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1119
timestamp 1666464484
transform 1 0 126672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1122
timestamp 1666464484
transform 1 0 127008 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1154
timestamp 1666464484
transform 1 0 130592 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1157
timestamp 1666464484
transform 1 0 130928 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1189
timestamp 1666464484
transform 1 0 134512 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1192
timestamp 1666464484
transform 1 0 134848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1224
timestamp 1666464484
transform 1 0 138432 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1227
timestamp 1666464484
transform 1 0 138768 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1259
timestamp 1666464484
transform 1 0 142352 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_1262
timestamp 1666464484
transform 1 0 142688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1270
timestamp 1666464484
transform 1 0 143584 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1274
timestamp 1666464484
transform 1 0 144032 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1278
timestamp 1666464484
transform 1 0 144480 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1294
timestamp 1666464484
transform 1 0 146272 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1297
timestamp 1666464484
transform 1 0 146608 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1312
timestamp 1666464484
transform 1 0 148288 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1666464484
transform -1 0 148624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1666464484
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1666464484
transform -1 0 148624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1666464484
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1666464484
transform -1 0 148624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1666464484
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1666464484
transform -1 0 148624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1666464484
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1666464484
transform -1 0 148624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1666464484
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1666464484
transform -1 0 148624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1666464484
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1666464484
transform -1 0 148624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1666464484
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1666464484
transform -1 0 148624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1666464484
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1666464484
transform -1 0 148624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1666464484
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1666464484
transform -1 0 148624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1666464484
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1666464484
transform -1 0 148624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1666464484
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1666464484
transform -1 0 148624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1666464484
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1666464484
transform -1 0 148624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1666464484
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1666464484
transform -1 0 148624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1666464484
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1666464484
transform -1 0 148624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1666464484
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1666464484
transform -1 0 148624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1666464484
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1666464484
transform -1 0 148624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1666464484
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1666464484
transform -1 0 148624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1666464484
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1666464484
transform -1 0 148624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1666464484
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1666464484
transform -1 0 148624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1666464484
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1666464484
transform -1 0 148624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1666464484
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1666464484
transform -1 0 148624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1666464484
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1666464484
transform -1 0 148624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1666464484
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1666464484
transform -1 0 148624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1666464484
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1666464484
transform -1 0 148624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1666464484
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1666464484
transform -1 0 148624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1666464484
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1666464484
transform -1 0 148624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1666464484
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1666464484
transform -1 0 148624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1666464484
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1666464484
transform -1 0 148624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1666464484
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1666464484
transform -1 0 148624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1666464484
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1666464484
transform -1 0 148624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1666464484
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1666464484
transform -1 0 148624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1666464484
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1666464484
transform -1 0 148624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1666464484
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1666464484
transform -1 0 148624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1666464484
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1666464484
transform -1 0 148624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1666464484
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1666464484
transform -1 0 148624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1666464484
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1666464484
transform -1 0 148624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1666464484
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1666464484
transform -1 0 148624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1666464484
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1666464484
transform -1 0 148624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1666464484
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1666464484
transform -1 0 148624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1666464484
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1666464484
transform -1 0 148624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1666464484
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1666464484
transform -1 0 148624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1666464484
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1666464484
transform -1 0 148624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1666464484
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1666464484
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1666464484
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1666464484
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1666464484
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1666464484
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1666464484
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1666464484
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1666464484
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1666464484
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1666464484
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1666464484
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1666464484
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1666464484
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1666464484
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1666464484
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1666464484
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1666464484
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1666464484
transform 1 0 79744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1666464484
transform 1 0 83664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1666464484
transform 1 0 87584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1666464484
transform 1 0 91504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1666464484
transform 1 0 95424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1666464484
transform 1 0 99344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1666464484
transform 1 0 103264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1666464484
transform 1 0 107184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1666464484
transform 1 0 111104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1666464484
transform 1 0 115024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1666464484
transform 1 0 118944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1666464484
transform 1 0 122864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1666464484
transform 1 0 126784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1666464484
transform 1 0 130704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1666464484
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1666464484
transform 1 0 138544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1666464484
transform 1 0 142464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1666464484
transform 1 0 146384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1666464484
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1666464484
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1666464484
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1666464484
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1666464484
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1666464484
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1666464484
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1666464484
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1666464484
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1666464484
transform 1 0 80864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1666464484
transform 1 0 88816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1666464484
transform 1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1666464484
transform 1 0 104720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1666464484
transform 1 0 112672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1666464484
transform 1 0 120624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1666464484
transform 1 0 128576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1666464484
transform 1 0 136528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1666464484
transform 1 0 144480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1666464484
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1666464484
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1666464484
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1666464484
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1666464484
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1666464484
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1666464484
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1666464484
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1666464484
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1666464484
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1666464484
transform 1 0 84784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1666464484
transform 1 0 92736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1666464484
transform 1 0 100688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1666464484
transform 1 0 108640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1666464484
transform 1 0 116592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1666464484
transform 1 0 124544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1666464484
transform 1 0 132496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1666464484
transform 1 0 140448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1666464484
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1666464484
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1666464484
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1666464484
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1666464484
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1666464484
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1666464484
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1666464484
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1666464484
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1666464484
transform 1 0 80864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1666464484
transform 1 0 88816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1666464484
transform 1 0 96768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1666464484
transform 1 0 104720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1666464484
transform 1 0 112672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1666464484
transform 1 0 120624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1666464484
transform 1 0 128576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1666464484
transform 1 0 136528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1666464484
transform 1 0 144480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1666464484
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1666464484
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1666464484
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1666464484
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1666464484
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1666464484
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1666464484
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1666464484
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1666464484
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1666464484
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1666464484
transform 1 0 84784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1666464484
transform 1 0 92736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1666464484
transform 1 0 100688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1666464484
transform 1 0 108640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1666464484
transform 1 0 116592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1666464484
transform 1 0 124544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1666464484
transform 1 0 132496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1666464484
transform 1 0 140448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1666464484
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1666464484
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1666464484
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1666464484
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1666464484
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1666464484
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1666464484
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1666464484
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1666464484
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1666464484
transform 1 0 80864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1666464484
transform 1 0 88816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1666464484
transform 1 0 96768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1666464484
transform 1 0 104720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1666464484
transform 1 0 112672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1666464484
transform 1 0 120624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1666464484
transform 1 0 128576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1666464484
transform 1 0 136528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1666464484
transform 1 0 144480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1666464484
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1666464484
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1666464484
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1666464484
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1666464484
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1666464484
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1666464484
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1666464484
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1666464484
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1666464484
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1666464484
transform 1 0 84784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1666464484
transform 1 0 92736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1666464484
transform 1 0 100688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1666464484
transform 1 0 108640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1666464484
transform 1 0 116592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1666464484
transform 1 0 124544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1666464484
transform 1 0 132496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1666464484
transform 1 0 140448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1666464484
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1666464484
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1666464484
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1666464484
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1666464484
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1666464484
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1666464484
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1666464484
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1666464484
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1666464484
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1666464484
transform 1 0 88816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1666464484
transform 1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1666464484
transform 1 0 104720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1666464484
transform 1 0 112672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1666464484
transform 1 0 120624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1666464484
transform 1 0 128576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1666464484
transform 1 0 136528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1666464484
transform 1 0 144480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1666464484
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1666464484
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1666464484
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1666464484
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1666464484
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1666464484
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1666464484
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1666464484
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1666464484
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1666464484
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1666464484
transform 1 0 84784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1666464484
transform 1 0 92736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1666464484
transform 1 0 100688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1666464484
transform 1 0 108640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1666464484
transform 1 0 116592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1666464484
transform 1 0 124544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1666464484
transform 1 0 132496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1666464484
transform 1 0 140448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1666464484
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1666464484
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1666464484
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1666464484
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1666464484
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1666464484
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1666464484
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1666464484
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1666464484
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1666464484
transform 1 0 80864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1666464484
transform 1 0 88816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1666464484
transform 1 0 96768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1666464484
transform 1 0 104720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1666464484
transform 1 0 112672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1666464484
transform 1 0 120624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1666464484
transform 1 0 128576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1666464484
transform 1 0 136528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1666464484
transform 1 0 144480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1666464484
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1666464484
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1666464484
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1666464484
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1666464484
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1666464484
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1666464484
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1666464484
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1666464484
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1666464484
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1666464484
transform 1 0 84784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1666464484
transform 1 0 92736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1666464484
transform 1 0 100688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1666464484
transform 1 0 108640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1666464484
transform 1 0 116592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1666464484
transform 1 0 124544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1666464484
transform 1 0 132496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1666464484
transform 1 0 140448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1666464484
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1666464484
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1666464484
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1666464484
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1666464484
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1666464484
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1666464484
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1666464484
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1666464484
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1666464484
transform 1 0 80864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1666464484
transform 1 0 88816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1666464484
transform 1 0 96768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1666464484
transform 1 0 104720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1666464484
transform 1 0 112672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1666464484
transform 1 0 120624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1666464484
transform 1 0 128576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1666464484
transform 1 0 136528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1666464484
transform 1 0 144480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1666464484
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1666464484
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1666464484
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1666464484
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1666464484
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1666464484
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1666464484
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1666464484
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1666464484
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1666464484
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1666464484
transform 1 0 84784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1666464484
transform 1 0 92736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1666464484
transform 1 0 100688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1666464484
transform 1 0 108640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1666464484
transform 1 0 116592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1666464484
transform 1 0 124544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1666464484
transform 1 0 132496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1666464484
transform 1 0 140448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1666464484
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1666464484
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1666464484
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1666464484
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1666464484
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1666464484
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1666464484
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1666464484
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1666464484
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1666464484
transform 1 0 80864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1666464484
transform 1 0 88816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1666464484
transform 1 0 96768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1666464484
transform 1 0 104720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1666464484
transform 1 0 112672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1666464484
transform 1 0 120624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1666464484
transform 1 0 128576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1666464484
transform 1 0 136528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1666464484
transform 1 0 144480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1666464484
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1666464484
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1666464484
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1666464484
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1666464484
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1666464484
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1666464484
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1666464484
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1666464484
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1666464484
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1666464484
transform 1 0 84784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1666464484
transform 1 0 92736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1666464484
transform 1 0 100688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1666464484
transform 1 0 108640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1666464484
transform 1 0 116592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1666464484
transform 1 0 124544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1666464484
transform 1 0 132496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1666464484
transform 1 0 140448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1666464484
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1666464484
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1666464484
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1666464484
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1666464484
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1666464484
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1666464484
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1666464484
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1666464484
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1666464484
transform 1 0 80864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1666464484
transform 1 0 88816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1666464484
transform 1 0 96768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1666464484
transform 1 0 104720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1666464484
transform 1 0 112672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1666464484
transform 1 0 120624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1666464484
transform 1 0 128576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1666464484
transform 1 0 136528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1666464484
transform 1 0 144480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1666464484
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1666464484
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1666464484
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1666464484
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1666464484
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1666464484
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1666464484
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1666464484
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1666464484
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1666464484
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1666464484
transform 1 0 84784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1666464484
transform 1 0 92736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1666464484
transform 1 0 100688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1666464484
transform 1 0 108640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1666464484
transform 1 0 116592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1666464484
transform 1 0 124544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1666464484
transform 1 0 132496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1666464484
transform 1 0 140448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1666464484
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1666464484
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1666464484
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1666464484
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1666464484
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1666464484
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1666464484
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1666464484
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1666464484
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1666464484
transform 1 0 80864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1666464484
transform 1 0 88816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1666464484
transform 1 0 96768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1666464484
transform 1 0 104720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1666464484
transform 1 0 112672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1666464484
transform 1 0 120624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1666464484
transform 1 0 128576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1666464484
transform 1 0 136528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1666464484
transform 1 0 144480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1666464484
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1666464484
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1666464484
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1666464484
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1666464484
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1666464484
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1666464484
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1666464484
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1666464484
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1666464484
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1666464484
transform 1 0 84784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1666464484
transform 1 0 92736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1666464484
transform 1 0 100688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1666464484
transform 1 0 108640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1666464484
transform 1 0 116592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1666464484
transform 1 0 124544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1666464484
transform 1 0 132496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1666464484
transform 1 0 140448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1666464484
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1666464484
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1666464484
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1666464484
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1666464484
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1666464484
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1666464484
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1666464484
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1666464484
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1666464484
transform 1 0 80864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1666464484
transform 1 0 88816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1666464484
transform 1 0 96768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1666464484
transform 1 0 104720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1666464484
transform 1 0 112672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1666464484
transform 1 0 120624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1666464484
transform 1 0 128576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1666464484
transform 1 0 136528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1666464484
transform 1 0 144480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1666464484
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1666464484
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1666464484
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1666464484
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1666464484
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1666464484
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1666464484
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1666464484
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1666464484
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1666464484
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1666464484
transform 1 0 84784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1666464484
transform 1 0 92736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1666464484
transform 1 0 100688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1666464484
transform 1 0 108640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1666464484
transform 1 0 116592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1666464484
transform 1 0 124544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1666464484
transform 1 0 132496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1666464484
transform 1 0 140448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1666464484
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1666464484
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1666464484
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1666464484
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1666464484
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1666464484
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1666464484
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1666464484
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1666464484
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1666464484
transform 1 0 80864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1666464484
transform 1 0 88816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1666464484
transform 1 0 96768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1666464484
transform 1 0 104720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1666464484
transform 1 0 112672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1666464484
transform 1 0 120624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1666464484
transform 1 0 128576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1666464484
transform 1 0 136528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1666464484
transform 1 0 144480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1666464484
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1666464484
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1666464484
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1666464484
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1666464484
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1666464484
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1666464484
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1666464484
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1666464484
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1666464484
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1666464484
transform 1 0 84784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1666464484
transform 1 0 92736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1666464484
transform 1 0 100688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1666464484
transform 1 0 108640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1666464484
transform 1 0 116592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1666464484
transform 1 0 124544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1666464484
transform 1 0 132496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1666464484
transform 1 0 140448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1666464484
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1666464484
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1666464484
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1666464484
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1666464484
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1666464484
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1666464484
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1666464484
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1666464484
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1666464484
transform 1 0 80864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1666464484
transform 1 0 88816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1666464484
transform 1 0 96768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1666464484
transform 1 0 104720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1666464484
transform 1 0 112672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1666464484
transform 1 0 120624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1666464484
transform 1 0 128576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1666464484
transform 1 0 136528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1666464484
transform 1 0 144480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1666464484
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1666464484
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1666464484
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1666464484
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1666464484
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1666464484
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1666464484
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1666464484
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1666464484
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1666464484
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1666464484
transform 1 0 84784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1666464484
transform 1 0 92736 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1666464484
transform 1 0 100688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1666464484
transform 1 0 108640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1666464484
transform 1 0 116592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1666464484
transform 1 0 124544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1666464484
transform 1 0 132496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1666464484
transform 1 0 140448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1666464484
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1666464484
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1666464484
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1666464484
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1666464484
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1666464484
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1666464484
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1666464484
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1666464484
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1666464484
transform 1 0 80864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1666464484
transform 1 0 88816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1666464484
transform 1 0 96768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1666464484
transform 1 0 104720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1666464484
transform 1 0 112672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1666464484
transform 1 0 120624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1666464484
transform 1 0 128576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1666464484
transform 1 0 136528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1666464484
transform 1 0 144480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1666464484
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1666464484
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1666464484
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1666464484
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1666464484
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1666464484
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1666464484
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1666464484
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1666464484
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1666464484
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1666464484
transform 1 0 84784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1666464484
transform 1 0 92736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1666464484
transform 1 0 100688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1666464484
transform 1 0 108640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1666464484
transform 1 0 116592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1666464484
transform 1 0 124544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1666464484
transform 1 0 132496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1666464484
transform 1 0 140448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1666464484
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1666464484
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1666464484
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1666464484
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1666464484
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1666464484
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1666464484
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1666464484
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1666464484
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1666464484
transform 1 0 80864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1666464484
transform 1 0 88816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1666464484
transform 1 0 96768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1666464484
transform 1 0 104720 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1666464484
transform 1 0 112672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1666464484
transform 1 0 120624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1666464484
transform 1 0 128576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1666464484
transform 1 0 136528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1666464484
transform 1 0 144480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1666464484
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1666464484
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1666464484
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1666464484
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1666464484
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1666464484
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1666464484
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1666464484
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1666464484
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1666464484
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1666464484
transform 1 0 84784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1666464484
transform 1 0 92736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1666464484
transform 1 0 100688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1666464484
transform 1 0 108640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1666464484
transform 1 0 116592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1666464484
transform 1 0 124544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1666464484
transform 1 0 132496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1666464484
transform 1 0 140448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1666464484
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1666464484
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1666464484
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1666464484
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1666464484
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1666464484
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1666464484
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1666464484
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1666464484
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1666464484
transform 1 0 80864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1666464484
transform 1 0 88816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1666464484
transform 1 0 96768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1666464484
transform 1 0 104720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1666464484
transform 1 0 112672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1666464484
transform 1 0 120624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1666464484
transform 1 0 128576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1666464484
transform 1 0 136528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1666464484
transform 1 0 144480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1666464484
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1666464484
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1666464484
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1666464484
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1666464484
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1666464484
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1666464484
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1666464484
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1666464484
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1666464484
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1666464484
transform 1 0 84784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1666464484
transform 1 0 92736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1666464484
transform 1 0 100688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1666464484
transform 1 0 108640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1666464484
transform 1 0 116592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1666464484
transform 1 0 124544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1666464484
transform 1 0 132496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1666464484
transform 1 0 140448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1666464484
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1666464484
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1666464484
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1666464484
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1666464484
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1666464484
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1666464484
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1666464484
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1666464484
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1666464484
transform 1 0 80864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1666464484
transform 1 0 88816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1666464484
transform 1 0 96768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1666464484
transform 1 0 104720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1666464484
transform 1 0 112672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1666464484
transform 1 0 120624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1666464484
transform 1 0 128576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1666464484
transform 1 0 136528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1666464484
transform 1 0 144480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1666464484
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1666464484
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1666464484
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1666464484
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1666464484
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1666464484
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1666464484
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1666464484
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1666464484
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1666464484
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1666464484
transform 1 0 84784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1666464484
transform 1 0 92736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1666464484
transform 1 0 100688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1666464484
transform 1 0 108640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1666464484
transform 1 0 116592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1666464484
transform 1 0 124544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1666464484
transform 1 0 132496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1666464484
transform 1 0 140448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1666464484
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1666464484
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1666464484
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1666464484
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1666464484
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1666464484
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1666464484
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1666464484
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1666464484
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1666464484
transform 1 0 80864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1666464484
transform 1 0 88816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1666464484
transform 1 0 96768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1666464484
transform 1 0 104720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1666464484
transform 1 0 112672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1666464484
transform 1 0 120624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1666464484
transform 1 0 128576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1666464484
transform 1 0 136528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1666464484
transform 1 0 144480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1666464484
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1666464484
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1666464484
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1666464484
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1666464484
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1666464484
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1666464484
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1666464484
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1666464484
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1666464484
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1666464484
transform 1 0 84784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1666464484
transform 1 0 92736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1666464484
transform 1 0 100688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1666464484
transform 1 0 108640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1666464484
transform 1 0 116592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1666464484
transform 1 0 124544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1666464484
transform 1 0 132496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1666464484
transform 1 0 140448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1666464484
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1666464484
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1666464484
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1666464484
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1666464484
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1666464484
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1666464484
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1666464484
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1666464484
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1666464484
transform 1 0 80864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1666464484
transform 1 0 88816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1666464484
transform 1 0 96768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1666464484
transform 1 0 104720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1666464484
transform 1 0 112672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1666464484
transform 1 0 120624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1666464484
transform 1 0 128576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1666464484
transform 1 0 136528 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1666464484
transform 1 0 144480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1666464484
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1666464484
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1666464484
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1666464484
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1666464484
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1666464484
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1666464484
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1666464484
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1666464484
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1666464484
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1666464484
transform 1 0 84784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1666464484
transform 1 0 92736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1666464484
transform 1 0 100688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1666464484
transform 1 0 108640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1666464484
transform 1 0 116592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1666464484
transform 1 0 124544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1666464484
transform 1 0 132496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1666464484
transform 1 0 140448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1666464484
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1666464484
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1666464484
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1666464484
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1666464484
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1666464484
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1666464484
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1666464484
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1666464484
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1666464484
transform 1 0 80864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1666464484
transform 1 0 88816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1666464484
transform 1 0 96768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1666464484
transform 1 0 104720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1666464484
transform 1 0 112672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1666464484
transform 1 0 120624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1666464484
transform 1 0 128576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1666464484
transform 1 0 136528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1666464484
transform 1 0 144480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1666464484
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1666464484
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1666464484
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1666464484
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1666464484
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1666464484
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1666464484
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1666464484
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1666464484
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1666464484
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1666464484
transform 1 0 84784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1666464484
transform 1 0 92736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1666464484
transform 1 0 100688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1666464484
transform 1 0 108640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1666464484
transform 1 0 116592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1666464484
transform 1 0 124544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1666464484
transform 1 0 132496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1666464484
transform 1 0 140448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1666464484
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1666464484
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1666464484
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1666464484
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1666464484
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1666464484
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1666464484
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1666464484
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1666464484
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1666464484
transform 1 0 80864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1666464484
transform 1 0 88816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1666464484
transform 1 0 96768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1666464484
transform 1 0 104720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1666464484
transform 1 0 112672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1666464484
transform 1 0 120624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1666464484
transform 1 0 128576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1666464484
transform 1 0 136528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1666464484
transform 1 0 144480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1666464484
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1666464484
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1666464484
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1666464484
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1666464484
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1666464484
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1666464484
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1666464484
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1666464484
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1666464484
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1666464484
transform 1 0 84784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1666464484
transform 1 0 92736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1666464484
transform 1 0 100688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1666464484
transform 1 0 108640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1666464484
transform 1 0 116592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1666464484
transform 1 0 124544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1666464484
transform 1 0 132496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1666464484
transform 1 0 140448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1666464484
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1666464484
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1666464484
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1666464484
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1666464484
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1666464484
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1666464484
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1666464484
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1666464484
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1666464484
transform 1 0 80864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1666464484
transform 1 0 88816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1666464484
transform 1 0 96768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1666464484
transform 1 0 104720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1666464484
transform 1 0 112672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1666464484
transform 1 0 120624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1666464484
transform 1 0 128576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1666464484
transform 1 0 136528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1666464484
transform 1 0 144480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1666464484
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1666464484
transform 1 0 9184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1666464484
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1666464484
transform 1 0 17024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1666464484
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1666464484
transform 1 0 24864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1666464484
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1666464484
transform 1 0 32704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1666464484
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1666464484
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1666464484
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1666464484
transform 1 0 48384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1666464484
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1666464484
transform 1 0 56224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1666464484
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1666464484
transform 1 0 64064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1666464484
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1666464484
transform 1 0 71904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1666464484
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1666464484
transform 1 0 79744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1666464484
transform 1 0 83664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1666464484
transform 1 0 87584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1666464484
transform 1 0 91504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1666464484
transform 1 0 95424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1666464484
transform 1 0 99344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1666464484
transform 1 0 103264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1666464484
transform 1 0 107184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1666464484
transform 1 0 111104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1666464484
transform 1 0 115024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1666464484
transform 1 0 118944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1666464484
transform 1 0 122864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1666464484
transform 1 0 126784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1666464484
transform 1 0 130704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1666464484
transform 1 0 134624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1666464484
transform 1 0 138544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1666464484
transform 1 0 142464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1666464484
transform 1 0 146384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _042_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 135072 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _043_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 129808 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _044_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 123536 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _045_
timestamp 1666464484
transform 1 0 123424 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _046_
timestamp 1666464484
transform -1 0 124880 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _047_
timestamp 1666464484
transform 1 0 124880 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _048_
timestamp 1666464484
transform -1 0 125664 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _049_
timestamp 1666464484
transform 1 0 125776 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _050_
timestamp 1666464484
transform -1 0 127568 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _051_
timestamp 1666464484
transform 1 0 127792 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _052_
timestamp 1666464484
transform -1 0 131824 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _053_
timestamp 1666464484
transform -1 0 130368 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _054_
timestamp 1666464484
transform 1 0 130032 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _055_
timestamp 1666464484
transform -1 0 131040 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _056_
timestamp 1666464484
transform 1 0 130928 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _057_
timestamp 1666464484
transform -1 0 132720 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _058_
timestamp 1666464484
transform 1 0 132832 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _059_
timestamp 1666464484
transform -1 0 133168 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _060_
timestamp 1666464484
transform 1 0 133728 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _061_
timestamp 1666464484
transform 1 0 135520 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _062_
timestamp 1666464484
transform -1 0 136976 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _063_
timestamp 1666464484
transform 1 0 137312 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _064_
timestamp 1666464484
transform -1 0 138544 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _065_
timestamp 1666464484
transform 1 0 138992 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _066_
timestamp 1666464484
transform -1 0 140560 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _067_
timestamp 1666464484
transform 1 0 140336 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _068_
timestamp 1666464484
transform -1 0 140560 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _069_
timestamp 1666464484
transform 1 0 141232 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _070_
timestamp 1666464484
transform -1 0 134288 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _071_
timestamp 1666464484
transform -1 0 144480 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _072_
timestamp 1666464484
transform 1 0 143584 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _073_
timestamp 1666464484
transform -1 0 142464 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _074_
timestamp 1666464484
transform 1 0 142128 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _075_
timestamp 1666464484
transform -1 0 142464 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _076_
timestamp 1666464484
transform 1 0 142688 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _077_
timestamp 1666464484
transform 1 0 113008 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _078_
timestamp 1666464484
transform 1 0 113008 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _079_
timestamp 1666464484
transform -1 0 127568 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _080_
timestamp 1666464484
transform -1 0 102816 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _081_
timestamp 1666464484
transform -1 0 99792 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _082_
timestamp 1666464484
transform 1 0 99120 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _083_
timestamp 1666464484
transform -1 0 99232 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _084_
timestamp 1666464484
transform 1 0 99344 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _085_
timestamp 1666464484
transform -1 0 101360 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _086_
timestamp 1666464484
transform 1 0 100240 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _087_
timestamp 1666464484
transform -1 0 101696 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _088_
timestamp 1666464484
transform 1 0 101360 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _089_
timestamp 1666464484
transform -1 0 104160 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _090_
timestamp 1666464484
transform -1 0 103600 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _091_
timestamp 1666464484
transform 1 0 103824 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _092_
timestamp 1666464484
transform -1 0 105280 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _093_
timestamp 1666464484
transform 1 0 105392 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _094_
timestamp 1666464484
transform -1 0 105168 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _095_
timestamp 1666464484
transform 1 0 105056 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _096_
timestamp 1666464484
transform -1 0 106736 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _097_
timestamp 1666464484
transform 1 0 106288 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _098_
timestamp 1666464484
transform -1 0 111440 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _099_
timestamp 1666464484
transform -1 0 110880 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _100_
timestamp 1666464484
transform 1 0 109872 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _101_
timestamp 1666464484
transform -1 0 113120 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _102_
timestamp 1666464484
transform 1 0 113568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _103_
timestamp 1666464484
transform -1 0 111888 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _104_
timestamp 1666464484
transform 1 0 111664 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _105_
timestamp 1666464484
transform -1 0 112448 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _106_
timestamp 1666464484
transform 1 0 112672 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _107_
timestamp 1666464484
transform -1 0 117824 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _108_
timestamp 1666464484
transform 1 0 115360 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _109_
timestamp 1666464484
transform 1 0 115808 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _110_
timestamp 1666464484
transform -1 0 117376 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _111_
timestamp 1666464484
transform 1 0 118048 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _112_
timestamp 1666464484
transform -1 0 119280 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _113_
timestamp 1666464484
transform 1 0 118944 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _114_
timestamp 1666464484
transform -1 0 120960 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _115_
timestamp 1666464484
transform 1 0 119840 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _116_
timestamp 1666464484
transform -1 0 75712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _117_
timestamp 1666464484
transform -1 0 78400 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _118_
timestamp 1666464484
transform -1 0 80192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _119_
timestamp 1666464484
transform -1 0 81088 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _120_
timestamp 1666464484
transform -1 0 83440 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _121_
timestamp 1666464484
transform -1 0 84448 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _122_
timestamp 1666464484
transform -1 0 86128 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _123_
timestamp 1666464484
transform -1 0 87808 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _124_
timestamp 1666464484
transform -1 0 89488 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _125_
timestamp 1666464484
transform 1 0 76832 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_
timestamp 1666464484
transform 1 0 78624 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _127_
timestamp 1666464484
transform 1 0 81200 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _128_
timestamp 1666464484
transform 1 0 81872 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _129_
timestamp 1666464484
transform 1 0 84336 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _130_
timestamp 1666464484
transform -1 0 86688 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1666464484
transform 1 0 87696 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _132_
timestamp 1666464484
transform 1 0 89152 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _133_
timestamp 1666464484
transform 1 0 90272 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _134_
timestamp 1666464484
transform -1 0 73920 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _135_
timestamp 1666464484
transform 1 0 75152 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1666464484
transform -1 0 148288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1666464484
transform -1 0 147392 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1666464484
transform -1 0 148288 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1666464484
transform -1 0 148288 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1666464484
transform -1 0 148288 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1666464484
transform -1 0 148288 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1666464484
transform -1 0 148288 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1666464484
transform -1 0 148288 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1666464484
transform -1 0 148288 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1666464484
transform -1 0 148288 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1666464484
transform -1 0 147392 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1666464484
transform 1 0 22064 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1666464484
transform 1 0 38864 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1666464484
transform 1 0 40880 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1666464484
transform 1 0 42224 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1666464484
transform 1 0 43680 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1666464484
transform 1 0 45584 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1666464484
transform 1 0 47264 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1666464484
transform 1 0 48944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1666464484
transform 1 0 50624 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1666464484
transform 1 0 52640 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1666464484
transform 1 0 53984 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1666464484
transform 1 0 23744 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1666464484
transform 1 0 55440 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1666464484
transform 1 0 57344 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1666464484
transform 1 0 59024 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1666464484
transform 1 0 60704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1666464484
transform 1 0 62384 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1666464484
transform 1 0 64400 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1666464484
transform 1 0 65744 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1666464484
transform 1 0 67200 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1666464484
transform 1 0 69104 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1666464484
transform 1 0 70784 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1666464484
transform 1 0 25424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1666464484
transform 1 0 72352 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1666464484
transform 1 0 74144 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1666464484
transform 1 0 27104 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1666464484
transform 1 0 29120 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1666464484
transform 1 0 30464 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1666464484
transform 1 0 31920 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1666464484
transform 1 0 33824 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1666464484
transform 1 0 35504 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1666464484
transform 1 0 37184 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1666464484
transform 1 0 93632 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1666464484
transform 1 0 109312 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1666464484
transform -1 0 114016 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1666464484
transform -1 0 114912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1666464484
transform 1 0 114464 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1666464484
transform -1 0 117936 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1666464484
transform 1 0 118160 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1666464484
transform 1 0 119504 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1666464484
transform 1 0 121184 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1666464484
transform 1 0 122080 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1666464484
transform -1 0 125776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1666464484
transform 1 0 94528 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1666464484
transform -1 0 127792 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1666464484
transform 1 0 127792 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1666464484
transform 1 0 129584 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1666464484
transform -1 0 133616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1666464484
transform -1 0 134512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1666464484
transform 1 0 134624 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1666464484
transform 1 0 137200 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input63
timestamp 1666464484
transform -1 0 141456 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1666464484
transform -1 0 142352 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input65
timestamp 1666464484
transform 1 0 142688 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input66
timestamp 1666464484
transform 1 0 95984 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input67
timestamp 1666464484
transform -1 0 144256 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input68
timestamp 1666464484
transform -1 0 145376 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input69
timestamp 1666464484
transform 1 0 97216 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input70
timestamp 1666464484
transform 1 0 99344 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input71
timestamp 1666464484
transform 1 0 101584 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input72
timestamp 1666464484
transform 1 0 102480 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input73
timestamp 1666464484
transform -1 0 106176 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1666464484
transform -1 0 107072 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1666464484
transform 1 0 107744 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output76 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 8512 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output77
timestamp 1666464484
transform -1 0 9072 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output78
timestamp 1666464484
transform -1 0 11200 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output79
timestamp 1666464484
transform -1 0 12992 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output80
timestamp 1666464484
transform -1 0 15120 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output81
timestamp 1666464484
transform -1 0 16912 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output82
timestamp 1666464484
transform -1 0 19152 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output83
timestamp 1666464484
transform -1 0 20272 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output84
timestamp 1666464484
transform -1 0 22848 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output85
timestamp 1666464484
transform 1 0 77952 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output86
timestamp 1666464484
transform 1 0 80080 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output87
timestamp 1666464484
transform 1 0 81872 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output88
timestamp 1666464484
transform 1 0 82544 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output89
timestamp 1666464484
transform -1 0 85792 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output90
timestamp 1666464484
transform 1 0 85904 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output91
timestamp 1666464484
transform 1 0 87920 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output92
timestamp 1666464484
transform 1 0 89712 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output93
timestamp 1666464484
transform 1 0 91840 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output94
timestamp 1666464484
transform -1 0 7168 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output95
timestamp 1666464484
transform 1 0 76160 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output96
timestamp 1666464484
transform 1 0 146720 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output97
timestamp 1666464484
transform 1 0 146720 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output98
timestamp 1666464484
transform 1 0 146720 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output99
timestamp 1666464484
transform 1 0 146720 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output100
timestamp 1666464484
transform 1 0 146720 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output101
timestamp 1666464484
transform 1 0 146720 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output102
timestamp 1666464484
transform 1 0 146720 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output103
timestamp 1666464484
transform 1 0 146720 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output104
timestamp 1666464484
transform 1 0 146720 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output105
timestamp 1666464484
transform 1 0 146720 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output106
timestamp 1666464484
transform 1 0 146720 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output107
timestamp 1666464484
transform 1 0 146720 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output108
timestamp 1666464484
transform 1 0 146720 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output109
timestamp 1666464484
transform 1 0 146720 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output110
timestamp 1666464484
transform 1 0 146720 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output111
timestamp 1666464484
transform 1 0 146720 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output112
timestamp 1666464484
transform 1 0 146720 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output113
timestamp 1666464484
transform 1 0 146720 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output114
timestamp 1666464484
transform 1 0 146720 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output115
timestamp 1666464484
transform 1 0 146720 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output116
timestamp 1666464484
transform 1 0 146720 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output117
timestamp 1666464484
transform 1 0 144704 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output118
timestamp 1666464484
transform 1 0 146720 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output119
timestamp 1666464484
transform 1 0 144928 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output120
timestamp 1666464484
transform 1 0 144928 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output121
timestamp 1666464484
transform 1 0 146720 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output122
timestamp 1666464484
transform 1 0 146720 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output123
timestamp 1666464484
transform 1 0 146720 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output124
timestamp 1666464484
transform 1 0 146720 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output125
timestamp 1666464484
transform 1 0 146720 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output126
timestamp 1666464484
transform 1 0 146720 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output127
timestamp 1666464484
transform 1 0 146720 0 1 18816
box -86 -86 1654 870
<< labels >>
flabel metal3 s 149200 2016 150000 2128 0 FreeSans 448 0 0 0 addr[0]
port 0 nsew signal input
flabel metal3 s 149200 2912 150000 3024 0 FreeSans 448 0 0 0 addr[1]
port 1 nsew signal input
flabel metal3 s 149200 3808 150000 3920 0 FreeSans 448 0 0 0 addr[2]
port 2 nsew signal input
flabel metal3 s 149200 4704 150000 4816 0 FreeSans 448 0 0 0 addr[3]
port 3 nsew signal input
flabel metal3 s 149200 5600 150000 5712 0 FreeSans 448 0 0 0 addr[4]
port 4 nsew signal input
flabel metal3 s 149200 6496 150000 6608 0 FreeSans 448 0 0 0 addr[5]
port 5 nsew signal input
flabel metal3 s 149200 7392 150000 7504 0 FreeSans 448 0 0 0 addr[6]
port 6 nsew signal input
flabel metal3 s 149200 8288 150000 8400 0 FreeSans 448 0 0 0 addr[7]
port 7 nsew signal input
flabel metal3 s 149200 9184 150000 9296 0 FreeSans 448 0 0 0 addr[8]
port 8 nsew signal input
flabel metal3 s 149200 10080 150000 10192 0 FreeSans 448 0 0 0 addr[9]
port 9 nsew signal input
flabel metal2 s 6832 0 6944 800 0 FreeSans 448 90 0 0 addr_mem0[0]
port 10 nsew signal tristate
flabel metal2 s 8512 0 8624 800 0 FreeSans 448 90 0 0 addr_mem0[1]
port 11 nsew signal tristate
flabel metal2 s 10192 0 10304 800 0 FreeSans 448 90 0 0 addr_mem0[2]
port 12 nsew signal tristate
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 addr_mem0[3]
port 13 nsew signal tristate
flabel metal2 s 13552 0 13664 800 0 FreeSans 448 90 0 0 addr_mem0[4]
port 14 nsew signal tristate
flabel metal2 s 15232 0 15344 800 0 FreeSans 448 90 0 0 addr_mem0[5]
port 15 nsew signal tristate
flabel metal2 s 16912 0 17024 800 0 FreeSans 448 90 0 0 addr_mem0[6]
port 16 nsew signal tristate
flabel metal2 s 18592 0 18704 800 0 FreeSans 448 90 0 0 addr_mem0[7]
port 17 nsew signal tristate
flabel metal2 s 20272 0 20384 800 0 FreeSans 448 90 0 0 addr_mem0[8]
port 18 nsew signal tristate
flabel metal2 s 77392 0 77504 800 0 FreeSans 448 90 0 0 addr_mem1[0]
port 19 nsew signal tristate
flabel metal2 s 79072 0 79184 800 0 FreeSans 448 90 0 0 addr_mem1[1]
port 20 nsew signal tristate
flabel metal2 s 80752 0 80864 800 0 FreeSans 448 90 0 0 addr_mem1[2]
port 21 nsew signal tristate
flabel metal2 s 82432 0 82544 800 0 FreeSans 448 90 0 0 addr_mem1[3]
port 22 nsew signal tristate
flabel metal2 s 84112 0 84224 800 0 FreeSans 448 90 0 0 addr_mem1[4]
port 23 nsew signal tristate
flabel metal2 s 85792 0 85904 800 0 FreeSans 448 90 0 0 addr_mem1[5]
port 24 nsew signal tristate
flabel metal2 s 87472 0 87584 800 0 FreeSans 448 90 0 0 addr_mem1[6]
port 25 nsew signal tristate
flabel metal2 s 89152 0 89264 800 0 FreeSans 448 90 0 0 addr_mem1[7]
port 26 nsew signal tristate
flabel metal2 s 90832 0 90944 800 0 FreeSans 448 90 0 0 addr_mem1[8]
port 27 nsew signal tristate
flabel metal3 s 149200 1120 150000 1232 0 FreeSans 448 0 0 0 csb
port 28 nsew signal input
flabel metal2 s 5152 0 5264 800 0 FreeSans 448 90 0 0 csb_mem0
port 29 nsew signal tristate
flabel metal2 s 75712 0 75824 800 0 FreeSans 448 90 0 0 csb_mem1
port 30 nsew signal tristate
flabel metal3 s 149200 10976 150000 11088 0 FreeSans 448 0 0 0 dout[0]
port 31 nsew signal tristate
flabel metal3 s 149200 19936 150000 20048 0 FreeSans 448 0 0 0 dout[10]
port 32 nsew signal tristate
flabel metal3 s 149200 20832 150000 20944 0 FreeSans 448 0 0 0 dout[11]
port 33 nsew signal tristate
flabel metal3 s 149200 21728 150000 21840 0 FreeSans 448 0 0 0 dout[12]
port 34 nsew signal tristate
flabel metal3 s 149200 22624 150000 22736 0 FreeSans 448 0 0 0 dout[13]
port 35 nsew signal tristate
flabel metal3 s 149200 23520 150000 23632 0 FreeSans 448 0 0 0 dout[14]
port 36 nsew signal tristate
flabel metal3 s 149200 24416 150000 24528 0 FreeSans 448 0 0 0 dout[15]
port 37 nsew signal tristate
flabel metal3 s 149200 25312 150000 25424 0 FreeSans 448 0 0 0 dout[16]
port 38 nsew signal tristate
flabel metal3 s 149200 26208 150000 26320 0 FreeSans 448 0 0 0 dout[17]
port 39 nsew signal tristate
flabel metal3 s 149200 27104 150000 27216 0 FreeSans 448 0 0 0 dout[18]
port 40 nsew signal tristate
flabel metal3 s 149200 28000 150000 28112 0 FreeSans 448 0 0 0 dout[19]
port 41 nsew signal tristate
flabel metal3 s 149200 11872 150000 11984 0 FreeSans 448 0 0 0 dout[1]
port 42 nsew signal tristate
flabel metal3 s 149200 28896 150000 29008 0 FreeSans 448 0 0 0 dout[20]
port 43 nsew signal tristate
flabel metal3 s 149200 29792 150000 29904 0 FreeSans 448 0 0 0 dout[21]
port 44 nsew signal tristate
flabel metal3 s 149200 30688 150000 30800 0 FreeSans 448 0 0 0 dout[22]
port 45 nsew signal tristate
flabel metal3 s 149200 31584 150000 31696 0 FreeSans 448 0 0 0 dout[23]
port 46 nsew signal tristate
flabel metal3 s 149200 32480 150000 32592 0 FreeSans 448 0 0 0 dout[24]
port 47 nsew signal tristate
flabel metal3 s 149200 33376 150000 33488 0 FreeSans 448 0 0 0 dout[25]
port 48 nsew signal tristate
flabel metal3 s 149200 34272 150000 34384 0 FreeSans 448 0 0 0 dout[26]
port 49 nsew signal tristate
flabel metal3 s 149200 35168 150000 35280 0 FreeSans 448 0 0 0 dout[27]
port 50 nsew signal tristate
flabel metal3 s 149200 36064 150000 36176 0 FreeSans 448 0 0 0 dout[28]
port 51 nsew signal tristate
flabel metal3 s 149200 36960 150000 37072 0 FreeSans 448 0 0 0 dout[29]
port 52 nsew signal tristate
flabel metal3 s 149200 12768 150000 12880 0 FreeSans 448 0 0 0 dout[2]
port 53 nsew signal tristate
flabel metal3 s 149200 37856 150000 37968 0 FreeSans 448 0 0 0 dout[30]
port 54 nsew signal tristate
flabel metal3 s 149200 38752 150000 38864 0 FreeSans 448 0 0 0 dout[31]
port 55 nsew signal tristate
flabel metal3 s 149200 13664 150000 13776 0 FreeSans 448 0 0 0 dout[3]
port 56 nsew signal tristate
flabel metal3 s 149200 14560 150000 14672 0 FreeSans 448 0 0 0 dout[4]
port 57 nsew signal tristate
flabel metal3 s 149200 15456 150000 15568 0 FreeSans 448 0 0 0 dout[5]
port 58 nsew signal tristate
flabel metal3 s 149200 16352 150000 16464 0 FreeSans 448 0 0 0 dout[6]
port 59 nsew signal tristate
flabel metal3 s 149200 17248 150000 17360 0 FreeSans 448 0 0 0 dout[7]
port 60 nsew signal tristate
flabel metal3 s 149200 18144 150000 18256 0 FreeSans 448 0 0 0 dout[8]
port 61 nsew signal tristate
flabel metal3 s 149200 19040 150000 19152 0 FreeSans 448 0 0 0 dout[9]
port 62 nsew signal tristate
flabel metal2 s 21952 0 22064 800 0 FreeSans 448 90 0 0 dout_mem0[0]
port 63 nsew signal input
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 dout_mem0[10]
port 64 nsew signal input
flabel metal2 s 40432 0 40544 800 0 FreeSans 448 90 0 0 dout_mem0[11]
port 65 nsew signal input
flabel metal2 s 42112 0 42224 800 0 FreeSans 448 90 0 0 dout_mem0[12]
port 66 nsew signal input
flabel metal2 s 43792 0 43904 800 0 FreeSans 448 90 0 0 dout_mem0[13]
port 67 nsew signal input
flabel metal2 s 45472 0 45584 800 0 FreeSans 448 90 0 0 dout_mem0[14]
port 68 nsew signal input
flabel metal2 s 47152 0 47264 800 0 FreeSans 448 90 0 0 dout_mem0[15]
port 69 nsew signal input
flabel metal2 s 48832 0 48944 800 0 FreeSans 448 90 0 0 dout_mem0[16]
port 70 nsew signal input
flabel metal2 s 50512 0 50624 800 0 FreeSans 448 90 0 0 dout_mem0[17]
port 71 nsew signal input
flabel metal2 s 52192 0 52304 800 0 FreeSans 448 90 0 0 dout_mem0[18]
port 72 nsew signal input
flabel metal2 s 53872 0 53984 800 0 FreeSans 448 90 0 0 dout_mem0[19]
port 73 nsew signal input
flabel metal2 s 23632 0 23744 800 0 FreeSans 448 90 0 0 dout_mem0[1]
port 74 nsew signal input
flabel metal2 s 55552 0 55664 800 0 FreeSans 448 90 0 0 dout_mem0[20]
port 75 nsew signal input
flabel metal2 s 57232 0 57344 800 0 FreeSans 448 90 0 0 dout_mem0[21]
port 76 nsew signal input
flabel metal2 s 58912 0 59024 800 0 FreeSans 448 90 0 0 dout_mem0[22]
port 77 nsew signal input
flabel metal2 s 60592 0 60704 800 0 FreeSans 448 90 0 0 dout_mem0[23]
port 78 nsew signal input
flabel metal2 s 62272 0 62384 800 0 FreeSans 448 90 0 0 dout_mem0[24]
port 79 nsew signal input
flabel metal2 s 63952 0 64064 800 0 FreeSans 448 90 0 0 dout_mem0[25]
port 80 nsew signal input
flabel metal2 s 65632 0 65744 800 0 FreeSans 448 90 0 0 dout_mem0[26]
port 81 nsew signal input
flabel metal2 s 67312 0 67424 800 0 FreeSans 448 90 0 0 dout_mem0[27]
port 82 nsew signal input
flabel metal2 s 68992 0 69104 800 0 FreeSans 448 90 0 0 dout_mem0[28]
port 83 nsew signal input
flabel metal2 s 70672 0 70784 800 0 FreeSans 448 90 0 0 dout_mem0[29]
port 84 nsew signal input
flabel metal2 s 25312 0 25424 800 0 FreeSans 448 90 0 0 dout_mem0[2]
port 85 nsew signal input
flabel metal2 s 72352 0 72464 800 0 FreeSans 448 90 0 0 dout_mem0[30]
port 86 nsew signal input
flabel metal2 s 74032 0 74144 800 0 FreeSans 448 90 0 0 dout_mem0[31]
port 87 nsew signal input
flabel metal2 s 26992 0 27104 800 0 FreeSans 448 90 0 0 dout_mem0[3]
port 88 nsew signal input
flabel metal2 s 28672 0 28784 800 0 FreeSans 448 90 0 0 dout_mem0[4]
port 89 nsew signal input
flabel metal2 s 30352 0 30464 800 0 FreeSans 448 90 0 0 dout_mem0[5]
port 90 nsew signal input
flabel metal2 s 32032 0 32144 800 0 FreeSans 448 90 0 0 dout_mem0[6]
port 91 nsew signal input
flabel metal2 s 33712 0 33824 800 0 FreeSans 448 90 0 0 dout_mem0[7]
port 92 nsew signal input
flabel metal2 s 35392 0 35504 800 0 FreeSans 448 90 0 0 dout_mem0[8]
port 93 nsew signal input
flabel metal2 s 37072 0 37184 800 0 FreeSans 448 90 0 0 dout_mem0[9]
port 94 nsew signal input
flabel metal2 s 92512 0 92624 800 0 FreeSans 448 90 0 0 dout_mem1[0]
port 95 nsew signal input
flabel metal2 s 109312 0 109424 800 0 FreeSans 448 90 0 0 dout_mem1[10]
port 96 nsew signal input
flabel metal2 s 110992 0 111104 800 0 FreeSans 448 90 0 0 dout_mem1[11]
port 97 nsew signal input
flabel metal2 s 112672 0 112784 800 0 FreeSans 448 90 0 0 dout_mem1[12]
port 98 nsew signal input
flabel metal2 s 114352 0 114464 800 0 FreeSans 448 90 0 0 dout_mem1[13]
port 99 nsew signal input
flabel metal2 s 116032 0 116144 800 0 FreeSans 448 90 0 0 dout_mem1[14]
port 100 nsew signal input
flabel metal2 s 117712 0 117824 800 0 FreeSans 448 90 0 0 dout_mem1[15]
port 101 nsew signal input
flabel metal2 s 119392 0 119504 800 0 FreeSans 448 90 0 0 dout_mem1[16]
port 102 nsew signal input
flabel metal2 s 121072 0 121184 800 0 FreeSans 448 90 0 0 dout_mem1[17]
port 103 nsew signal input
flabel metal2 s 122752 0 122864 800 0 FreeSans 448 90 0 0 dout_mem1[18]
port 104 nsew signal input
flabel metal2 s 124432 0 124544 800 0 FreeSans 448 90 0 0 dout_mem1[19]
port 105 nsew signal input
flabel metal2 s 94192 0 94304 800 0 FreeSans 448 90 0 0 dout_mem1[1]
port 106 nsew signal input
flabel metal2 s 126112 0 126224 800 0 FreeSans 448 90 0 0 dout_mem1[20]
port 107 nsew signal input
flabel metal2 s 127792 0 127904 800 0 FreeSans 448 90 0 0 dout_mem1[21]
port 108 nsew signal input
flabel metal2 s 129472 0 129584 800 0 FreeSans 448 90 0 0 dout_mem1[22]
port 109 nsew signal input
flabel metal2 s 131152 0 131264 800 0 FreeSans 448 90 0 0 dout_mem1[23]
port 110 nsew signal input
flabel metal2 s 132832 0 132944 800 0 FreeSans 448 90 0 0 dout_mem1[24]
port 111 nsew signal input
flabel metal2 s 134512 0 134624 800 0 FreeSans 448 90 0 0 dout_mem1[25]
port 112 nsew signal input
flabel metal2 s 136192 0 136304 800 0 FreeSans 448 90 0 0 dout_mem1[26]
port 113 nsew signal input
flabel metal2 s 137872 0 137984 800 0 FreeSans 448 90 0 0 dout_mem1[27]
port 114 nsew signal input
flabel metal2 s 139552 0 139664 800 0 FreeSans 448 90 0 0 dout_mem1[28]
port 115 nsew signal input
flabel metal2 s 141232 0 141344 800 0 FreeSans 448 90 0 0 dout_mem1[29]
port 116 nsew signal input
flabel metal2 s 95872 0 95984 800 0 FreeSans 448 90 0 0 dout_mem1[2]
port 117 nsew signal input
flabel metal2 s 142912 0 143024 800 0 FreeSans 448 90 0 0 dout_mem1[30]
port 118 nsew signal input
flabel metal2 s 144592 0 144704 800 0 FreeSans 448 90 0 0 dout_mem1[31]
port 119 nsew signal input
flabel metal2 s 97552 0 97664 800 0 FreeSans 448 90 0 0 dout_mem1[3]
port 120 nsew signal input
flabel metal2 s 99232 0 99344 800 0 FreeSans 448 90 0 0 dout_mem1[4]
port 121 nsew signal input
flabel metal2 s 100912 0 101024 800 0 FreeSans 448 90 0 0 dout_mem1[5]
port 122 nsew signal input
flabel metal2 s 102592 0 102704 800 0 FreeSans 448 90 0 0 dout_mem1[6]
port 123 nsew signal input
flabel metal2 s 104272 0 104384 800 0 FreeSans 448 90 0 0 dout_mem1[7]
port 124 nsew signal input
flabel metal2 s 105952 0 106064 800 0 FreeSans 448 90 0 0 dout_mem1[8]
port 125 nsew signal input
flabel metal2 s 107632 0 107744 800 0 FreeSans 448 90 0 0 dout_mem1[9]
port 126 nsew signal input
flabel metal4 s 19594 3076 19914 36908 0 FreeSans 1280 90 0 0 vdd
port 127 nsew power bidirectional
flabel metal4 s 56414 3076 56734 36908 0 FreeSans 1280 90 0 0 vdd
port 127 nsew power bidirectional
flabel metal4 s 93234 3076 93554 36908 0 FreeSans 1280 90 0 0 vdd
port 127 nsew power bidirectional
flabel metal4 s 130054 3076 130374 36908 0 FreeSans 1280 90 0 0 vdd
port 127 nsew power bidirectional
flabel metal4 s 38004 3076 38324 36908 0 FreeSans 1280 90 0 0 vss
port 128 nsew ground bidirectional
flabel metal4 s 74824 3076 75144 36908 0 FreeSans 1280 90 0 0 vss
port 128 nsew ground bidirectional
flabel metal4 s 111644 3076 111964 36908 0 FreeSans 1280 90 0 0 vss
port 128 nsew ground bidirectional
flabel metal4 s 148464 3076 148784 36908 0 FreeSans 1280 90 0 0 vss
port 128 nsew ground bidirectional
rlabel metal1 74984 36848 74984 36848 0 vdd
rlabel via1 75064 36064 75064 36064 0 vss
rlabel metal2 123256 4760 123256 4760 0 _000_
rlabel metal2 124600 4368 124600 4368 0 _001_
rlabel metal2 125440 4536 125440 4536 0 _002_
rlabel metal3 127624 4536 127624 4536 0 _003_
rlabel metal3 129528 4312 129528 4312 0 _004_
rlabel metal2 130032 3752 130032 3752 0 _005_
rlabel metal2 130760 5208 130760 5208 0 _006_
rlabel metal2 132440 4368 132440 4368 0 _007_
rlabel metal3 133392 4536 133392 4536 0 _008_
rlabel metal2 139608 3920 139608 3920 0 _009_
rlabel metal2 136696 3920 136696 3920 0 _010_
rlabel metal2 138264 4592 138264 4592 0 _011_
rlabel metal2 140336 3752 140336 3752 0 _012_
rlabel metal2 140224 4536 140224 4536 0 _013_
rlabel metal2 143528 4592 143528 4592 0 _014_
rlabel metal2 144200 3920 144200 3920 0 _015_
rlabel metal2 142240 5320 142240 5320 0 _016_
rlabel metal3 142520 4536 142520 4536 0 _017_
rlabel metal2 113288 5040 113288 5040 0 _018_
rlabel metal2 117880 5432 117880 5432 0 _019_
rlabel metal2 100632 4648 100632 4648 0 _020_
rlabel metal2 99456 4536 99456 4536 0 _021_
rlabel metal3 99232 11256 99232 11256 0 _022_
rlabel metal2 101024 3752 101024 3752 0 _023_
rlabel metal2 101416 6468 101416 6468 0 _024_
rlabel metal2 104216 4648 104216 4648 0 _025_
rlabel metal2 103656 4312 103656 4312 0 _026_
rlabel metal2 105000 4368 105000 4368 0 _027_
rlabel metal2 104888 5600 104888 5600 0 _028_
rlabel metal2 106456 4760 106456 4760 0 _029_
rlabel metal3 110264 4312 110264 4312 0 _030_
rlabel metal2 110600 3920 110600 3920 0 _031_
rlabel metal2 112784 3752 112784 3752 0 _032_
rlabel metal2 111832 4536 111832 4536 0 _033_
rlabel metal3 112504 4984 112504 4984 0 _034_
rlabel metal2 118440 3976 118440 3976 0 _035_
rlabel metal2 115640 4368 115640 4368 0 _036_
rlabel metal3 117656 4536 117656 4536 0 _037_
rlabel metal2 119056 4536 119056 4536 0 _038_
rlabel metal2 120680 4144 120680 4144 0 _039_
rlabel metal2 134624 5208 134624 5208 0 _040_
rlabel metal2 124040 3920 124040 3920 0 _041_
rlabel metal2 148120 2744 148120 2744 0 addr[0]
rlabel metal2 147112 3640 147112 3640 0 addr[1]
rlabel metal2 148120 4088 148120 4088 0 addr[2]
rlabel metal2 148120 4928 148120 4928 0 addr[3]
rlabel metal2 148120 5768 148120 5768 0 addr[4]
rlabel metal3 148666 6552 148666 6552 0 addr[5]
rlabel metal2 148120 7784 148120 7784 0 addr[6]
rlabel metal3 148666 8344 148666 8344 0 addr[7]
rlabel metal2 148120 9464 148120 9464 0 addr[8]
rlabel metal2 148120 10360 148120 10360 0 addr[9]
rlabel metal2 6888 854 6888 854 0 addr_mem0[0]
rlabel metal2 8568 2198 8568 2198 0 addr_mem0[1]
rlabel metal2 10248 2198 10248 2198 0 addr_mem0[2]
rlabel metal2 11928 2086 11928 2086 0 addr_mem0[3]
rlabel metal2 13608 2198 13608 2198 0 addr_mem0[4]
rlabel metal2 15288 2086 15288 2086 0 addr_mem0[5]
rlabel metal2 16968 2478 16968 2478 0 addr_mem0[6]
rlabel metal2 18648 2086 18648 2086 0 addr_mem0[7]
rlabel metal2 20328 2086 20328 2086 0 addr_mem0[8]
rlabel metal2 77448 2030 77448 2030 0 addr_mem1[0]
rlabel metal2 79128 2086 79128 2086 0 addr_mem1[1]
rlabel metal2 80808 2142 80808 2142 0 addr_mem1[2]
rlabel metal2 82488 2086 82488 2086 0 addr_mem1[3]
rlabel metal2 84168 2086 84168 2086 0 addr_mem1[4]
rlabel metal2 85848 2478 85848 2478 0 addr_mem1[5]
rlabel metal2 87528 2086 87528 2086 0 addr_mem1[6]
rlabel metal2 89208 2086 89208 2086 0 addr_mem1[7]
rlabel metal2 90888 2030 90888 2030 0 addr_mem1[8]
rlabel metal2 147224 2296 147224 2296 0 csb
rlabel metal2 5208 2086 5208 2086 0 csb_mem0
rlabel metal2 75768 2086 75768 2086 0 csb_mem1
rlabel metal2 147784 11200 147784 11200 0 dout[0]
rlabel metal2 147784 20440 147784 20440 0 dout[10]
rlabel metal2 147784 21168 147784 21168 0 dout[11]
rlabel metal2 147784 22064 147784 22064 0 dout[12]
rlabel metal2 147784 22848 147784 22848 0 dout[13]
rlabel metal2 147784 23744 147784 23744 0 dout[14]
rlabel metal2 147784 24528 147784 24528 0 dout[15]
rlabel metal3 148498 25368 148498 25368 0 dout[16]
rlabel metal2 147784 26600 147784 26600 0 dout[17]
rlabel metal2 147784 27440 147784 27440 0 dout[18]
rlabel metal2 147784 28336 147784 28336 0 dout[19]
rlabel metal2 147784 11984 147784 11984 0 dout[1]
rlabel metal2 147784 29120 147784 29120 0 dout[20]
rlabel metal2 147784 30016 147784 30016 0 dout[21]
rlabel metal2 147784 30800 147784 30800 0 dout[22]
rlabel metal3 148498 31640 148498 31640 0 dout[23]
rlabel metal2 147784 32872 147784 32872 0 dout[24]
rlabel metal2 147784 33824 147784 33824 0 dout[25]
rlabel metal2 147784 34552 147784 34552 0 dout[26]
rlabel metal2 147784 35448 147784 35448 0 dout[27]
rlabel metal2 147784 36288 147784 36288 0 dout[28]
rlabel metal2 145880 36792 145880 36792 0 dout[29]
rlabel metal3 148498 12824 148498 12824 0 dout[2]
rlabel metal2 145992 36848 145992 36848 0 dout[30]
rlabel metal2 146104 36904 146104 36904 0 dout[31]
rlabel metal2 147784 14056 147784 14056 0 dout[3]
rlabel metal2 147784 14896 147784 14896 0 dout[4]
rlabel metal2 147784 15736 147784 15736 0 dout[5]
rlabel metal2 147784 16632 147784 16632 0 dout[6]
rlabel metal2 147784 17472 147784 17472 0 dout[7]
rlabel metal2 147784 18256 147784 18256 0 dout[8]
rlabel metal3 148498 19096 148498 19096 0 dout[9]
rlabel metal2 21896 4200 21896 4200 0 dout_mem0[0]
rlabel metal2 38696 3416 38696 3416 0 dout_mem0[10]
rlabel metal2 40432 3416 40432 3416 0 dout_mem0[11]
rlabel metal2 42056 3416 42056 3416 0 dout_mem0[12]
rlabel metal2 43848 2086 43848 2086 0 dout_mem0[13]
rlabel metal2 45416 3416 45416 3416 0 dout_mem0[14]
rlabel metal2 47096 3416 47096 3416 0 dout_mem0[15]
rlabel metal2 49000 3416 49000 3416 0 dout_mem0[16]
rlabel metal2 50456 3416 50456 3416 0 dout_mem0[17]
rlabel metal2 52192 3416 52192 3416 0 dout_mem0[18]
rlabel metal2 53816 3416 53816 3416 0 dout_mem0[19]
rlabel metal2 23576 3416 23576 3416 0 dout_mem0[1]
rlabel metal2 55608 2086 55608 2086 0 dout_mem0[20]
rlabel metal2 57176 3416 57176 3416 0 dout_mem0[21]
rlabel metal2 58856 3416 58856 3416 0 dout_mem0[22]
rlabel metal2 60760 3416 60760 3416 0 dout_mem0[23]
rlabel metal2 62216 3416 62216 3416 0 dout_mem0[24]
rlabel metal2 63952 3416 63952 3416 0 dout_mem0[25]
rlabel metal2 65576 3416 65576 3416 0 dout_mem0[26]
rlabel metal2 67368 2086 67368 2086 0 dout_mem0[27]
rlabel metal2 68936 3416 68936 3416 0 dout_mem0[28]
rlabel metal2 70616 3416 70616 3416 0 dout_mem0[29]
rlabel metal2 25480 3416 25480 3416 0 dout_mem0[2]
rlabel metal2 72464 3416 72464 3416 0 dout_mem0[30]
rlabel metal2 74200 3416 74200 3416 0 dout_mem0[31]
rlabel metal2 26936 3416 26936 3416 0 dout_mem0[3]
rlabel metal2 28672 3416 28672 3416 0 dout_mem0[4]
rlabel metal2 30296 3416 30296 3416 0 dout_mem0[5]
rlabel metal2 32088 2086 32088 2086 0 dout_mem0[6]
rlabel metal2 33656 3416 33656 3416 0 dout_mem0[7]
rlabel metal2 35336 3416 35336 3416 0 dout_mem0[8]
rlabel metal2 37240 3416 37240 3416 0 dout_mem0[9]
rlabel metal3 93184 3528 93184 3528 0 dout_mem1[0]
rlabel metal2 109424 4312 109424 4312 0 dout_mem1[10]
rlabel metal3 112448 3416 112448 3416 0 dout_mem1[11]
rlabel metal2 114184 5712 114184 5712 0 dout_mem1[12]
rlabel metal2 114632 4928 114632 4928 0 dout_mem1[13]
rlabel metal3 116928 3416 116928 3416 0 dout_mem1[14]
rlabel metal2 118328 4592 118328 4592 0 dout_mem1[15]
rlabel metal2 119560 4312 119560 4312 0 dout_mem1[16]
rlabel metal2 121240 3416 121240 3416 0 dout_mem1[17]
rlabel metal3 122528 3416 122528 3416 0 dout_mem1[18]
rlabel metal3 125048 3416 125048 3416 0 dout_mem1[19]
rlabel metal2 94472 3416 94472 3416 0 dout_mem1[1]
rlabel metal3 126840 3528 126840 3528 0 dout_mem1[20]
rlabel metal2 127904 4312 127904 4312 0 dout_mem1[21]
rlabel metal2 129416 5768 129416 5768 0 dout_mem1[22]
rlabel metal3 132328 3416 132328 3416 0 dout_mem1[23]
rlabel metal2 134232 2128 134232 2128 0 dout_mem1[24]
rlabel metal2 134680 4312 134680 4312 0 dout_mem1[25]
rlabel metal3 136808 3416 136808 3416 0 dout_mem1[26]
rlabel metal3 139552 3528 139552 3528 0 dout_mem1[27]
rlabel metal3 140952 3416 140952 3416 0 dout_mem1[28]
rlabel metal2 142856 4256 142856 4256 0 dout_mem1[29]
rlabel metal2 96040 3416 96040 3416 0 dout_mem1[2]
rlabel metal3 143528 4312 143528 4312 0 dout_mem1[30]
rlabel metal2 144872 3528 144872 3528 0 dout_mem1[31]
rlabel metal2 97496 4312 97496 4312 0 dout_mem1[3]
rlabel metal2 99176 5096 99176 5096 0 dout_mem1[4]
rlabel metal2 101752 2072 101752 2072 0 dout_mem1[5]
rlabel metal2 102648 2086 102648 2086 0 dout_mem1[6]
rlabel metal3 105224 3416 105224 3416 0 dout_mem1[7]
rlabel metal3 106456 3528 106456 3528 0 dout_mem1[8]
rlabel metal2 107800 3416 107800 3416 0 dout_mem1[9]
rlabel metal2 77672 5936 77672 5936 0 net1
rlabel metal2 147672 10696 147672 10696 0 net10
rlabel metal3 119112 4984 119112 4984 0 net100
rlabel metal2 118552 5880 118552 5880 0 net101
rlabel metal2 146888 24640 146888 24640 0 net102
rlabel metal2 146888 25368 146888 25368 0 net103
rlabel metal2 123984 4984 123984 4984 0 net104
rlabel metal2 125384 6272 125384 6272 0 net105
rlabel metal3 142800 28616 142800 28616 0 net106
rlabel metal2 99624 8904 99624 8904 0 net107
rlabel metal3 146664 29400 146664 29400 0 net108
rlabel metal3 137816 4592 137816 4592 0 net109
rlabel metal2 76104 5376 76104 5376 0 net11
rlabel metal3 146664 30968 146664 30968 0 net110
rlabel metal2 146888 31640 146888 31640 0 net111
rlabel metal3 146608 33320 146608 33320 0 net112
rlabel metal2 137816 5880 137816 5880 0 net113
rlabel metal2 139496 5824 139496 5824 0 net114
rlabel metal2 145432 33936 145432 33936 0 net115
rlabel metal3 142800 36232 142800 36232 0 net116
rlabel metal2 144200 36232 144200 36232 0 net117
rlabel metal2 99848 12096 99848 12096 0 net118
rlabel metal3 143472 35560 143472 35560 0 net119
rlabel metal2 22568 5656 22568 5656 0 net12
rlabel metal2 144536 34104 144536 34104 0 net120
rlabel metal2 100744 13440 100744 13440 0 net121
rlabel metal2 101864 14112 101864 14112 0 net122
rlabel metal2 146888 15960 146888 15960 0 net123
rlabel metal2 116648 13552 116648 13552 0 net124
rlabel metal2 119224 15848 119224 15848 0 net125
rlabel metal2 146888 18368 146888 18368 0 net126
rlabel metal3 146608 19208 146608 19208 0 net127
rlabel metal3 40936 3304 40936 3304 0 net13
rlabel metal3 111384 4536 111384 4536 0 net14
rlabel metal2 111048 5096 111048 5096 0 net15
rlabel metal2 44184 2240 44184 2240 0 net16
rlabel metal2 46088 2296 46088 2296 0 net17
rlabel metal2 47768 2072 47768 2072 0 net18
rlabel metal2 49448 2352 49448 2352 0 net19
rlabel metal2 78904 2968 78904 2968 0 net2
rlabel metal2 51128 5488 51128 5488 0 net20
rlabel metal2 53144 5880 53144 5880 0 net21
rlabel metal2 124376 2800 124376 2800 0 net22
rlabel metal2 24248 2408 24248 2408 0 net23
rlabel metal2 125944 5264 125944 5264 0 net24
rlabel metal2 64120 2128 64120 2128 0 net25
rlabel metal3 128520 6552 128520 6552 0 net26
rlabel metal2 121016 3136 121016 3136 0 net27
rlabel metal2 62888 3136 62888 3136 0 net28
rlabel metal2 64904 2912 64904 2912 0 net29
rlabel metal3 146944 4536 146944 4536 0 net3
rlabel metal3 95816 4032 95816 4032 0 net30
rlabel metal2 67704 2688 67704 2688 0 net31
rlabel metal2 69608 2744 69608 2744 0 net32
rlabel metal2 71288 5096 71288 5096 0 net33
rlabel metal3 28336 3304 28336 3304 0 net34
rlabel metal2 72856 3528 72856 3528 0 net35
rlabel metal2 74648 3080 74648 3080 0 net36
rlabel metal2 27608 3136 27608 3136 0 net37
rlabel metal2 29624 3080 29624 3080 0 net38
rlabel metal2 30968 3024 30968 3024 0 net39
rlabel metal2 147784 4816 147784 4816 0 net4
rlabel metal2 32424 2912 32424 2912 0 net40
rlabel metal2 34328 2856 34328 2856 0 net41
rlabel metal2 36008 4928 36008 4928 0 net42
rlabel metal3 38416 3304 38416 3304 0 net43
rlabel metal2 94136 2800 94136 2800 0 net44
rlabel metal2 112504 4088 112504 4088 0 net45
rlabel metal3 112392 3304 112392 3304 0 net46
rlabel metal2 114072 3640 114072 3640 0 net47
rlabel metal2 115976 3808 115976 3808 0 net48
rlabel metal2 116928 4088 116928 4088 0 net49
rlabel metal2 85400 5264 85400 5264 0 net5
rlabel metal2 118664 3752 118664 3752 0 net50
rlabel metal2 120344 4088 120344 4088 0 net51
rlabel metal2 121688 3696 121688 3696 0 net52
rlabel metal2 122584 3416 122584 3416 0 net53
rlabel metal2 125272 3752 125272 3752 0 net54
rlabel metal3 97104 3304 97104 3304 0 net55
rlabel metal2 127232 3416 127232 3416 0 net56
rlabel metal2 129752 3808 129752 3808 0 net57
rlabel metal2 130424 4760 130424 4760 0 net58
rlabel metal3 132608 3304 132608 3304 0 net59
rlabel metal2 147784 6384 147784 6384 0 net6
rlabel metal2 134008 3248 134008 3248 0 net60
rlabel metal2 136360 4088 136360 4088 0 net61
rlabel metal2 137704 3696 137704 3696 0 net62
rlabel metal2 140952 3136 140952 3136 0 net63
rlabel metal3 140952 3304 140952 3304 0 net64
rlabel metal3 143528 3752 143528 3752 0 net65
rlabel metal2 96488 3416 96488 3416 0 net66
rlabel metal2 143752 4592 143752 4592 0 net67
rlabel metal3 143472 3304 143472 3304 0 net68
rlabel metal2 100744 4088 100744 4088 0 net69
rlabel metal2 147784 7616 147784 7616 0 net7
rlabel metal3 100464 4312 100464 4312 0 net70
rlabel metal2 102088 3696 102088 3696 0 net71
rlabel metal2 102984 3416 102984 3416 0 net72
rlabel metal2 105672 3136 105672 3136 0 net73
rlabel metal2 106568 3752 106568 3752 0 net74
rlabel metal2 108248 3416 108248 3416 0 net75
rlabel metal2 75208 4200 75208 4200 0 net76
rlabel metal2 77896 5152 77896 5152 0 net77
rlabel metal3 11592 4536 11592 4536 0 net78
rlabel metal3 13272 4536 13272 4536 0 net79
rlabel metal2 90776 7168 90776 7168 0 net8
rlabel metal2 15064 3528 15064 3528 0 net80
rlabel metal3 17136 3528 17136 3528 0 net81
rlabel metal2 18984 4368 18984 4368 0 net82
rlabel metal2 21672 5376 21672 5376 0 net83
rlabel metal2 22680 3584 22680 3584 0 net84
rlabel metal2 77336 3976 77336 3976 0 net85
rlabel metal2 79184 4424 79184 4424 0 net86
rlabel metal2 81704 3976 81704 3976 0 net87
rlabel metal2 82376 4592 82376 4592 0 net88
rlabel metal2 84840 3976 84840 3976 0 net89
rlabel metal2 147672 9184 147672 9184 0 net9
rlabel metal2 86184 3864 86184 3864 0 net90
rlabel metal2 88200 3976 88200 3976 0 net91
rlabel metal2 89656 3976 89656 3976 0 net92
rlabel metal2 90776 3976 90776 3976 0 net93
rlabel metal2 6720 3528 6720 3528 0 net94
rlabel metal2 75768 4424 75768 4424 0 net95
rlabel metal2 115976 9576 115976 9576 0 net96
rlabel metal3 146608 20776 146608 20776 0 net97
rlabel metal2 146888 21504 146888 21504 0 net98
rlabel metal3 146608 22344 146608 22344 0 net99
<< properties >>
string FIXED_BBOX 0 0 150000 40000
<< end >>
