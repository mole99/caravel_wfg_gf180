VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wfg_top
  CLASS BLOCK ;
  FOREIGN wfg_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 800.000 ;
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.680 4.000 30.240 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.160 4.000 48.720 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.640 4.000 67.200 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 85.120 4.000 85.680 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 103.600 4.000 104.160 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 122.080 4.000 122.640 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.560 4.000 141.120 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 159.040 4.000 159.600 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 177.520 4.000 178.080 ;
    END
  END addr1[8]
  PIN addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 196.000 4.000 196.560 ;
    END
  END addr1[9]
  PIN csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.200 4.000 11.760 ;
    END
  END csb1
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.480 4.000 215.040 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 399.280 4.000 399.840 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 417.760 4.000 418.320 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 436.240 4.000 436.800 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 454.720 4.000 455.280 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 473.200 4.000 473.760 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 491.680 4.000 492.240 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 510.160 4.000 510.720 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 528.640 4.000 529.200 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 547.120 4.000 547.680 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 565.600 4.000 566.160 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.960 4.000 233.520 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 584.080 4.000 584.640 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 602.560 4.000 603.120 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 621.040 4.000 621.600 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 639.520 4.000 640.080 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 658.000 4.000 658.560 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 676.480 4.000 677.040 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 694.960 4.000 695.520 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 713.440 4.000 714.000 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 731.920 4.000 732.480 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 750.400 4.000 750.960 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 251.440 4.000 252.000 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 768.880 4.000 769.440 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 787.360 4.000 787.920 ;
    END
  END dout1[31]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 269.920 4.000 270.480 ;
    END
  END dout1[3]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 288.400 4.000 288.960 ;
    END
  END dout1[4]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 306.880 4.000 307.440 ;
    END
  END dout1[5]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 325.360 4.000 325.920 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 343.840 4.000 344.400 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.320 4.000 362.880 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.800 4.000 381.360 ;
    END
  END dout1[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 616.560 796.000 617.120 800.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 790.160 796.000 790.720 800.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 796.000 634.480 800.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 651.280 796.000 651.840 800.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 796.000 669.200 800.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 686.000 796.000 686.560 800.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 703.360 796.000 703.920 800.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.720 796.000 721.280 800.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 738.080 796.000 738.640 800.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 755.440 796.000 756.000 800.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 796.000 773.360 800.000 ;
    END
  END io_oeb[9]
  PIN io_wbs_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END io_wbs_ack
  PIN io_wbs_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END io_wbs_adr[0]
  PIN io_wbs_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 0.000 286.160 4.000 ;
    END
  END io_wbs_adr[10]
  PIN io_wbs_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 0.000 309.680 4.000 ;
    END
  END io_wbs_adr[11]
  PIN io_wbs_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 0.000 333.200 4.000 ;
    END
  END io_wbs_adr[12]
  PIN io_wbs_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 0.000 356.720 4.000 ;
    END
  END io_wbs_adr[13]
  PIN io_wbs_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 0.000 380.240 4.000 ;
    END
  END io_wbs_adr[14]
  PIN io_wbs_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 0.000 403.760 4.000 ;
    END
  END io_wbs_adr[15]
  PIN io_wbs_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 0.000 427.280 4.000 ;
    END
  END io_wbs_adr[16]
  PIN io_wbs_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 0.000 450.800 4.000 ;
    END
  END io_wbs_adr[17]
  PIN io_wbs_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 0.000 474.320 4.000 ;
    END
  END io_wbs_adr[18]
  PIN io_wbs_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 0.000 497.840 4.000 ;
    END
  END io_wbs_adr[19]
  PIN io_wbs_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END io_wbs_adr[1]
  PIN io_wbs_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 0.000 521.360 4.000 ;
    END
  END io_wbs_adr[20]
  PIN io_wbs_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 0.000 544.880 4.000 ;
    END
  END io_wbs_adr[21]
  PIN io_wbs_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 0.000 568.400 4.000 ;
    END
  END io_wbs_adr[22]
  PIN io_wbs_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 0.000 591.920 4.000 ;
    END
  END io_wbs_adr[23]
  PIN io_wbs_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 0.000 615.440 4.000 ;
    END
  END io_wbs_adr[24]
  PIN io_wbs_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 0.000 638.960 4.000 ;
    END
  END io_wbs_adr[25]
  PIN io_wbs_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 0.000 662.480 4.000 ;
    END
  END io_wbs_adr[26]
  PIN io_wbs_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 0.000 686.000 4.000 ;
    END
  END io_wbs_adr[27]
  PIN io_wbs_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 708.960 0.000 709.520 4.000 ;
    END
  END io_wbs_adr[28]
  PIN io_wbs_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 0.000 733.040 4.000 ;
    END
  END io_wbs_adr[29]
  PIN io_wbs_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END io_wbs_adr[2]
  PIN io_wbs_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 756.000 0.000 756.560 4.000 ;
    END
  END io_wbs_adr[30]
  PIN io_wbs_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 0.000 780.080 4.000 ;
    END
  END io_wbs_adr[31]
  PIN io_wbs_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 0.000 121.520 4.000 ;
    END
  END io_wbs_adr[3]
  PIN io_wbs_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END io_wbs_adr[4]
  PIN io_wbs_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END io_wbs_adr[5]
  PIN io_wbs_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END io_wbs_adr[6]
  PIN io_wbs_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 0.000 215.600 4.000 ;
    END
  END io_wbs_adr[7]
  PIN io_wbs_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 4.000 ;
    END
  END io_wbs_adr[8]
  PIN io_wbs_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 0.000 262.640 4.000 ;
    END
  END io_wbs_adr[9]
  PIN io_wbs_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 11.200 0.000 11.760 4.000 ;
    END
  END io_wbs_clk
  PIN io_wbs_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 0.000 19.600 4.000 ;
    END
  END io_wbs_cyc
  PIN io_wbs_datrd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 0.000 58.800 4.000 ;
    END
  END io_wbs_datrd[0]
  PIN io_wbs_datrd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 0.000 294.000 4.000 ;
    END
  END io_wbs_datrd[10]
  PIN io_wbs_datrd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 0.000 317.520 4.000 ;
    END
  END io_wbs_datrd[11]
  PIN io_wbs_datrd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 0.000 341.040 4.000 ;
    END
  END io_wbs_datrd[12]
  PIN io_wbs_datrd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 0.000 364.560 4.000 ;
    END
  END io_wbs_datrd[13]
  PIN io_wbs_datrd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 0.000 388.080 4.000 ;
    END
  END io_wbs_datrd[14]
  PIN io_wbs_datrd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 0.000 411.600 4.000 ;
    END
  END io_wbs_datrd[15]
  PIN io_wbs_datrd[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 434.560 0.000 435.120 4.000 ;
    END
  END io_wbs_datrd[16]
  PIN io_wbs_datrd[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 0.000 458.640 4.000 ;
    END
  END io_wbs_datrd[17]
  PIN io_wbs_datrd[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 0.000 482.160 4.000 ;
    END
  END io_wbs_datrd[18]
  PIN io_wbs_datrd[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 0.000 505.680 4.000 ;
    END
  END io_wbs_datrd[19]
  PIN io_wbs_datrd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 0.000 82.320 4.000 ;
    END
  END io_wbs_datrd[1]
  PIN io_wbs_datrd[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 528.640 0.000 529.200 4.000 ;
    END
  END io_wbs_datrd[20]
  PIN io_wbs_datrd[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 552.160 0.000 552.720 4.000 ;
    END
  END io_wbs_datrd[21]
  PIN io_wbs_datrd[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 0.000 576.240 4.000 ;
    END
  END io_wbs_datrd[22]
  PIN io_wbs_datrd[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 0.000 599.760 4.000 ;
    END
  END io_wbs_datrd[23]
  PIN io_wbs_datrd[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 622.720 0.000 623.280 4.000 ;
    END
  END io_wbs_datrd[24]
  PIN io_wbs_datrd[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 646.240 0.000 646.800 4.000 ;
    END
  END io_wbs_datrd[25]
  PIN io_wbs_datrd[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 669.760 0.000 670.320 4.000 ;
    END
  END io_wbs_datrd[26]
  PIN io_wbs_datrd[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 693.280 0.000 693.840 4.000 ;
    END
  END io_wbs_datrd[27]
  PIN io_wbs_datrd[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 716.800 0.000 717.360 4.000 ;
    END
  END io_wbs_datrd[28]
  PIN io_wbs_datrd[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 740.320 0.000 740.880 4.000 ;
    END
  END io_wbs_datrd[29]
  PIN io_wbs_datrd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 0.000 105.840 4.000 ;
    END
  END io_wbs_datrd[2]
  PIN io_wbs_datrd[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 763.840 0.000 764.400 4.000 ;
    END
  END io_wbs_datrd[30]
  PIN io_wbs_datrd[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 787.360 0.000 787.920 4.000 ;
    END
  END io_wbs_datrd[31]
  PIN io_wbs_datrd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 4.000 ;
    END
  END io_wbs_datrd[3]
  PIN io_wbs_datrd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 0.000 152.880 4.000 ;
    END
  END io_wbs_datrd[4]
  PIN io_wbs_datrd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 0.000 176.400 4.000 ;
    END
  END io_wbs_datrd[5]
  PIN io_wbs_datrd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 0.000 199.920 4.000 ;
    END
  END io_wbs_datrd[6]
  PIN io_wbs_datrd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 4.000 ;
    END
  END io_wbs_datrd[7]
  PIN io_wbs_datrd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 0.000 246.960 4.000 ;
    END
  END io_wbs_datrd[8]
  PIN io_wbs_datrd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 0.000 270.480 4.000 ;
    END
  END io_wbs_datrd[9]
  PIN io_wbs_datwr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 4.000 ;
    END
  END io_wbs_datwr[0]
  PIN io_wbs_datwr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 301.280 0.000 301.840 4.000 ;
    END
  END io_wbs_datwr[10]
  PIN io_wbs_datwr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 0.000 325.360 4.000 ;
    END
  END io_wbs_datwr[11]
  PIN io_wbs_datwr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 0.000 348.880 4.000 ;
    END
  END io_wbs_datwr[12]
  PIN io_wbs_datwr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.840 0.000 372.400 4.000 ;
    END
  END io_wbs_datwr[13]
  PIN io_wbs_datwr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 395.360 0.000 395.920 4.000 ;
    END
  END io_wbs_datwr[14]
  PIN io_wbs_datwr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 0.000 419.440 4.000 ;
    END
  END io_wbs_datwr[15]
  PIN io_wbs_datwr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 442.400 0.000 442.960 4.000 ;
    END
  END io_wbs_datwr[16]
  PIN io_wbs_datwr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 465.920 0.000 466.480 4.000 ;
    END
  END io_wbs_datwr[17]
  PIN io_wbs_datwr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 489.440 0.000 490.000 4.000 ;
    END
  END io_wbs_datwr[18]
  PIN io_wbs_datwr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 512.960 0.000 513.520 4.000 ;
    END
  END io_wbs_datwr[19]
  PIN io_wbs_datwr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 0.000 90.160 4.000 ;
    END
  END io_wbs_datwr[1]
  PIN io_wbs_datwr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 536.480 0.000 537.040 4.000 ;
    END
  END io_wbs_datwr[20]
  PIN io_wbs_datwr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 560.000 0.000 560.560 4.000 ;
    END
  END io_wbs_datwr[21]
  PIN io_wbs_datwr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 583.520 0.000 584.080 4.000 ;
    END
  END io_wbs_datwr[22]
  PIN io_wbs_datwr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 607.040 0.000 607.600 4.000 ;
    END
  END io_wbs_datwr[23]
  PIN io_wbs_datwr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 630.560 0.000 631.120 4.000 ;
    END
  END io_wbs_datwr[24]
  PIN io_wbs_datwr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 654.080 0.000 654.640 4.000 ;
    END
  END io_wbs_datwr[25]
  PIN io_wbs_datwr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 677.600 0.000 678.160 4.000 ;
    END
  END io_wbs_datwr[26]
  PIN io_wbs_datwr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 701.120 0.000 701.680 4.000 ;
    END
  END io_wbs_datwr[27]
  PIN io_wbs_datwr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 724.640 0.000 725.200 4.000 ;
    END
  END io_wbs_datwr[28]
  PIN io_wbs_datwr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 748.160 0.000 748.720 4.000 ;
    END
  END io_wbs_datwr[29]
  PIN io_wbs_datwr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 0.000 113.680 4.000 ;
    END
  END io_wbs_datwr[2]
  PIN io_wbs_datwr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 771.680 0.000 772.240 4.000 ;
    END
  END io_wbs_datwr[30]
  PIN io_wbs_datwr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 795.200 0.000 795.760 4.000 ;
    END
  END io_wbs_datwr[31]
  PIN io_wbs_datwr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 0.000 137.200 4.000 ;
    END
  END io_wbs_datwr[3]
  PIN io_wbs_datwr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 0.000 160.720 4.000 ;
    END
  END io_wbs_datwr[4]
  PIN io_wbs_datwr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 0.000 184.240 4.000 ;
    END
  END io_wbs_datwr[5]
  PIN io_wbs_datwr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 0.000 207.760 4.000 ;
    END
  END io_wbs_datwr[6]
  PIN io_wbs_datwr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 0.000 231.280 4.000 ;
    END
  END io_wbs_datwr[7]
  PIN io_wbs_datwr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 0.000 254.800 4.000 ;
    END
  END io_wbs_datwr[8]
  PIN io_wbs_datwr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 0.000 278.320 4.000 ;
    END
  END io_wbs_datwr[9]
  PIN io_wbs_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END io_wbs_rst
  PIN io_wbs_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 0.000 35.280 4.000 ;
    END
  END io_wbs_stb
  PIN io_wbs_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 0.000 43.120 4.000 ;
    END
  END io_wbs_we
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 784.300 ;
    END
  END vss
  PIN wfg_drive_pat_dout_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.040 796.000 61.600 800.000 ;
    END
  END wfg_drive_pat_dout_o[0]
  PIN wfg_drive_pat_dout_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.640 796.000 235.200 800.000 ;
    END
  END wfg_drive_pat_dout_o[10]
  PIN wfg_drive_pat_dout_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 796.000 252.560 800.000 ;
    END
  END wfg_drive_pat_dout_o[11]
  PIN wfg_drive_pat_dout_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.360 796.000 269.920 800.000 ;
    END
  END wfg_drive_pat_dout_o[12]
  PIN wfg_drive_pat_dout_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 796.000 287.280 800.000 ;
    END
  END wfg_drive_pat_dout_o[13]
  PIN wfg_drive_pat_dout_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.080 796.000 304.640 800.000 ;
    END
  END wfg_drive_pat_dout_o[14]
  PIN wfg_drive_pat_dout_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 796.000 322.000 800.000 ;
    END
  END wfg_drive_pat_dout_o[15]
  PIN wfg_drive_pat_dout_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.800 796.000 339.360 800.000 ;
    END
  END wfg_drive_pat_dout_o[16]
  PIN wfg_drive_pat_dout_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 796.000 356.720 800.000 ;
    END
  END wfg_drive_pat_dout_o[17]
  PIN wfg_drive_pat_dout_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 373.520 796.000 374.080 800.000 ;
    END
  END wfg_drive_pat_dout_o[18]
  PIN wfg_drive_pat_dout_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 796.000 391.440 800.000 ;
    END
  END wfg_drive_pat_dout_o[19]
  PIN wfg_drive_pat_dout_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 796.000 78.960 800.000 ;
    END
  END wfg_drive_pat_dout_o[1]
  PIN wfg_drive_pat_dout_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 408.240 796.000 408.800 800.000 ;
    END
  END wfg_drive_pat_dout_o[20]
  PIN wfg_drive_pat_dout_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 425.600 796.000 426.160 800.000 ;
    END
  END wfg_drive_pat_dout_o[21]
  PIN wfg_drive_pat_dout_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 442.960 796.000 443.520 800.000 ;
    END
  END wfg_drive_pat_dout_o[22]
  PIN wfg_drive_pat_dout_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 796.000 460.880 800.000 ;
    END
  END wfg_drive_pat_dout_o[23]
  PIN wfg_drive_pat_dout_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.680 796.000 478.240 800.000 ;
    END
  END wfg_drive_pat_dout_o[24]
  PIN wfg_drive_pat_dout_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 495.040 796.000 495.600 800.000 ;
    END
  END wfg_drive_pat_dout_o[25]
  PIN wfg_drive_pat_dout_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 512.400 796.000 512.960 800.000 ;
    END
  END wfg_drive_pat_dout_o[26]
  PIN wfg_drive_pat_dout_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 796.000 530.320 800.000 ;
    END
  END wfg_drive_pat_dout_o[27]
  PIN wfg_drive_pat_dout_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.120 796.000 547.680 800.000 ;
    END
  END wfg_drive_pat_dout_o[28]
  PIN wfg_drive_pat_dout_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 796.000 565.040 800.000 ;
    END
  END wfg_drive_pat_dout_o[29]
  PIN wfg_drive_pat_dout_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.760 796.000 96.320 800.000 ;
    END
  END wfg_drive_pat_dout_o[2]
  PIN wfg_drive_pat_dout_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.840 796.000 582.400 800.000 ;
    END
  END wfg_drive_pat_dout_o[30]
  PIN wfg_drive_pat_dout_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 796.000 599.760 800.000 ;
    END
  END wfg_drive_pat_dout_o[31]
  PIN wfg_drive_pat_dout_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 796.000 113.680 800.000 ;
    END
  END wfg_drive_pat_dout_o[3]
  PIN wfg_drive_pat_dout_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.480 796.000 131.040 800.000 ;
    END
  END wfg_drive_pat_dout_o[4]
  PIN wfg_drive_pat_dout_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 796.000 148.400 800.000 ;
    END
  END wfg_drive_pat_dout_o[5]
  PIN wfg_drive_pat_dout_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 165.200 796.000 165.760 800.000 ;
    END
  END wfg_drive_pat_dout_o[6]
  PIN wfg_drive_pat_dout_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 796.000 183.120 800.000 ;
    END
  END wfg_drive_pat_dout_o[7]
  PIN wfg_drive_pat_dout_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.920 796.000 200.480 800.000 ;
    END
  END wfg_drive_pat_dout_o[8]
  PIN wfg_drive_pat_dout_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 796.000 217.840 800.000 ;
    END
  END wfg_drive_pat_dout_o[9]
  PIN wfg_drive_spi_cs_no
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 8.960 796.000 9.520 800.000 ;
    END
  END wfg_drive_spi_cs_no
  PIN wfg_drive_spi_sclk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.320 796.000 26.880 800.000 ;
    END
  END wfg_drive_spi_sclk_o
  PIN wfg_drive_spi_sdo_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 796.000 44.240 800.000 ;
    END
  END wfg_drive_spi_sdo_o
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 797.350 788.890 ;
      LAYER Metal2 ;
        RECT 0.140 795.700 8.660 796.000 ;
        RECT 9.820 795.700 26.020 796.000 ;
        RECT 27.180 795.700 43.380 796.000 ;
        RECT 44.540 795.700 60.740 796.000 ;
        RECT 61.900 795.700 78.100 796.000 ;
        RECT 79.260 795.700 95.460 796.000 ;
        RECT 96.620 795.700 112.820 796.000 ;
        RECT 113.980 795.700 130.180 796.000 ;
        RECT 131.340 795.700 147.540 796.000 ;
        RECT 148.700 795.700 164.900 796.000 ;
        RECT 166.060 795.700 182.260 796.000 ;
        RECT 183.420 795.700 199.620 796.000 ;
        RECT 200.780 795.700 216.980 796.000 ;
        RECT 218.140 795.700 234.340 796.000 ;
        RECT 235.500 795.700 251.700 796.000 ;
        RECT 252.860 795.700 269.060 796.000 ;
        RECT 270.220 795.700 286.420 796.000 ;
        RECT 287.580 795.700 303.780 796.000 ;
        RECT 304.940 795.700 321.140 796.000 ;
        RECT 322.300 795.700 338.500 796.000 ;
        RECT 339.660 795.700 355.860 796.000 ;
        RECT 357.020 795.700 373.220 796.000 ;
        RECT 374.380 795.700 390.580 796.000 ;
        RECT 391.740 795.700 407.940 796.000 ;
        RECT 409.100 795.700 425.300 796.000 ;
        RECT 426.460 795.700 442.660 796.000 ;
        RECT 443.820 795.700 460.020 796.000 ;
        RECT 461.180 795.700 477.380 796.000 ;
        RECT 478.540 795.700 494.740 796.000 ;
        RECT 495.900 795.700 512.100 796.000 ;
        RECT 513.260 795.700 529.460 796.000 ;
        RECT 530.620 795.700 546.820 796.000 ;
        RECT 547.980 795.700 564.180 796.000 ;
        RECT 565.340 795.700 581.540 796.000 ;
        RECT 582.700 795.700 598.900 796.000 ;
        RECT 600.060 795.700 616.260 796.000 ;
        RECT 617.420 795.700 633.620 796.000 ;
        RECT 634.780 795.700 650.980 796.000 ;
        RECT 652.140 795.700 668.340 796.000 ;
        RECT 669.500 795.700 685.700 796.000 ;
        RECT 686.860 795.700 703.060 796.000 ;
        RECT 704.220 795.700 720.420 796.000 ;
        RECT 721.580 795.700 737.780 796.000 ;
        RECT 738.940 795.700 755.140 796.000 ;
        RECT 756.300 795.700 772.500 796.000 ;
        RECT 773.660 795.700 789.860 796.000 ;
        RECT 791.020 795.700 797.300 796.000 ;
        RECT 0.140 4.300 797.300 795.700 ;
        RECT 0.140 4.000 3.060 4.300 ;
        RECT 4.220 4.000 10.900 4.300 ;
        RECT 12.060 4.000 18.740 4.300 ;
        RECT 19.900 4.000 26.580 4.300 ;
        RECT 27.740 4.000 34.420 4.300 ;
        RECT 35.580 4.000 42.260 4.300 ;
        RECT 43.420 4.000 50.100 4.300 ;
        RECT 51.260 4.000 57.940 4.300 ;
        RECT 59.100 4.000 65.780 4.300 ;
        RECT 66.940 4.000 73.620 4.300 ;
        RECT 74.780 4.000 81.460 4.300 ;
        RECT 82.620 4.000 89.300 4.300 ;
        RECT 90.460 4.000 97.140 4.300 ;
        RECT 98.300 4.000 104.980 4.300 ;
        RECT 106.140 4.000 112.820 4.300 ;
        RECT 113.980 4.000 120.660 4.300 ;
        RECT 121.820 4.000 128.500 4.300 ;
        RECT 129.660 4.000 136.340 4.300 ;
        RECT 137.500 4.000 144.180 4.300 ;
        RECT 145.340 4.000 152.020 4.300 ;
        RECT 153.180 4.000 159.860 4.300 ;
        RECT 161.020 4.000 167.700 4.300 ;
        RECT 168.860 4.000 175.540 4.300 ;
        RECT 176.700 4.000 183.380 4.300 ;
        RECT 184.540 4.000 191.220 4.300 ;
        RECT 192.380 4.000 199.060 4.300 ;
        RECT 200.220 4.000 206.900 4.300 ;
        RECT 208.060 4.000 214.740 4.300 ;
        RECT 215.900 4.000 222.580 4.300 ;
        RECT 223.740 4.000 230.420 4.300 ;
        RECT 231.580 4.000 238.260 4.300 ;
        RECT 239.420 4.000 246.100 4.300 ;
        RECT 247.260 4.000 253.940 4.300 ;
        RECT 255.100 4.000 261.780 4.300 ;
        RECT 262.940 4.000 269.620 4.300 ;
        RECT 270.780 4.000 277.460 4.300 ;
        RECT 278.620 4.000 285.300 4.300 ;
        RECT 286.460 4.000 293.140 4.300 ;
        RECT 294.300 4.000 300.980 4.300 ;
        RECT 302.140 4.000 308.820 4.300 ;
        RECT 309.980 4.000 316.660 4.300 ;
        RECT 317.820 4.000 324.500 4.300 ;
        RECT 325.660 4.000 332.340 4.300 ;
        RECT 333.500 4.000 340.180 4.300 ;
        RECT 341.340 4.000 348.020 4.300 ;
        RECT 349.180 4.000 355.860 4.300 ;
        RECT 357.020 4.000 363.700 4.300 ;
        RECT 364.860 4.000 371.540 4.300 ;
        RECT 372.700 4.000 379.380 4.300 ;
        RECT 380.540 4.000 387.220 4.300 ;
        RECT 388.380 4.000 395.060 4.300 ;
        RECT 396.220 4.000 402.900 4.300 ;
        RECT 404.060 4.000 410.740 4.300 ;
        RECT 411.900 4.000 418.580 4.300 ;
        RECT 419.740 4.000 426.420 4.300 ;
        RECT 427.580 4.000 434.260 4.300 ;
        RECT 435.420 4.000 442.100 4.300 ;
        RECT 443.260 4.000 449.940 4.300 ;
        RECT 451.100 4.000 457.780 4.300 ;
        RECT 458.940 4.000 465.620 4.300 ;
        RECT 466.780 4.000 473.460 4.300 ;
        RECT 474.620 4.000 481.300 4.300 ;
        RECT 482.460 4.000 489.140 4.300 ;
        RECT 490.300 4.000 496.980 4.300 ;
        RECT 498.140 4.000 504.820 4.300 ;
        RECT 505.980 4.000 512.660 4.300 ;
        RECT 513.820 4.000 520.500 4.300 ;
        RECT 521.660 4.000 528.340 4.300 ;
        RECT 529.500 4.000 536.180 4.300 ;
        RECT 537.340 4.000 544.020 4.300 ;
        RECT 545.180 4.000 551.860 4.300 ;
        RECT 553.020 4.000 559.700 4.300 ;
        RECT 560.860 4.000 567.540 4.300 ;
        RECT 568.700 4.000 575.380 4.300 ;
        RECT 576.540 4.000 583.220 4.300 ;
        RECT 584.380 4.000 591.060 4.300 ;
        RECT 592.220 4.000 598.900 4.300 ;
        RECT 600.060 4.000 606.740 4.300 ;
        RECT 607.900 4.000 614.580 4.300 ;
        RECT 615.740 4.000 622.420 4.300 ;
        RECT 623.580 4.000 630.260 4.300 ;
        RECT 631.420 4.000 638.100 4.300 ;
        RECT 639.260 4.000 645.940 4.300 ;
        RECT 647.100 4.000 653.780 4.300 ;
        RECT 654.940 4.000 661.620 4.300 ;
        RECT 662.780 4.000 669.460 4.300 ;
        RECT 670.620 4.000 677.300 4.300 ;
        RECT 678.460 4.000 685.140 4.300 ;
        RECT 686.300 4.000 692.980 4.300 ;
        RECT 694.140 4.000 700.820 4.300 ;
        RECT 701.980 4.000 708.660 4.300 ;
        RECT 709.820 4.000 716.500 4.300 ;
        RECT 717.660 4.000 724.340 4.300 ;
        RECT 725.500 4.000 732.180 4.300 ;
        RECT 733.340 4.000 740.020 4.300 ;
        RECT 741.180 4.000 747.860 4.300 ;
        RECT 749.020 4.000 755.700 4.300 ;
        RECT 756.860 4.000 763.540 4.300 ;
        RECT 764.700 4.000 771.380 4.300 ;
        RECT 772.540 4.000 779.220 4.300 ;
        RECT 780.380 4.000 787.060 4.300 ;
        RECT 788.220 4.000 794.900 4.300 ;
        RECT 796.060 4.000 797.300 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 788.220 797.350 792.260 ;
        RECT 4.300 787.060 797.350 788.220 ;
        RECT 0.090 769.740 797.350 787.060 ;
        RECT 4.300 768.580 797.350 769.740 ;
        RECT 0.090 751.260 797.350 768.580 ;
        RECT 4.300 750.100 797.350 751.260 ;
        RECT 0.090 732.780 797.350 750.100 ;
        RECT 4.300 731.620 797.350 732.780 ;
        RECT 0.090 714.300 797.350 731.620 ;
        RECT 4.300 713.140 797.350 714.300 ;
        RECT 0.090 695.820 797.350 713.140 ;
        RECT 4.300 694.660 797.350 695.820 ;
        RECT 0.090 677.340 797.350 694.660 ;
        RECT 4.300 676.180 797.350 677.340 ;
        RECT 0.090 658.860 797.350 676.180 ;
        RECT 4.300 657.700 797.350 658.860 ;
        RECT 0.090 640.380 797.350 657.700 ;
        RECT 4.300 639.220 797.350 640.380 ;
        RECT 0.090 621.900 797.350 639.220 ;
        RECT 4.300 620.740 797.350 621.900 ;
        RECT 0.090 603.420 797.350 620.740 ;
        RECT 4.300 602.260 797.350 603.420 ;
        RECT 0.090 584.940 797.350 602.260 ;
        RECT 4.300 583.780 797.350 584.940 ;
        RECT 0.090 566.460 797.350 583.780 ;
        RECT 4.300 565.300 797.350 566.460 ;
        RECT 0.090 547.980 797.350 565.300 ;
        RECT 4.300 546.820 797.350 547.980 ;
        RECT 0.090 529.500 797.350 546.820 ;
        RECT 4.300 528.340 797.350 529.500 ;
        RECT 0.090 511.020 797.350 528.340 ;
        RECT 4.300 509.860 797.350 511.020 ;
        RECT 0.090 492.540 797.350 509.860 ;
        RECT 4.300 491.380 797.350 492.540 ;
        RECT 0.090 474.060 797.350 491.380 ;
        RECT 4.300 472.900 797.350 474.060 ;
        RECT 0.090 455.580 797.350 472.900 ;
        RECT 4.300 454.420 797.350 455.580 ;
        RECT 0.090 437.100 797.350 454.420 ;
        RECT 4.300 435.940 797.350 437.100 ;
        RECT 0.090 418.620 797.350 435.940 ;
        RECT 4.300 417.460 797.350 418.620 ;
        RECT 0.090 400.140 797.350 417.460 ;
        RECT 4.300 398.980 797.350 400.140 ;
        RECT 0.090 381.660 797.350 398.980 ;
        RECT 4.300 380.500 797.350 381.660 ;
        RECT 0.090 363.180 797.350 380.500 ;
        RECT 4.300 362.020 797.350 363.180 ;
        RECT 0.090 344.700 797.350 362.020 ;
        RECT 4.300 343.540 797.350 344.700 ;
        RECT 0.090 326.220 797.350 343.540 ;
        RECT 4.300 325.060 797.350 326.220 ;
        RECT 0.090 307.740 797.350 325.060 ;
        RECT 4.300 306.580 797.350 307.740 ;
        RECT 0.090 289.260 797.350 306.580 ;
        RECT 4.300 288.100 797.350 289.260 ;
        RECT 0.090 270.780 797.350 288.100 ;
        RECT 4.300 269.620 797.350 270.780 ;
        RECT 0.090 252.300 797.350 269.620 ;
        RECT 4.300 251.140 797.350 252.300 ;
        RECT 0.090 233.820 797.350 251.140 ;
        RECT 4.300 232.660 797.350 233.820 ;
        RECT 0.090 215.340 797.350 232.660 ;
        RECT 4.300 214.180 797.350 215.340 ;
        RECT 0.090 196.860 797.350 214.180 ;
        RECT 4.300 195.700 797.350 196.860 ;
        RECT 0.090 178.380 797.350 195.700 ;
        RECT 4.300 177.220 797.350 178.380 ;
        RECT 0.090 159.900 797.350 177.220 ;
        RECT 4.300 158.740 797.350 159.900 ;
        RECT 0.090 141.420 797.350 158.740 ;
        RECT 4.300 140.260 797.350 141.420 ;
        RECT 0.090 122.940 797.350 140.260 ;
        RECT 4.300 121.780 797.350 122.940 ;
        RECT 0.090 104.460 797.350 121.780 ;
        RECT 4.300 103.300 797.350 104.460 ;
        RECT 0.090 85.980 797.350 103.300 ;
        RECT 4.300 84.820 797.350 85.980 ;
        RECT 0.090 67.500 797.350 84.820 ;
        RECT 4.300 66.340 797.350 67.500 ;
        RECT 0.090 49.020 797.350 66.340 ;
        RECT 4.300 47.860 797.350 49.020 ;
        RECT 0.090 30.540 797.350 47.860 ;
        RECT 4.300 29.380 797.350 30.540 ;
        RECT 0.090 12.060 797.350 29.380 ;
        RECT 4.300 10.900 797.350 12.060 ;
        RECT 0.090 4.620 797.350 10.900 ;
      LAYER Metal4 ;
        RECT 4.620 15.080 21.940 774.950 ;
        RECT 24.140 15.080 98.740 774.950 ;
        RECT 100.940 15.080 175.540 774.950 ;
        RECT 177.740 15.080 252.340 774.950 ;
        RECT 254.540 15.080 329.140 774.950 ;
        RECT 331.340 15.080 405.940 774.950 ;
        RECT 408.140 15.080 482.740 774.950 ;
        RECT 484.940 15.080 559.540 774.950 ;
        RECT 561.740 15.080 636.340 774.950 ;
        RECT 638.540 15.080 713.140 774.950 ;
        RECT 715.340 15.080 779.380 774.950 ;
        RECT 4.620 5.690 779.380 15.080 ;
  END
END wfg_top
END LIBRARY

