* NGSPICE file created from wb_memory.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

.subckt wb_memory addr_mem0[0] addr_mem0[1] addr_mem0[2] addr_mem0[3] addr_mem0[4]
+ addr_mem0[5] addr_mem0[6] addr_mem0[7] addr_mem0[8] addr_mem1[0] addr_mem1[1] addr_mem1[2]
+ addr_mem1[3] addr_mem1[4] addr_mem1[5] addr_mem1[6] addr_mem1[7] addr_mem1[8] csb_mem0
+ csb_mem1 din_mem0[0] din_mem0[10] din_mem0[11] din_mem0[12] din_mem0[13] din_mem0[14]
+ din_mem0[15] din_mem0[16] din_mem0[17] din_mem0[18] din_mem0[19] din_mem0[1] din_mem0[20]
+ din_mem0[21] din_mem0[22] din_mem0[23] din_mem0[24] din_mem0[25] din_mem0[26] din_mem0[27]
+ din_mem0[28] din_mem0[29] din_mem0[2] din_mem0[30] din_mem0[31] din_mem0[3] din_mem0[4]
+ din_mem0[5] din_mem0[6] din_mem0[7] din_mem0[8] din_mem0[9] din_mem1[0] din_mem1[10]
+ din_mem1[11] din_mem1[12] din_mem1[13] din_mem1[14] din_mem1[15] din_mem1[16] din_mem1[17]
+ din_mem1[18] din_mem1[19] din_mem1[1] din_mem1[20] din_mem1[21] din_mem1[22] din_mem1[23]
+ din_mem1[24] din_mem1[25] din_mem1[26] din_mem1[27] din_mem1[28] din_mem1[29] din_mem1[2]
+ din_mem1[30] din_mem1[31] din_mem1[3] din_mem1[4] din_mem1[5] din_mem1[6] din_mem1[7]
+ din_mem1[8] din_mem1[9] dout_mem0[0] dout_mem0[10] dout_mem0[11] dout_mem0[12] dout_mem0[13]
+ dout_mem0[14] dout_mem0[15] dout_mem0[16] dout_mem0[17] dout_mem0[18] dout_mem0[19]
+ dout_mem0[1] dout_mem0[20] dout_mem0[21] dout_mem0[22] dout_mem0[23] dout_mem0[24]
+ dout_mem0[25] dout_mem0[26] dout_mem0[27] dout_mem0[28] dout_mem0[29] dout_mem0[2]
+ dout_mem0[30] dout_mem0[31] dout_mem0[3] dout_mem0[4] dout_mem0[5] dout_mem0[6]
+ dout_mem0[7] dout_mem0[8] dout_mem0[9] dout_mem1[0] dout_mem1[10] dout_mem1[11]
+ dout_mem1[12] dout_mem1[13] dout_mem1[14] dout_mem1[15] dout_mem1[16] dout_mem1[17]
+ dout_mem1[18] dout_mem1[19] dout_mem1[1] dout_mem1[20] dout_mem1[21] dout_mem1[22]
+ dout_mem1[23] dout_mem1[24] dout_mem1[25] dout_mem1[26] dout_mem1[27] dout_mem1[28]
+ dout_mem1[29] dout_mem1[2] dout_mem1[30] dout_mem1[31] dout_mem1[3] dout_mem1[4]
+ dout_mem1[5] dout_mem1[6] dout_mem1[7] dout_mem1[8] dout_mem1[9] io_wbs_ack io_wbs_adr[0]
+ io_wbs_adr[10] io_wbs_adr[11] io_wbs_adr[12] io_wbs_adr[13] io_wbs_adr[14] io_wbs_adr[15]
+ io_wbs_adr[16] io_wbs_adr[17] io_wbs_adr[18] io_wbs_adr[19] io_wbs_adr[1] io_wbs_adr[20]
+ io_wbs_adr[21] io_wbs_adr[22] io_wbs_adr[23] io_wbs_adr[24] io_wbs_adr[25] io_wbs_adr[26]
+ io_wbs_adr[27] io_wbs_adr[28] io_wbs_adr[29] io_wbs_adr[2] io_wbs_adr[30] io_wbs_adr[31]
+ io_wbs_adr[3] io_wbs_adr[4] io_wbs_adr[5] io_wbs_adr[6] io_wbs_adr[7] io_wbs_adr[8]
+ io_wbs_adr[9] io_wbs_clk io_wbs_cyc io_wbs_datrd[0] io_wbs_datrd[10] io_wbs_datrd[11]
+ io_wbs_datrd[12] io_wbs_datrd[13] io_wbs_datrd[14] io_wbs_datrd[15] io_wbs_datrd[16]
+ io_wbs_datrd[17] io_wbs_datrd[18] io_wbs_datrd[19] io_wbs_datrd[1] io_wbs_datrd[20]
+ io_wbs_datrd[21] io_wbs_datrd[22] io_wbs_datrd[23] io_wbs_datrd[24] io_wbs_datrd[25]
+ io_wbs_datrd[26] io_wbs_datrd[27] io_wbs_datrd[28] io_wbs_datrd[29] io_wbs_datrd[2]
+ io_wbs_datrd[30] io_wbs_datrd[31] io_wbs_datrd[3] io_wbs_datrd[4] io_wbs_datrd[5]
+ io_wbs_datrd[6] io_wbs_datrd[7] io_wbs_datrd[8] io_wbs_datrd[9] io_wbs_datwr[0]
+ io_wbs_datwr[10] io_wbs_datwr[11] io_wbs_datwr[12] io_wbs_datwr[13] io_wbs_datwr[14]
+ io_wbs_datwr[15] io_wbs_datwr[16] io_wbs_datwr[17] io_wbs_datwr[18] io_wbs_datwr[19]
+ io_wbs_datwr[1] io_wbs_datwr[20] io_wbs_datwr[21] io_wbs_datwr[22] io_wbs_datwr[23]
+ io_wbs_datwr[24] io_wbs_datwr[25] io_wbs_datwr[26] io_wbs_datwr[27] io_wbs_datwr[28]
+ io_wbs_datwr[29] io_wbs_datwr[2] io_wbs_datwr[30] io_wbs_datwr[31] io_wbs_datwr[3]
+ io_wbs_datwr[4] io_wbs_datwr[5] io_wbs_datwr[6] io_wbs_datwr[7] io_wbs_datwr[8]
+ io_wbs_datwr[9] io_wbs_rst io_wbs_sel[0] io_wbs_sel[1] io_wbs_sel[2] io_wbs_sel[3]
+ io_wbs_stb io_wbs_we vdd vss web_mem0 web_mem1 wmask_mem0[0] wmask_mem0[1] wmask_mem0[2]
+ wmask_mem0[3] wmask_mem1[0] wmask_mem1[1] wmask_mem1[2] wmask_mem1[3]
XFILLER_39_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__189__I1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input108_I io_wbs_rst vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input73_I io_wbs_adr[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__190__S _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_432_ net105 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__429__I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_294_ _158_ _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_363_ _062_ _027_ clknet_2_3__leaf_io_wbs_clk net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_3_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__275__S _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__185__S _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_415_ net90 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_346_ _045_ _010_ clknet_2_0__leaf_io_wbs_clk net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_277_ _148_ _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_0_io_wbs_clk_I io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwb_memory_240 csb_mem0 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__261__I0 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput231 net231 web_mem1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput220 net220 io_wbs_datrd[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input36_I dout_mem1[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_200_ _071_ _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__252__I0 net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__442__I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__243__I0 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_329_ _166_ _029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__234__I0 net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__351__CLK clknet_2_2__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__437__I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__193__S _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__278__S _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__450__I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input66_I io_wbs_adr[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output222_I net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_431_ net104 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__445__I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_362_ _061_ _026_ clknet_2_2__leaf_io_wbs_clk net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_293_ _157_ _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_414_ net89 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_345_ _044_ _009_ clknet_2_0__leaf_io_wbs_clk net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_276_ net220 _147_ _145_ _148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__261__I1 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwb_memory_241 csb_mem1 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput232 net232 wmask_mem0[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput221 net221 io_wbs_datrd[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput210 net210 io_wbs_datrd[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input29_I dout_mem0[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__196__S _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__252__I1 _130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__243__I1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_328_ _166_ _028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_259_ net227 _134_ _135_ _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__234__I1 _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__453__I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input96_I io_wbs_datwr[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__448__I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__341__CLK clknet_2_0__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input11_I dout_mem0[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput110 io_wbs_sel[1] net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__178__I _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__364__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I dout_mem0[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input59_I dout_mem1[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__199__S _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_430_ net103 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_292_ net108 _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_361_ _060_ _025_ clknet_2_3__leaf_io_wbs_clk net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_42_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__461__I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input113_I io_wbs_stb vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output165_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_413_ net88 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__456__I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_275_ net23 net55 _139_ _147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_344_ _043_ _008_ clknet_2_1__leaf_io_wbs_clk net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput200 net200 io_wbs_datrd[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput233 net233 wmask_mem0[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput222 net222 io_wbs_datrd[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput211 net211 io_wbs_datrd[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_4_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__186__I _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_189_ net19 net51 _077_ _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_327_ _166_ _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_258_ _104_ _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input41_I dout_mem1[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output128_I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input89_I io_wbs_datwr[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__464__I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output195_I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput111 io_wbs_sel[2] net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput100 io_wbs_datwr[31] net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__459__I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output208_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_291_ _156_ net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_360_ _059_ _024_ clknet_2_2__leaf_io_wbs_clk net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input106_I io_wbs_datwr[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input71_I io_wbs_adr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__354__CLK clknet_2_2__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_412_ net86 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__255__I0 net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_343_ _042_ _007_ clknet_2_1__leaf_io_wbs_clk net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_274_ _146_ _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput234 net234 wmask_mem0[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__382__I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput223 net223 io_wbs_datrd[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput201 net201 io_wbs_datrd[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput212 net212 io_wbs_datrd[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__237__I0 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__292__I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_326_ _166_ _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_257_ net30 net62 _129_ _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_188_ _084_ _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__377__I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__219__I0 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input34_I dout_mem1[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_309_ _162_ _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output140_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output238_I net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__390__I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput112 io_wbs_sel[3] net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput101 io_wbs_datwr[3] net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__385__I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__295__I _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__282__I1 _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_290_ web_mem _069_ _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__273__I1 _144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input64_I dout_mem1[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_411_ net85 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__255__I1 _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_342_ _041_ _006_ clknet_2_0__leaf_io_wbs_clk net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_2_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_273_ net223 _144_ _145_ _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__182__I0 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput235 net235 wmask_mem0[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput202 net202 io_wbs_datrd[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput224 net224 io_wbs_datrd[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput213 net213 io_wbs_datrd[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__237__I1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_325_ _157_ _166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_187_ net217 _082_ _083_ _084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_256_ _133_ _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__393__I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__344__CLK clknet_2_1__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input27_I dout_mem0[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__367__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_308_ _162_ _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_239_ _121_ _050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__388__I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__298__I _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input94_I io_wbs_datwr[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput102 io_wbs_datwr[4] net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput113 io_wbs_stb net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_3__f_io_wbs_clk_I clknet_0_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input1_I dout_mem0[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__396__I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input57_I dout_mem1[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output213_I net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_410_ net84 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_341_ _040_ _005_ clknet_2_0__leaf_io_wbs_clk net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_272_ operation _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput236 net236 wmask_mem1[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput203 net203 io_wbs_datrd[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput225 net225 io_wbs_datrd[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput214 net214 io_wbs_datrd[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input111_I io_wbs_sel[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output163_I net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_255_ net228 _132_ _125_ _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_324_ _165_ _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_186_ _071_ _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_169_ net25 net57 _069_ _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_238_ net202 _120_ _115_ _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_307_ _162_ _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output126_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__399__I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input87_I io_wbs_datwr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__357__CLK clknet_2_2__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput103 io_wbs_datwr[5] net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput114 io_wbs_we net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_5_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output193_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__208__S _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output206_I net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_271_ net26 net58 _139_ _144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_340_ _039_ _004_ clknet_2_1__leaf_io_wbs_clk net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput237 net237 wmask_mem1[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput215 net215 io_wbs_datrd[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput226 net226 io_wbs_datrd[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput204 net204 io_wbs_datrd[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__200__I _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input104_I io_wbs_datwr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_185_ net20 net52 _077_ _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_254_ net31 net63 _129_ _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_323_ _165_ _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_306_ _162_ _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_237_ net5 net37 _119_ _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_168_ net66 _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__289__A1 _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input32_I dout_mem0[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output119_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput104 io_wbs_datwr[6] net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_output236_I net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__276__I1 _147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__224__S _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__347__CLK clknet_2_0__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__185__I0 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_270_ _143_ _041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__219__S _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_399_ net104 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput205 net205 io_wbs_datrd[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput216 net216 io_wbs_datrd[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput238 net238 wmask_mem1[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput227 net227 io_wbs_datrd[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_4_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input62_I dout_mem1[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output149_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_322_ _165_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_253_ _131_ _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_184_ _081_ _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__301__I _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_305_ _160_ _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_236_ _097_ _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__206__I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__289__A2 _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input25_I dout_mem0[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_219_ net10 net42 _098_ _107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__227__S _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput105 io_wbs_datwr[7] net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output131_I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output229_I net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input92_I io_wbs_datwr[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__194__I1 _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__240__S _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__304__I _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__185__I1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_398_ net103 net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput239 net239 wmask_mem1[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput206 net206 io_wbs_datrd[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xclkbuf_2_2__f_io_wbs_clk clknet_0_io_wbs_clk clknet_2_2__leaf_io_wbs_clk vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xoutput228 net228 io_wbs_datrd[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput217 net217 io_wbs_datrd[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input55_I dout_mem1[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output211_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_321_ _165_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_252_ net229 _130_ _125_ _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_183_ net218 _080_ _072_ _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__402__I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_304_ _161_ _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_235_ _118_ _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__312__I _163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__222__I _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input18_I dout_mem0[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__243__S _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__212__I0 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__307__I _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_218_ _106_ _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__203__I0 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput106 io_wbs_datwr[8] net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_5_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output124_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__238__S _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__359__D _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input85_I io_wbs_datwr[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__410__I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__370__CLK clknet_2_1__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__320__I _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__230__I _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output191_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__405__I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_397_ net102 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__251__S _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput207 net207 io_wbs_datrd[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput229 net229 io_wbs_datrd[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput218 net218 io_wbs_datrd[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__315__I _160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input48_I dout_mem1[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output204_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_182_ net21 net53 _077_ _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_251_ net32 net64 _129_ _130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_320_ _157_ _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_449_ net92 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__367__D _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input102_I io_wbs_datwr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output154_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_303_ _161_ _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_234_ net203 _117_ _115_ _118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__413__I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__212__I1 _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_217_ net208 _103_ _105_ _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__279__I1 _149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__203__I1 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input30_I dout_mem0[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput107 io_wbs_datwr[9] net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_5_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__408__I net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__254__S _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__318__I _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__197__I0 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input78_I io_wbs_datwr[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__179__I0 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__421__I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_396_ net101 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput208 net208 io_wbs_datrd[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput219 net219 io_wbs_datrd[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_36_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__360__CLK clknet_2_2__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_250_ _097_ _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__416__I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_181_ _079_ _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_448_ net91 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_379_ net71 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__262__S _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__236__I _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input60_I dout_mem1[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__172__S _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output147_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_302_ _161_ _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_233_ net6 net38 _109_ _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__257__S _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_216_ _104_ _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput108 io_wbs_rst net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_0_io_wbs_clk io_wbs_clk clknet_0_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input23_I dout_mem0[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__424__I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__197__I1 _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput90 io_wbs_datwr[22] net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__180__S _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__244__I _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__419__I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__265__S _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input90_I io_wbs_datwr[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__175__S _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output177_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_464_ net112 net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_395_ net98 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput209 net209 io_wbs_datrd[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__251__I0 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_180_ net219 _078_ _072_ _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__432__I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_447_ net90 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_378_ net70 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__233__I0 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input53_I dout_mem1[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__427__I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_301_ _161_ _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_232_ _116_ _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__224__I0 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__337__I _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__350__CLK clknet_2_2__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__273__S _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__183__S _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_215_ operation _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__268__S _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput109 io_wbs_sel[0] net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input16_I dout_mem0[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__440__I net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I dout_mem0[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput80 io_wbs_datwr[13] net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput91 io_wbs_datwr[23] net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output122_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__435__I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__170__I operation vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__281__S _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input83_I io_wbs_datwr[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_463_ net111 net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_394_ net87 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__276__S _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__251__I1 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_377_ net69 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_446_ net89 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__233__I1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input46_I dout_mem1[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_300_ _160_ _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_231_ net204 _114_ _115_ _116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__224__I1 _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__443__I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_429_ net102 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 dout_mem0[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input100_I io_wbs_datwr[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output152_I net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__438__I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_214_ net11 net43 _098_ _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__258__I _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__194__S _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__340__CLK clknet_2_1__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput190 net190 din_mem1[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__168__I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__279__S _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__363__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput81 io_wbs_datwr[14] net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput70 io_wbs_adr[5] net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput92 io_wbs_datwr[24] net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__189__S _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__451__I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input76_I io_wbs_datwr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_393_ net76 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_462_ net110 net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__446__I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_445_ net88 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_376_ net68 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input39_I dout_mem1[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__197__S _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_230_ _104_ _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_428_ net101 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_359_ _058_ _023_ clknet_2_3__leaf_io_wbs_clk net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput2 dout_mem0[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__454__I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_213_ _102_ _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput191 net191 din_mem1[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput180 net180 din_mem1[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__449__I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput60 dout_mem1[5] net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput82 io_wbs_datwr[15] net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput71 io_wbs_adr[6] net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput93 io_wbs_datwr[25] net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input21_I dout_mem0[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__281__I0 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input69_I io_wbs_adr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__254__I0 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_461_ net109 net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_392_ net65 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__462__I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__353__CLK clknet_2_2__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output175_I net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_444_ net86 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__457__I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__227__I0 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_375_ net67 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__192__I _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__209__I0 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_427_ net98 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_358_ _057_ _022_ clknet_2_3__leaf_io_wbs_clk net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_289_ _155_ _069_ net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 dout_mem0[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input51_I dout_mem1[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output138_I net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_212_ net210 _101_ _093_ _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__380__I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input99_I io_wbs_datwr[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput181 net181 din_mem1[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput170 net170 din_mem1[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput192 net192 din_mem1[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__375__I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput50 dout_mem1[25] net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput61 dout_mem1[6] net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput72 io_wbs_adr[7] net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput83 io_wbs_datwr[16] net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput94 io_wbs_datwr[26] net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input14_I dout_mem0[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__281__I1 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I dout_mem0[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_460_ net112 net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_391_ net74 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output120_I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__254__I1 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output218_I net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__245__I1 _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input81_I io_wbs_datwr[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__172__I0 net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_443_ net85 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__227__I1 _112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__383__I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__293__I _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__209__I1 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__343__CLK clknet_2_1__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_426_ net87 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_357_ _056_ _021_ clknet_2_2__leaf_io_wbs_clk net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_288_ web_mem _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__378__I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 dout_mem0[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__366__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input44_I dout_mem1[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__288__I web_mem vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_211_ net13 net45 _098_ _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_409_ net83 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput182 net182 din_mem1[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput160 net160 din_mem0[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput193 net193 din_mem1[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput171 net171 din_mem1[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output150_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput40 dout_mem1[16] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput51 dout_mem1[26] net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput62 dout_mem1[7] net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__391__I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput84 io_wbs_datwr[17] net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput73 io_wbs_adr[8] net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput95 io_wbs_datwr[27] net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__386__I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_390_ net73 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__296__I _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__190__I1 _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input109_I io_wbs_sel[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input74_I io_wbs_adr[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__172__I1 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output230_I net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_442_ net84 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_425_ net76 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_287_ net113 net75 net114 _153_ _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_356_ _055_ _020_ clknet_2_3__leaf_io_wbs_clk net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput5 dout_mem0[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__394__I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input37_I dout_mem1[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_210_ _100_ _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_408_ net82 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_339_ _038_ _003_ clknet_2_1__leaf_io_wbs_clk net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__389__I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput161 net161 din_mem0[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput150 net150 din_mem0[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput183 net183 din_mem1[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput172 net172 din_mem1[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput194 net194 din_mem1[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output143_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__299__I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__203__S _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__356__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__275__I0 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput52 dout_mem1[27] net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput63 dout_mem1[8] net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput30 dout_mem0[7] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput41 dout_mem1[17] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput85 io_wbs_datwr[18] net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput74 io_wbs_adr[9] net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput96 io_wbs_datwr[28] net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__257__I0 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__248__I0 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__397__I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input67_I io_wbs_adr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_441_ net83 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_372_ _000_ _036_ clknet_2_1__leaf_io_wbs_clk operation vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__211__S _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_424_ net100 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_355_ _054_ _019_ clknet_2_3__leaf_io_wbs_clk net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_286_ _154_ _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 dout_mem0[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_407_ net81 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_338_ _037_ _002_ clknet_2_1__leaf_io_wbs_clk net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_269_ net224 _142_ _135_ _143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput173 net173 din_mem1[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput195 net195 din_mem1[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput140 net140 din_mem0[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput162 net162 din_mem0[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput184 net184 din_mem1[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput151 net151 din_mem0[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output136_I net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__275__I1 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput20 dout_mem0[27] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput31 dout_mem0[8] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput42 dout_mem1[18] net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput53 dout_mem1[28] net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput64 dout_mem1[9] net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput86 io_wbs_datwr[19] net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput75 io_wbs_cyc net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput97 io_wbs_datwr[29] net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_38_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__266__I1 _140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input97_I io_wbs_datwr[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__257__I1 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__214__S _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__193__I0 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__248__I1 _127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I dout_mem0[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__346__CLK clknet_2_0__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__175__I0 net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I dout_mem0[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__369__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_440_ net82 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_371_ _001_ _035_ clknet_2_1__leaf_io_wbs_clk web_mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input114_I io_wbs_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output166_I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_423_ net99 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_354_ _053_ _018_ clknet_2_2__leaf_io_wbs_clk net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_41_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_285_ net113 net75 _153_ _154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput7 dout_mem0[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_406_ net80 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_337_ _158_ _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__217__S _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_268_ net27 net59 _139_ _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_199_ net16 net48 _087_ _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input42_I dout_mem1[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput163 net163 din_mem0[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput185 net185 din_mem1[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput174 net174 din_mem1[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput196 net196 din_mem1[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput130 net130 addr_mem1[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput152 net152 din_mem0[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput141 net141 din_mem0[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output129_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput54 dout_mem1[29] net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput21 dout_mem0[28] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput10 dout_mem0[18] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput32 dout_mem0[9] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput43 dout_mem1[19] net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput65 io_wbs_adr[10] net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput76 io_wbs_datwr[0] net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput87 io_wbs_datwr[1] net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput98 io_wbs_datwr[2] net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__193__I1 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output196_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__175__I1 _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_370_ operation _034_ clknet_2_1__leaf_io_wbs_clk net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_5_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input107_I io_wbs_datwr[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input72_I io_wbs_adr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output159_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_422_ net97 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_284_ _071_ net197 _153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_353_ _052_ _017_ clknet_2_2__leaf_io_wbs_clk net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__359__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 dout_mem0[16] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_39_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__302__I _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__220__I0 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__211__I0 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_405_ net79 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_336_ _158_ _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_267_ _141_ _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__233__S _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_198_ _091_ _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__207__I _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput186 net186 din_mem1[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput142 net142 din_mem0[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput164 net164 din_mem0[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput120 net120 addr_mem0[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput175 net175 din_mem1[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input35_I dout_mem1[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput131 net131 addr_mem1[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput153 net153 din_mem0[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput197 net197 io_wbs_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput55 dout_mem1[2] net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput33 dout_mem1[0] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput44 dout_mem1[1] net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput22 dout_mem0[29] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput11 dout_mem0[19] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput88 io_wbs_datwr[20] net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput66 io_wbs_adr[11] net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_319_ _164_ _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput77 io_wbs_datwr[10] net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput99 io_wbs_datwr[30] net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output239_I net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__400__I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__310__I _160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__305__I _160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__241__S _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__215__I operation vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_2_0__f_io_wbs_clk_I clknet_0_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input65_I io_wbs_adr[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_421_ net96 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output221_I net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_352_ _051_ _016_ clknet_2_3__leaf_io_wbs_clk net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_283_ _152_ _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput9 dout_mem0[17] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__403__I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__220__I1 _107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_404_ net78 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_335_ _158_ _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_266_ net225 _140_ _135_ _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_197_ net214 _090_ _083_ _091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__313__I _163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__278__I1 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput132 net132 addr_mem1[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput121 net121 addr_mem0[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput143 net143 din_mem0[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__370__D operation vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput187 net187 din_mem1[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput165 net165 din_mem1[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput154 net154 din_mem0[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput176 net176 din_mem1[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input28_I dout_mem0[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput198 net198 io_wbs_datrd[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__269__I1 _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__349__CLK clknet_2_1__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__308__I _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput34 dout_mem1[10] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput23 dout_mem0[2] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput12 dout_mem0[1] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput45 dout_mem1[20] net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput56 dout_mem1[30] net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__196__I0 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput89 io_wbs_datwr[21] net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput78 io_wbs_datwr[11] net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput67 io_wbs_adr[2] net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_318_ _164_ _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_249_ _128_ _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__187__I0 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output134_I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__169__I0 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input95_I io_wbs_datwr[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__411__I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input10_I dout_mem0[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__406__I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__316__I _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I dout_mem0[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input58_I dout_mem1[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_2_1__f_io_wbs_clk clknet_0_io_wbs_clk clknet_2_1__leaf_io_wbs_clk vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_420_ net95 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output214_I net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_351_ _050_ _015_ clknet_2_2__leaf_io_wbs_clk net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_2_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_282_ net198 _151_ _145_ _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__247__S _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input112_I io_wbs_sel[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output164_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_403_ net77 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_334_ _167_ _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_196_ net17 net49 _087_ _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_265_ net28 net60 _139_ _140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput155 net155 din_mem0[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput144 net144 din_mem0[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput177 net177 din_mem1[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput122 net122 addr_mem0[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput133 net133 din_mem0[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput166 net166 din_mem1[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput188 net188 din_mem1[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput199 net199 io_wbs_datrd[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__414__I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput13 dout_mem0[20] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_317_ _164_ _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput46 dout_mem1[21] net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput57 dout_mem1[31] net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput35 dout_mem1[11] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput24 dout_mem0[30] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_179_ net22 net54 _077_ _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__196__I1 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput79 io_wbs_datwr[12] net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput68 io_wbs_adr[3] net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_248_ net199 _127_ _125_ _128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__187__I1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input40_I dout_mem1[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output127_I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__409__I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__319__I _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__169__I1 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__339__CLK clknet_2_1__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input88_I io_wbs_datwr[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__422__I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__417__I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output207_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_350_ _049_ _014_ clknet_2_2__leaf_io_wbs_clk net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_41_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_281_ net1 net33 _076_ _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__223__I0 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__214__I0 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input105_I io_wbs_datwr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input70_I io_wbs_adr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_264_ net66 _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_402_ net107 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_333_ _167_ _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_195_ _089_ _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__372__CLK clknet_2_1__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput178 net178 din_mem1[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput167 net167 din_mem1[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput156 net156 din_mem0[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput145 net145 din_mem0[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput134 net134 din_mem0[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput189 net189 din_mem1[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput123 net123 addr_mem0[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__430__I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__290__A1 web_mem vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput36 dout_mem1[12] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput25 dout_mem0[31] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput14 dout_mem0[21] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_247_ net2 net34 _119_ _127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_316_ _164_ _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_178_ _076_ _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput58 dout_mem1[3] net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput47 dout_mem1[22] net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput69 io_wbs_adr[4] net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input33_I dout_mem1[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__250__I _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__425__I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__271__S _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__335__I _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output237_I net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__266__S _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output187_I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__241__I1 _122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__223__I1 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_280_ _150_ _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__433__I net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input63_I dout_mem1[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__428__I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_401_ net106 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_263_ _138_ _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_332_ _167_ _031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_194_ net215 _088_ _083_ _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__199__I0 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput124 net124 addr_mem1[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput146 net146 din_mem0[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput168 net168 din_mem1[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput157 net157 din_mem0[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput135 net135 din_mem0[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput179 net179 din_mem1[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_3_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__290__A2 _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput48 dout_mem1[23] net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput59 dout_mem1[4] net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput15 dout_mem0[22] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput26 dout_mem0[3] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput37 dout_mem1[13] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_177_ net66 _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_315_ _160_ _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_246_ _126_ _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__269__S _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__179__S _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input26_I dout_mem0[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__362__CLK clknet_2_2__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__441__I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_229_ net7 net39 _109_ _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output132_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__436__I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__171__I _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__282__S _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input93_I io_wbs_datwr[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__187__S _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input56_I dout_mem1[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_400_ net105 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output212_I net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_331_ _167_ _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_193_ net18 net50 _087_ _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__444__I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_262_ net226 _137_ _135_ _138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput125 net125 addr_mem1[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput158 net158 din_mem0[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput147 net147 din_mem0[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput136 net136 din_mem0[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput169 net169 din_mem1[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input110_I io_wbs_sel[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__264__I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output162_I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__439__I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_314_ _163_ _017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput38 dout_mem1[14] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput27 dout_mem0[4] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput49 dout_mem1[24] net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput16 dout_mem0[23] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_245_ net200 _124_ _125_ _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_176_ _075_ _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input19_I dout_mem0[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__271__I0 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_228_ _113_ _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output125_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__452__I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__352__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input86_I io_wbs_datwr[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__272__I operation vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__447__I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__226__I0 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__217__I0 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__208__I0 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output192_I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__177__I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__358__RN _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I dout_mem1[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output205_I net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_330_ _157_ _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_192_ _076_ _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_261_ net29 net61 _129_ _137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__460__I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_459_ net111 net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput159 net159 din_mem0[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput115 net115 addr_mem0[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput126 net126 addr_mem1[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput148 net148 din_mem0[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput137 net137 din_mem0[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__284__A1 _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input103_I io_wbs_datwr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__455__I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_313_ _163_ _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_244_ _104_ _125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput17 dout_mem0[24] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput28 dout_mem0[5] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput39 dout_mem1[15] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_175_ net221 _074_ _072_ _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__271__I1 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_227_ net205 _112_ _105_ _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__262__I1 _137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input31_I dout_mem0[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__180__I0 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input79_I io_wbs_datwr[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__226__I1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__463__I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__217__I1 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__458__I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__342__CLK clknet_2_0__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__365__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_260_ _136_ _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_191_ _086_ _063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_389_ net72 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_458_ net110 net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput138 net138 din_mem0[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput116 net116 addr_mem0[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput149 net149 din_mem0[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput127 net127 addr_mem1[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__284__A2 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input61_I dout_mem1[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output148_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput18 dout_mem0[25] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_243_ net3 net35 _119_ _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_312_ _163_ _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput29 dout_mem0[6] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_174_ net24 net56 _069_ _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__381__I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_226_ net8 net40 _109_ _112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__376__I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input24_I dout_mem0[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_2_1__f_io_wbs_clk_I clknet_0_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_209_ net211 _099_ _093_ _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__180__I1 _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output130_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output228_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input91_I io_wbs_datwr[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output178_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__384__I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__294__I _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_190_ net216 _085_ _083_ _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_388_ net71 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_457_ net109 net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput128 net128 addr_mem1[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput117 net117 addr_mem0[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput139 net139 din_mem0[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__379__I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input54_I dout_mem1[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output210_I net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput19 dout_mem0[26] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_173_ _073_ _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_311_ _163_ _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_242_ _123_ _049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__355__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__265__I0 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output160_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_225_ _111_ _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__247__I0 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__392__I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input17_I dout_mem0[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__229__I0 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_208_ net14 net46 _098_ _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__387__I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I dout_mem0[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output123_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__297__I _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input84_I io_wbs_datwr[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output190_I net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_456_ net100 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_387_ net70 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput129 net129 addr_mem1[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput118 net118 addr_mem0[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__395__I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input47_I dout_mem1[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_310_ _160_ _163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output203_I net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_172_ net222 _070_ _072_ _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_241_ net201 _122_ _115_ _123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_439_ net81 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__265__I1 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input101_I io_wbs_datwr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output153_I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_224_ net206 _110_ _105_ _111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__247__I1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__183__I0 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__238__I1 _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__174__I0 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__229__I1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_207_ _097_ _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__345__CLK clknet_2_0__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__368__CLK clknet_2_2__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__398__I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input77_I io_wbs_datwr[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_455_ net99 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_386_ net69 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput119 net119 addr_mem0[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_240_ net4 net36 _119_ _122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_171_ _071_ _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_438_ net80 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_369_ _068_ _033_ clknet_2_3__leaf_io_wbs_clk net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output146_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_223_ net9 net41 _109_ _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__220__S _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__183__I1 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__174__I1 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_206_ net66 _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input22_I dout_mem0[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__358__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output176_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_454_ net97 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_385_ net68 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__223__S _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__201__I0 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__268__I0 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_3__f_io_wbs_clk clknet_0_io_wbs_clk clknet_2_3__leaf_io_wbs_clk vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_170_ operation _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_437_ net79 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_299_ net108 _160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_368_ _067_ _032_ clknet_2_2__leaf_io_wbs_clk net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input52_I dout_mem1[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output139_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_222_ _097_ _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__300__I _160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_205_ _096_ _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__231__S _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input15_I dout_mem0[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__226__S _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I dout_mem0[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output121_I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output219_I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input82_I io_wbs_datwr[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_453_ net96 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_384_ net67 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__303__I _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__201__I1 _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__360__D _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__268__I1 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__259__I1 _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_436_ net78 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__348__CLK clknet_2_0__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_298_ _159_ _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_367_ _066_ _031_ clknet_2_3__leaf_io_wbs_clk net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__234__S _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input45_I dout_mem1[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_221_ _108_ _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__229__S _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_419_ net94 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output151_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__401__I net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_204_ net212 _095_ _093_ _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__311__I _163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output199_I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__306__I _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__216__I _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__237__S _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__358__D _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input75_I io_wbs_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_452_ net95 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_383_ net65 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__404__I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_435_ net77 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_366_ _065_ _030_ clknet_2_3__leaf_io_wbs_clk net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_2_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_297_ _159_ _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__314__I _163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input38_I dout_mem1[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_220_ net207 _107_ _105_ _108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__309__I _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_418_ net93 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_349_ _048_ _013_ clknet_2_1__leaf_io_wbs_clk net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__366__D _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__338__CLK clknet_2_1__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_203_ net15 net47 _087_ _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__412__I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__240__I0 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__231__I0 net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input20_I dout_mem0[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__407__I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__317__I _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__204__I0 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input68_I io_wbs_adr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_451_ net94 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_382_ net74 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__371__CLK clknet_2_1__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__420__I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_434_ net107 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_365_ _064_ _029_ clknet_2_3__leaf_io_wbs_clk net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_296_ _159_ _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__330__I _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_2__f_io_wbs_clk_I clknet_0_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__415__I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_417_ net92 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__325__I _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_279_ net209 _149_ _145_ _150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_348_ _047_ _012_ clknet_2_0__leaf_io_wbs_clk net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__261__S _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input50_I dout_mem1[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output137_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_202_ _094_ _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input98_I io_wbs_datwr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__240__I1 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__231__I1 _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input13_I dout_mem0[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__423__I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input5_I dout_mem0[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__204__I1 _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output217_I net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_381_ net73 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_450_ net93 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__418__I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_2_0__f_io_wbs_clk clknet_0_io_wbs_clk clknet_2_0__leaf_io_wbs_clk vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_5_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__189__I0 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__174__S _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input80_I io_wbs_datwr[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output167_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_433_ net106 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_295_ _159_ _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_364_ _063_ _028_ clknet_2_3__leaf_io_wbs_clk net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__259__S _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__169__S _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__431__I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_416_ net91 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_278_ net12 net44 _076_ _149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_347_ _046_ _011_ clknet_2_0__leaf_io_wbs_clk net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__361__CLK clknet_2_3__leaf_io_wbs_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput230 net230 web_mem0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input43_I dout_mem1[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__426__I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_201_ net213 _092_ _093_ _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__336__I _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__182__S _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output197_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_380_ net72 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__434__I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

