// This is the unpowered netlist.
module wb_mux (io_wbs_ack,
    io_wbs_ack_0,
    io_wbs_ack_1,
    io_wbs_cyc,
    io_wbs_cyc_0,
    io_wbs_cyc_1,
    io_wbs_stb,
    io_wbs_stb_0,
    io_wbs_stb_1,
    io_wbs_we,
    io_wbs_we_0,
    io_wbs_we_1,
    io_wbs_adr,
    io_wbs_adr_0,
    io_wbs_adr_1,
    io_wbs_datrd,
    io_wbs_datrd_0,
    io_wbs_datrd_1,
    io_wbs_datwr,
    io_wbs_datwr_0,
    io_wbs_datwr_1,
    io_wbs_sel,
    io_wbs_sel_0,
    io_wbs_sel_1);
 output io_wbs_ack;
 input io_wbs_ack_0;
 input io_wbs_ack_1;
 input io_wbs_cyc;
 output io_wbs_cyc_0;
 output io_wbs_cyc_1;
 input io_wbs_stb;
 output io_wbs_stb_0;
 output io_wbs_stb_1;
 input io_wbs_we;
 output io_wbs_we_0;
 output io_wbs_we_1;
 input [31:0] io_wbs_adr;
 output [31:0] io_wbs_adr_0;
 output [31:0] io_wbs_adr_1;
 output [31:0] io_wbs_datrd;
 input [31:0] io_wbs_datrd_0;
 input [31:0] io_wbs_datrd_1;
 input [31:0] io_wbs_datwr;
 output [31:0] io_wbs_datwr_0;
 output [31:0] io_wbs_datwr_1;
 input [3:0] io_wbs_sel;
 output [3:0] io_wbs_sel_0;
 output [3:0] io_wbs_sel_1;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _100_ (.I(net2),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _101_ (.A1(net16),
    .A2(net15),
    .A3(net18),
    .A4(net17),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _102_ (.A1(net27),
    .A2(net26),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _103_ (.A1(net24),
    .A2(net23),
    .A3(_001_),
    .A4(_002_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _104_ (.A1(net11),
    .A2(net10),
    .A3(net13),
    .A4(net12),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _105_ (.A1(net20),
    .A2(net19),
    .A3(net22),
    .A4(net21),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _106_ (.A1(_004_),
    .A2(_005_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _107_ (.A1(net9),
    .A2(net8),
    .A3(net7),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _108_ (.A1(net6),
    .A2(_003_),
    .A3(_006_),
    .A4(_007_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _109_ (.I(_008_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _110_ (.I(_009_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _111_ (.I(_010_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _112_ (.I(net6),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _113_ (.A1(_012_),
    .A2(_003_),
    .A3(_006_),
    .A4(_007_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _114_ (.I(_013_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _115_ (.I(_014_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _116_ (.I(_015_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _117_ (.I(net1),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _118_ (.A1(_000_),
    .A2(_011_),
    .B1(_016_),
    .B2(_017_),
    .ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _119_ (.I(net68),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _120_ (.I(net36),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _121_ (.A1(_018_),
    .A2(_011_),
    .B1(_016_),
    .B2(_019_),
    .ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _122_ (.I(net79),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _123_ (.I(_008_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _124_ (.I(_021_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _125_ (.I(_013_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _126_ (.I(_023_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _127_ (.I(net47),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _128_ (.A1(_020_),
    .A2(_022_),
    .B1(_024_),
    .B2(_025_),
    .ZN(net216));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _129_ (.I(net90),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _130_ (.I(net58),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _131_ (.A1(_026_),
    .A2(_022_),
    .B1(_024_),
    .B2(_027_),
    .ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _132_ (.I(net93),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _133_ (.I(net61),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _134_ (.A1(_028_),
    .A2(_022_),
    .B1(_024_),
    .B2(_029_),
    .ZN(net230));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _135_ (.I(net94),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _136_ (.I(net62),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _137_ (.A1(_030_),
    .A2(_022_),
    .B1(_024_),
    .B2(_031_),
    .ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _138_ (.I(net95),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _139_ (.I(_021_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _140_ (.I(_023_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _141_ (.I(net63),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _142_ (.A1(_032_),
    .A2(_033_),
    .B1(_034_),
    .B2(_035_),
    .ZN(net232));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _143_ (.I(net96),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _144_ (.I(net64),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _145_ (.A1(_036_),
    .A2(_033_),
    .B1(_034_),
    .B2(_037_),
    .ZN(net233));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _146_ (.I(net97),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _147_ (.I(net65),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _148_ (.A1(_038_),
    .A2(_033_),
    .B1(_034_),
    .B2(_039_),
    .ZN(net234));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _149_ (.I(net98),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _150_ (.I(net66),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _151_ (.A1(_040_),
    .A2(_033_),
    .B1(_034_),
    .B2(_041_),
    .ZN(net235));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _152_ (.I(net99),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _153_ (.I(_021_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _154_ (.I(_023_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _155_ (.I(net67),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _156_ (.A1(_042_),
    .A2(_043_),
    .B1(_044_),
    .B2(_045_),
    .ZN(net236));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _157_ (.I(net69),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _158_ (.I(net37),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _159_ (.A1(_046_),
    .A2(_043_),
    .B1(_044_),
    .B2(_047_),
    .ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _160_ (.I(net70),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _161_ (.I(net38),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _162_ (.A1(_048_),
    .A2(_043_),
    .B1(_044_),
    .B2(_049_),
    .ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _163_ (.I(net71),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _164_ (.I(net39),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _165_ (.A1(_050_),
    .A2(_043_),
    .B1(_044_),
    .B2(_051_),
    .ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _166_ (.I(net72),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _167_ (.I(_021_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _168_ (.I(_023_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _169_ (.I(net40),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _170_ (.A1(_052_),
    .A2(_053_),
    .B1(_054_),
    .B2(_055_),
    .ZN(net209));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _171_ (.I(net73),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _172_ (.I(net41),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _173_ (.A1(_056_),
    .A2(_053_),
    .B1(_054_),
    .B2(_057_),
    .ZN(net210));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _174_ (.I(net74),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _175_ (.I(net42),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _176_ (.A1(_058_),
    .A2(_053_),
    .B1(_054_),
    .B2(_059_),
    .ZN(net211));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _177_ (.I(net75),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _178_ (.I(net43),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _179_ (.A1(_060_),
    .A2(_053_),
    .B1(_054_),
    .B2(_061_),
    .ZN(net212));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _180_ (.I(net76),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _181_ (.I(_009_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _182_ (.I(_014_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _183_ (.I(net44),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _184_ (.A1(_062_),
    .A2(_063_),
    .B1(_064_),
    .B2(_065_),
    .ZN(net213));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _185_ (.I(net77),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _186_ (.I(net45),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _187_ (.A1(_066_),
    .A2(_063_),
    .B1(_064_),
    .B2(_067_),
    .ZN(net214));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _188_ (.I(net78),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _189_ (.I(net46),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _190_ (.A1(_068_),
    .A2(_063_),
    .B1(_064_),
    .B2(_069_),
    .ZN(net215));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _191_ (.I(net80),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _192_ (.I(net48),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _193_ (.A1(_070_),
    .A2(_063_),
    .B1(_064_),
    .B2(_071_),
    .ZN(net217));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _194_ (.I(net81),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _195_ (.I(_009_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _196_ (.I(_014_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _197_ (.I(net49),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _198_ (.A1(_072_),
    .A2(_073_),
    .B1(_074_),
    .B2(_075_),
    .ZN(net218));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _199_ (.I(net82),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _200_ (.I(net50),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _201_ (.A1(_076_),
    .A2(_073_),
    .B1(_074_),
    .B2(_077_),
    .ZN(net219));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _202_ (.I(net83),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _203_ (.I(net51),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _204_ (.A1(_078_),
    .A2(_073_),
    .B1(_074_),
    .B2(_079_),
    .ZN(net220));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _205_ (.I(net84),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _206_ (.I(net52),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _207_ (.A1(_080_),
    .A2(_073_),
    .B1(_074_),
    .B2(_081_),
    .ZN(net221));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _208_ (.I(net85),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _209_ (.I(_009_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _210_ (.I(_014_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _211_ (.I(net53),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _212_ (.A1(_082_),
    .A2(_083_),
    .B1(_084_),
    .B2(_085_),
    .ZN(net222));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _213_ (.I(net86),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _214_ (.I(net54),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _215_ (.A1(_086_),
    .A2(_083_),
    .B1(_084_),
    .B2(_087_),
    .ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _216_ (.I(net87),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _217_ (.I(net55),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _218_ (.A1(_088_),
    .A2(_083_),
    .B1(_084_),
    .B2(_089_),
    .ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _219_ (.I(net88),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _220_ (.I(net56),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _221_ (.A1(_090_),
    .A2(_083_),
    .B1(_084_),
    .B2(_091_),
    .ZN(net225));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _222_ (.I(net89),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _223_ (.I(net57),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _224_ (.A1(_092_),
    .A2(_010_),
    .B1(_015_),
    .B2(_093_),
    .ZN(net226));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _225_ (.I(net91),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _226_ (.I(net59),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _227_ (.A1(_094_),
    .A2(_010_),
    .B1(_015_),
    .B2(_095_),
    .ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _228_ (.I(net92),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _229_ (.I(net60),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _230_ (.A1(_096_),
    .A2(_010_),
    .B1(_015_),
    .B2(_097_),
    .ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _231_ (.I(net136),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _232_ (.A1(_098_),
    .A2(_016_),
    .ZN(net309));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _233_ (.I(net35),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _234_ (.A1(_099_),
    .A2(_016_),
    .ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _235_ (.A1(_098_),
    .A2(_011_),
    .ZN(net310));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _236_ (.A1(_099_),
    .A2(_011_),
    .ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _237_ (.I(net3),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _238_ (.I(net14),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _239_ (.I(net25),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _240_ (.I(net28),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _241_ (.I(net29),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _242_ (.I(net30),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _243_ (.I(net31),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _244_ (.I(net32),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _245_ (.I(net33),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _246_ (.I(net34),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _247_ (.I(net4),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _248_ (.I(net5),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _249_ (.I(net6),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _250_ (.I(net7),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _251_ (.I(net8),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _252_ (.I(net9),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _253_ (.I(net10),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _254_ (.I(net11),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _255_ (.I(net12),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _256_ (.I(net13),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _257_ (.I(net15),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _258_ (.I(net16),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _259_ (.I(net17),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _260_ (.I(net18),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _261_ (.I(net19),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _262_ (.I(net20),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _263_ (.I(net21),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _264_ (.I(net22),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _265_ (.I(net23),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _266_ (.I(net24),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _267_ (.I(net26),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _268_ (.I(net27),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _269_ (.I(net3),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _270_ (.I(net14),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _271_ (.I(net25),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _272_ (.I(net28),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _273_ (.I(net29),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _274_ (.I(net30),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _275_ (.I(net31),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _276_ (.I(net32),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _277_ (.I(net33),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _278_ (.I(net34),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _279_ (.I(net4),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _280_ (.I(net5),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _281_ (.I(net6),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _282_ (.I(net7),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _283_ (.I(net8),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _284_ (.I(net9),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _285_ (.I(net10),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _286_ (.I(net11),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _287_ (.I(net12),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _288_ (.I(net13),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _289_ (.I(net15),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _290_ (.I(net16),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _291_ (.I(net17),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _292_ (.I(net18),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _293_ (.I(net19),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _294_ (.I(net20),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _295_ (.I(net21),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _296_ (.I(net22),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _297_ (.I(net23),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _298_ (.I(net24),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _299_ (.I(net26),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _300_ (.I(net27),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _301_ (.I(net100),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _302_ (.I(net111),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _303_ (.I(net122),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _304_ (.I(net125),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _305_ (.I(net126),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _306_ (.I(net127),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _307_ (.I(net128),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _308_ (.I(net129),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _309_ (.I(net130),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _310_ (.I(net131),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _311_ (.I(net101),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _312_ (.I(net102),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _313_ (.I(net103),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _314_ (.I(net104),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _315_ (.I(net105),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _316_ (.I(net106),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _317_ (.I(net107),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _318_ (.I(net108),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _319_ (.I(net109),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _320_ (.I(net110),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _321_ (.I(net112),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _322_ (.I(net113),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _323_ (.I(net114),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _324_ (.I(net115),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _325_ (.I(net116),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _326_ (.I(net117),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _327_ (.I(net118),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _328_ (.I(net119),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _329_ (.I(net120),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _330_ (.I(net121),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _331_ (.I(net123),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _332_ (.I(net124),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _333_ (.I(net100),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _334_ (.I(net111),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _335_ (.I(net122),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _336_ (.I(net125),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _337_ (.I(net126),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _338_ (.I(net127),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _339_ (.I(net128),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _340_ (.I(net129),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _341_ (.I(net130),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _342_ (.I(net131),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _343_ (.I(net101),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _344_ (.I(net102),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _345_ (.I(net103),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _346_ (.I(net104),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _347_ (.I(net105),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _348_ (.I(net106),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _349_ (.I(net107),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _350_ (.I(net108),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _351_ (.I(net109),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _352_ (.I(net110),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _353_ (.I(net112),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _354_ (.I(net113),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _355_ (.I(net114),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _356_ (.I(net115),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _357_ (.I(net116),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _358_ (.I(net117),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _359_ (.I(net118),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _360_ (.I(net119),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _361_ (.I(net120),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _362_ (.I(net121),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _363_ (.I(net123),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _364_ (.I(net124),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _365_ (.I(net132),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _366_ (.I(net133),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _367_ (.I(net134),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _368_ (.I(net135),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _369_ (.I(net132),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _370_ (.I(net133),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _371_ (.I(net134),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _372_ (.I(net135),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _373_ (.I(net137),
    .Z(net311));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _374_ (.I(net137),
    .Z(net312));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_wbs_ack_0),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(io_wbs_ack_1),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_wbs_adr[0]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_wbs_adr[10]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(io_wbs_adr[11]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(io_wbs_adr[12]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input7 (.I(io_wbs_adr[13]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input8 (.I(io_wbs_adr[14]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input9 (.I(io_wbs_adr[15]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(io_wbs_adr[16]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(io_wbs_adr[17]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(io_wbs_adr[18]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(io_wbs_adr[19]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(io_wbs_adr[1]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(io_wbs_adr[20]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(io_wbs_adr[21]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(io_wbs_adr[22]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(io_wbs_adr[23]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input19 (.I(io_wbs_adr[24]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input20 (.I(io_wbs_adr[25]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input21 (.I(io_wbs_adr[26]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input22 (.I(io_wbs_adr[27]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input23 (.I(io_wbs_adr[28]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input24 (.I(io_wbs_adr[29]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input25 (.I(io_wbs_adr[2]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input26 (.I(io_wbs_adr[30]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input27 (.I(io_wbs_adr[31]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input28 (.I(io_wbs_adr[3]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input29 (.I(io_wbs_adr[4]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input30 (.I(io_wbs_adr[5]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input31 (.I(io_wbs_adr[6]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input32 (.I(io_wbs_adr[7]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input33 (.I(io_wbs_adr[8]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input34 (.I(io_wbs_adr[9]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input35 (.I(io_wbs_cyc),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input36 (.I(io_wbs_datrd_0[0]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input37 (.I(io_wbs_datrd_0[10]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input38 (.I(io_wbs_datrd_0[11]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input39 (.I(io_wbs_datrd_0[12]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input40 (.I(io_wbs_datrd_0[13]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input41 (.I(io_wbs_datrd_0[14]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input42 (.I(io_wbs_datrd_0[15]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input43 (.I(io_wbs_datrd_0[16]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input44 (.I(io_wbs_datrd_0[17]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input45 (.I(io_wbs_datrd_0[18]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input46 (.I(io_wbs_datrd_0[19]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input47 (.I(io_wbs_datrd_0[1]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input48 (.I(io_wbs_datrd_0[20]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input49 (.I(io_wbs_datrd_0[21]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input50 (.I(io_wbs_datrd_0[22]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input51 (.I(io_wbs_datrd_0[23]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input52 (.I(io_wbs_datrd_0[24]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input53 (.I(io_wbs_datrd_0[25]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input54 (.I(io_wbs_datrd_0[26]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input55 (.I(io_wbs_datrd_0[27]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input56 (.I(io_wbs_datrd_0[28]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input57 (.I(io_wbs_datrd_0[29]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input58 (.I(io_wbs_datrd_0[2]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input59 (.I(io_wbs_datrd_0[30]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input60 (.I(io_wbs_datrd_0[31]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input61 (.I(io_wbs_datrd_0[3]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input62 (.I(io_wbs_datrd_0[4]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input63 (.I(io_wbs_datrd_0[5]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input64 (.I(io_wbs_datrd_0[6]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input65 (.I(io_wbs_datrd_0[7]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input66 (.I(io_wbs_datrd_0[8]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input67 (.I(io_wbs_datrd_0[9]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input68 (.I(io_wbs_datrd_1[0]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input69 (.I(io_wbs_datrd_1[10]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input70 (.I(io_wbs_datrd_1[11]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input71 (.I(io_wbs_datrd_1[12]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input72 (.I(io_wbs_datrd_1[13]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input73 (.I(io_wbs_datrd_1[14]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input74 (.I(io_wbs_datrd_1[15]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input75 (.I(io_wbs_datrd_1[16]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input76 (.I(io_wbs_datrd_1[17]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input77 (.I(io_wbs_datrd_1[18]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input78 (.I(io_wbs_datrd_1[19]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input79 (.I(io_wbs_datrd_1[1]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input80 (.I(io_wbs_datrd_1[20]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input81 (.I(io_wbs_datrd_1[21]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input82 (.I(io_wbs_datrd_1[22]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input83 (.I(io_wbs_datrd_1[23]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input84 (.I(io_wbs_datrd_1[24]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input85 (.I(io_wbs_datrd_1[25]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input86 (.I(io_wbs_datrd_1[26]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input87 (.I(io_wbs_datrd_1[27]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input88 (.I(io_wbs_datrd_1[28]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input89 (.I(io_wbs_datrd_1[29]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input90 (.I(io_wbs_datrd_1[2]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input91 (.I(io_wbs_datrd_1[30]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input92 (.I(io_wbs_datrd_1[31]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input93 (.I(io_wbs_datrd_1[3]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input94 (.I(io_wbs_datrd_1[4]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input95 (.I(io_wbs_datrd_1[5]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input96 (.I(io_wbs_datrd_1[6]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input97 (.I(io_wbs_datrd_1[7]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input98 (.I(io_wbs_datrd_1[8]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input99 (.I(io_wbs_datrd_1[9]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input100 (.I(io_wbs_datwr[0]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input101 (.I(io_wbs_datwr[10]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input102 (.I(io_wbs_datwr[11]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input103 (.I(io_wbs_datwr[12]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input104 (.I(io_wbs_datwr[13]),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input105 (.I(io_wbs_datwr[14]),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input106 (.I(io_wbs_datwr[15]),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input107 (.I(io_wbs_datwr[16]),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input108 (.I(io_wbs_datwr[17]),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input109 (.I(io_wbs_datwr[18]),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input110 (.I(io_wbs_datwr[19]),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input111 (.I(io_wbs_datwr[1]),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input112 (.I(io_wbs_datwr[20]),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input113 (.I(io_wbs_datwr[21]),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input114 (.I(io_wbs_datwr[22]),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input115 (.I(io_wbs_datwr[23]),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input116 (.I(io_wbs_datwr[24]),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input117 (.I(io_wbs_datwr[25]),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input118 (.I(io_wbs_datwr[26]),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input119 (.I(io_wbs_datwr[27]),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input120 (.I(io_wbs_datwr[28]),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input121 (.I(io_wbs_datwr[29]),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input122 (.I(io_wbs_datwr[2]),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input123 (.I(io_wbs_datwr[30]),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input124 (.I(io_wbs_datwr[31]),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input125 (.I(io_wbs_datwr[3]),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input126 (.I(io_wbs_datwr[4]),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input127 (.I(io_wbs_datwr[5]),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input128 (.I(io_wbs_datwr[6]),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input129 (.I(io_wbs_datwr[7]),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input130 (.I(io_wbs_datwr[8]),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input131 (.I(io_wbs_datwr[9]),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input132 (.I(io_wbs_sel[0]),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input133 (.I(io_wbs_sel[1]),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input134 (.I(io_wbs_sel[2]),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input135 (.I(io_wbs_sel[3]),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input136 (.I(io_wbs_stb),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input137 (.I(io_wbs_we),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output138 (.I(net138),
    .Z(io_wbs_ack));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output139 (.I(net139),
    .Z(io_wbs_adr_0[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output140 (.I(net140),
    .Z(io_wbs_adr_0[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output141 (.I(net141),
    .Z(io_wbs_adr_0[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output142 (.I(net142),
    .Z(io_wbs_adr_0[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output143 (.I(net143),
    .Z(io_wbs_adr_0[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output144 (.I(net144),
    .Z(io_wbs_adr_0[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output145 (.I(net145),
    .Z(io_wbs_adr_0[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output146 (.I(net146),
    .Z(io_wbs_adr_0[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output147 (.I(net147),
    .Z(io_wbs_adr_0[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output148 (.I(net148),
    .Z(io_wbs_adr_0[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output149 (.I(net149),
    .Z(io_wbs_adr_0[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output150 (.I(net150),
    .Z(io_wbs_adr_0[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output151 (.I(net151),
    .Z(io_wbs_adr_0[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output152 (.I(net152),
    .Z(io_wbs_adr_0[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output153 (.I(net153),
    .Z(io_wbs_adr_0[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output154 (.I(net154),
    .Z(io_wbs_adr_0[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output155 (.I(net155),
    .Z(io_wbs_adr_0[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output156 (.I(net156),
    .Z(io_wbs_adr_0[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output157 (.I(net157),
    .Z(io_wbs_adr_0[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output158 (.I(net158),
    .Z(io_wbs_adr_0[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output159 (.I(net159),
    .Z(io_wbs_adr_0[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output160 (.I(net160),
    .Z(io_wbs_adr_0[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output161 (.I(net161),
    .Z(io_wbs_adr_0[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output162 (.I(net162),
    .Z(io_wbs_adr_0[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output163 (.I(net163),
    .Z(io_wbs_adr_0[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output164 (.I(net164),
    .Z(io_wbs_adr_0[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output165 (.I(net165),
    .Z(io_wbs_adr_0[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output166 (.I(net166),
    .Z(io_wbs_adr_0[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output167 (.I(net167),
    .Z(io_wbs_adr_0[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output168 (.I(net168),
    .Z(io_wbs_adr_0[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output169 (.I(net169),
    .Z(io_wbs_adr_0[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output170 (.I(net170),
    .Z(io_wbs_adr_0[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output171 (.I(net171),
    .Z(io_wbs_adr_1[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output172 (.I(net172),
    .Z(io_wbs_adr_1[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output173 (.I(net173),
    .Z(io_wbs_adr_1[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output174 (.I(net174),
    .Z(io_wbs_adr_1[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output175 (.I(net175),
    .Z(io_wbs_adr_1[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output176 (.I(net176),
    .Z(io_wbs_adr_1[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output177 (.I(net177),
    .Z(io_wbs_adr_1[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output178 (.I(net178),
    .Z(io_wbs_adr_1[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output179 (.I(net179),
    .Z(io_wbs_adr_1[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output180 (.I(net180),
    .Z(io_wbs_adr_1[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output181 (.I(net181),
    .Z(io_wbs_adr_1[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output182 (.I(net182),
    .Z(io_wbs_adr_1[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output183 (.I(net183),
    .Z(io_wbs_adr_1[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output184 (.I(net184),
    .Z(io_wbs_adr_1[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output185 (.I(net185),
    .Z(io_wbs_adr_1[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output186 (.I(net186),
    .Z(io_wbs_adr_1[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output187 (.I(net187),
    .Z(io_wbs_adr_1[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output188 (.I(net188),
    .Z(io_wbs_adr_1[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output189 (.I(net189),
    .Z(io_wbs_adr_1[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output190 (.I(net190),
    .Z(io_wbs_adr_1[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output191 (.I(net191),
    .Z(io_wbs_adr_1[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output192 (.I(net192),
    .Z(io_wbs_adr_1[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output193 (.I(net193),
    .Z(io_wbs_adr_1[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output194 (.I(net194),
    .Z(io_wbs_adr_1[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output195 (.I(net195),
    .Z(io_wbs_adr_1[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output196 (.I(net196),
    .Z(io_wbs_adr_1[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output197 (.I(net197),
    .Z(io_wbs_adr_1[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output198 (.I(net198),
    .Z(io_wbs_adr_1[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output199 (.I(net199),
    .Z(io_wbs_adr_1[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output200 (.I(net200),
    .Z(io_wbs_adr_1[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output201 (.I(net201),
    .Z(io_wbs_adr_1[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output202 (.I(net202),
    .Z(io_wbs_adr_1[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output203 (.I(net203),
    .Z(io_wbs_cyc_0));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output204 (.I(net204),
    .Z(io_wbs_cyc_1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output205 (.I(net205),
    .Z(io_wbs_datrd[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output206 (.I(net206),
    .Z(io_wbs_datrd[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output207 (.I(net207),
    .Z(io_wbs_datrd[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output208 (.I(net208),
    .Z(io_wbs_datrd[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output209 (.I(net209),
    .Z(io_wbs_datrd[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output210 (.I(net210),
    .Z(io_wbs_datrd[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output211 (.I(net211),
    .Z(io_wbs_datrd[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output212 (.I(net212),
    .Z(io_wbs_datrd[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output213 (.I(net213),
    .Z(io_wbs_datrd[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output214 (.I(net214),
    .Z(io_wbs_datrd[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output215 (.I(net215),
    .Z(io_wbs_datrd[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output216 (.I(net216),
    .Z(io_wbs_datrd[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output217 (.I(net217),
    .Z(io_wbs_datrd[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output218 (.I(net218),
    .Z(io_wbs_datrd[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output219 (.I(net219),
    .Z(io_wbs_datrd[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output220 (.I(net220),
    .Z(io_wbs_datrd[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output221 (.I(net221),
    .Z(io_wbs_datrd[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output222 (.I(net222),
    .Z(io_wbs_datrd[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output223 (.I(net223),
    .Z(io_wbs_datrd[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output224 (.I(net224),
    .Z(io_wbs_datrd[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output225 (.I(net225),
    .Z(io_wbs_datrd[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output226 (.I(net226),
    .Z(io_wbs_datrd[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output227 (.I(net227),
    .Z(io_wbs_datrd[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output228 (.I(net228),
    .Z(io_wbs_datrd[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output229 (.I(net229),
    .Z(io_wbs_datrd[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output230 (.I(net230),
    .Z(io_wbs_datrd[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output231 (.I(net231),
    .Z(io_wbs_datrd[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output232 (.I(net232),
    .Z(io_wbs_datrd[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output233 (.I(net233),
    .Z(io_wbs_datrd[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output234 (.I(net234),
    .Z(io_wbs_datrd[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output235 (.I(net235),
    .Z(io_wbs_datrd[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output236 (.I(net236),
    .Z(io_wbs_datrd[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output237 (.I(net237),
    .Z(io_wbs_datwr_0[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output238 (.I(net238),
    .Z(io_wbs_datwr_0[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output239 (.I(net239),
    .Z(io_wbs_datwr_0[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output240 (.I(net240),
    .Z(io_wbs_datwr_0[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output241 (.I(net241),
    .Z(io_wbs_datwr_0[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output242 (.I(net242),
    .Z(io_wbs_datwr_0[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output243 (.I(net243),
    .Z(io_wbs_datwr_0[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output244 (.I(net244),
    .Z(io_wbs_datwr_0[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output245 (.I(net245),
    .Z(io_wbs_datwr_0[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output246 (.I(net246),
    .Z(io_wbs_datwr_0[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output247 (.I(net247),
    .Z(io_wbs_datwr_0[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output248 (.I(net248),
    .Z(io_wbs_datwr_0[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output249 (.I(net249),
    .Z(io_wbs_datwr_0[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output250 (.I(net250),
    .Z(io_wbs_datwr_0[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output251 (.I(net251),
    .Z(io_wbs_datwr_0[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output252 (.I(net252),
    .Z(io_wbs_datwr_0[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output253 (.I(net253),
    .Z(io_wbs_datwr_0[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output254 (.I(net254),
    .Z(io_wbs_datwr_0[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output255 (.I(net255),
    .Z(io_wbs_datwr_0[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output256 (.I(net256),
    .Z(io_wbs_datwr_0[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output257 (.I(net257),
    .Z(io_wbs_datwr_0[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output258 (.I(net258),
    .Z(io_wbs_datwr_0[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output259 (.I(net259),
    .Z(io_wbs_datwr_0[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output260 (.I(net260),
    .Z(io_wbs_datwr_0[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output261 (.I(net261),
    .Z(io_wbs_datwr_0[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output262 (.I(net262),
    .Z(io_wbs_datwr_0[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output263 (.I(net263),
    .Z(io_wbs_datwr_0[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output264 (.I(net264),
    .Z(io_wbs_datwr_0[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output265 (.I(net265),
    .Z(io_wbs_datwr_0[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output266 (.I(net266),
    .Z(io_wbs_datwr_0[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output267 (.I(net267),
    .Z(io_wbs_datwr_0[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output268 (.I(net268),
    .Z(io_wbs_datwr_0[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output269 (.I(net269),
    .Z(io_wbs_datwr_1[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output270 (.I(net270),
    .Z(io_wbs_datwr_1[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output271 (.I(net271),
    .Z(io_wbs_datwr_1[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output272 (.I(net272),
    .Z(io_wbs_datwr_1[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output273 (.I(net273),
    .Z(io_wbs_datwr_1[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output274 (.I(net274),
    .Z(io_wbs_datwr_1[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output275 (.I(net275),
    .Z(io_wbs_datwr_1[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output276 (.I(net276),
    .Z(io_wbs_datwr_1[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output277 (.I(net277),
    .Z(io_wbs_datwr_1[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output278 (.I(net278),
    .Z(io_wbs_datwr_1[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output279 (.I(net279),
    .Z(io_wbs_datwr_1[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output280 (.I(net280),
    .Z(io_wbs_datwr_1[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output281 (.I(net281),
    .Z(io_wbs_datwr_1[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output282 (.I(net282),
    .Z(io_wbs_datwr_1[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output283 (.I(net283),
    .Z(io_wbs_datwr_1[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output284 (.I(net284),
    .Z(io_wbs_datwr_1[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output285 (.I(net285),
    .Z(io_wbs_datwr_1[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output286 (.I(net286),
    .Z(io_wbs_datwr_1[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output287 (.I(net287),
    .Z(io_wbs_datwr_1[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output288 (.I(net288),
    .Z(io_wbs_datwr_1[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output289 (.I(net289),
    .Z(io_wbs_datwr_1[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output290 (.I(net290),
    .Z(io_wbs_datwr_1[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output291 (.I(net291),
    .Z(io_wbs_datwr_1[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output292 (.I(net292),
    .Z(io_wbs_datwr_1[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output293 (.I(net293),
    .Z(io_wbs_datwr_1[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output294 (.I(net294),
    .Z(io_wbs_datwr_1[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output295 (.I(net295),
    .Z(io_wbs_datwr_1[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output296 (.I(net296),
    .Z(io_wbs_datwr_1[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output297 (.I(net297),
    .Z(io_wbs_datwr_1[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output298 (.I(net298),
    .Z(io_wbs_datwr_1[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output299 (.I(net299),
    .Z(io_wbs_datwr_1[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output300 (.I(net300),
    .Z(io_wbs_datwr_1[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output301 (.I(net301),
    .Z(io_wbs_sel_0[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output302 (.I(net302),
    .Z(io_wbs_sel_0[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output303 (.I(net303),
    .Z(io_wbs_sel_0[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output304 (.I(net304),
    .Z(io_wbs_sel_0[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output305 (.I(net305),
    .Z(io_wbs_sel_1[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output306 (.I(net306),
    .Z(io_wbs_sel_1[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output307 (.I(net307),
    .Z(io_wbs_sel_1[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output308 (.I(net308),
    .Z(io_wbs_sel_1[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output309 (.I(net309),
    .Z(io_wbs_stb_0));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output310 (.I(net310),
    .Z(io_wbs_stb_1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output311 (.I(net311),
    .Z(io_wbs_we_0));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output312 (.I(net312),
    .Z(io_wbs_we_1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__113__A2 (.I(_003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__A2 (.I(_003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__113__A3 (.I(_006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__A3 (.I(_006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__I (.I(_008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__109__I (.I(_008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__209__I (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__195__I (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__I (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__110__I (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__236__A2 (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__A2 (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__121__A2 (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__118__A2 (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__125__I (.I(_013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__114__I (.I(_013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__I (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__I (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__I (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__115__I (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__A2 (.I(_016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__A2 (.I(_016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__121__B1 (.I(_016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__118__B1 (.I(_016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__I (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__I (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__140__I (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__126__I (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_wbs_ack_0));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_wbs_ack_1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_wbs_adr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_wbs_adr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_wbs_adr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_wbs_adr[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_wbs_adr[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_wbs_adr[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_wbs_adr[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_wbs_adr[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_wbs_adr[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_wbs_adr[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_wbs_adr[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(io_wbs_adr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_wbs_adr[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(io_wbs_adr[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(io_wbs_adr[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(io_wbs_adr[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(io_wbs_adr[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(io_wbs_adr[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(io_wbs_adr[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(io_wbs_adr[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(io_wbs_adr[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(io_wbs_adr[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(io_wbs_adr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(io_wbs_adr[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(io_wbs_adr[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(io_wbs_adr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(io_wbs_adr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(io_wbs_adr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(io_wbs_adr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(io_wbs_adr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(io_wbs_adr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(io_wbs_adr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(io_wbs_cyc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(io_wbs_datrd_0[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(io_wbs_datrd_0[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(io_wbs_datrd_0[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(io_wbs_datrd_0[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(io_wbs_datrd_0[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(io_wbs_datrd_0[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(io_wbs_datrd_0[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(io_wbs_datrd_0[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(io_wbs_datrd_0[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(io_wbs_datrd_0[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(io_wbs_datrd_0[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(io_wbs_datrd_0[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(io_wbs_datrd_0[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(io_wbs_datrd_0[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(io_wbs_datrd_0[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(io_wbs_datrd_0[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(io_wbs_datrd_0[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(io_wbs_datrd_0[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(io_wbs_datrd_0[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(io_wbs_datrd_0[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(io_wbs_datrd_0[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(io_wbs_datrd_0[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(io_wbs_datrd_0[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(io_wbs_datrd_0[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(io_wbs_datrd_0[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(io_wbs_datrd_0[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(io_wbs_datrd_0[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(io_wbs_datrd_0[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(io_wbs_datrd_0[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(io_wbs_datrd_0[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(io_wbs_datrd_0[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(io_wbs_datrd_0[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(io_wbs_datrd_1[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(io_wbs_datrd_1[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(io_wbs_datrd_1[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(io_wbs_datrd_1[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(io_wbs_datrd_1[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(io_wbs_datrd_1[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(io_wbs_datrd_1[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(io_wbs_datrd_1[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(io_wbs_datrd_1[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(io_wbs_datrd_1[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(io_wbs_datrd_1[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(io_wbs_datrd_1[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(io_wbs_datrd_1[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(io_wbs_datrd_1[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(io_wbs_datrd_1[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(io_wbs_datrd_1[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(io_wbs_datrd_1[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(io_wbs_datrd_1[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(io_wbs_datrd_1[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(io_wbs_datrd_1[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(io_wbs_datrd_1[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(io_wbs_datrd_1[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(io_wbs_datrd_1[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(io_wbs_datrd_1[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(io_wbs_datrd_1[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(io_wbs_datrd_1[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(io_wbs_datrd_1[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(io_wbs_datrd_1[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(io_wbs_datrd_1[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(io_wbs_datrd_1[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input98_I (.I(io_wbs_datrd_1[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input99_I (.I(io_wbs_datrd_1[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input100_I (.I(io_wbs_datwr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input101_I (.I(io_wbs_datwr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input102_I (.I(io_wbs_datwr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input103_I (.I(io_wbs_datwr[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input104_I (.I(io_wbs_datwr[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input105_I (.I(io_wbs_datwr[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input106_I (.I(io_wbs_datwr[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input107_I (.I(io_wbs_datwr[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input108_I (.I(io_wbs_datwr[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input109_I (.I(io_wbs_datwr[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input110_I (.I(io_wbs_datwr[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input111_I (.I(io_wbs_datwr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input112_I (.I(io_wbs_datwr[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input113_I (.I(io_wbs_datwr[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input114_I (.I(io_wbs_datwr[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input115_I (.I(io_wbs_datwr[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input116_I (.I(io_wbs_datwr[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input117_I (.I(io_wbs_datwr[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input118_I (.I(io_wbs_datwr[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input119_I (.I(io_wbs_datwr[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input120_I (.I(io_wbs_datwr[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input121_I (.I(io_wbs_datwr[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input122_I (.I(io_wbs_datwr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input123_I (.I(io_wbs_datwr[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input124_I (.I(io_wbs_datwr[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input125_I (.I(io_wbs_datwr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input126_I (.I(io_wbs_datwr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input127_I (.I(io_wbs_datwr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input128_I (.I(io_wbs_datwr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input129_I (.I(io_wbs_datwr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input130_I (.I(io_wbs_datwr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input131_I (.I(io_wbs_datwr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input132_I (.I(io_wbs_sel[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input133_I (.I(io_wbs_sel[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input134_I (.I(io_wbs_sel[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input135_I (.I(io_wbs_sel[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input136_I (.I(io_wbs_stb));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input137_I (.I(io_wbs_we));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__117__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__100__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__280__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__248__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__112__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__250__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__107__A3 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__283__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__107__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__107__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__285__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__A4 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__288__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__A3 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__101__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__101__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__101__A4 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__101__A3 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__105__A2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__105__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__105__A4 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__105__A3 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__103__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__103__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__102__A2 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__102__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__158__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__164__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__186__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__189__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__127__I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__192__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__211__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__217__I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__130__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__133__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__141__I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__155__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__119__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__157__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__166__I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__171__I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__177__I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__122__I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__191__I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__194__I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__199__I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__202__I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__208__I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__213__I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__216__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__222__I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__129__I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__225__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__135__I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__143__I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__146__I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__318__I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__321__I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__323__I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__324__I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__326__I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__359__I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__330__I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__332__I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__339__I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__341__I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__372__I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__374__I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output138_I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output139_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output140_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output141_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output142_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output143_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output144_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output145_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output149_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output152_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output153_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output154_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output155_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output156_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output157_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output158_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output159_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output160_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output161_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output162_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output163_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output164_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output166_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output167_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output169_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output170_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output172_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output173_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output174_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output175_I (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output177_I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output180_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output185_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output186_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output188_I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output189_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output191_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output194_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output195_I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output204_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output205_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output206_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output207_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output208_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output209_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output210_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output211_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output212_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output213_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output214_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output215_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output216_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output217_I (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output218_I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output219_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output220_I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output221_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output222_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output223_I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output224_I (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output225_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output226_I (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output227_I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output228_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output229_I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output230_I (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output231_I (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output232_I (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output233_I (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output234_I (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output235_I (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output236_I (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output237_I (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output238_I (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output239_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output240_I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output241_I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output242_I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output243_I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output244_I (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output245_I (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output246_I (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output247_I (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output248_I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output249_I (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output250_I (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output251_I (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output252_I (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output253_I (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output254_I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output255_I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output256_I (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output257_I (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output258_I (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output259_I (.I(net259));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output260_I (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output261_I (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output262_I (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output263_I (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output264_I (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output265_I (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output266_I (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output267_I (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output268_I (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output269_I (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output270_I (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output271_I (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output272_I (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output273_I (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output274_I (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output275_I (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output276_I (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output277_I (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output278_I (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output279_I (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output280_I (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output281_I (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output282_I (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output283_I (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output284_I (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output285_I (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output286_I (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output287_I (.I(net287));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output288_I (.I(net288));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output289_I (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output290_I (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output291_I (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output292_I (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output293_I (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output294_I (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output295_I (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output296_I (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output297_I (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output298_I (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output299_I (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output300_I (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output305_I (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output306_I (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output307_I (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output308_I (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output310_I (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output312_I (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_687 ();
endmodule

