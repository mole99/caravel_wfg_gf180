magic
tech gf180mcuC
magscale 1 10
timestamp 1669807972
<< metal1 >>
rect 1344 76858 78624 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 78624 76858
rect 1344 76772 78624 76806
rect 1344 76074 78624 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 78624 76074
rect 1344 75988 78624 76022
rect 1344 75290 78624 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 78624 75290
rect 1344 75204 78624 75238
rect 3042 74846 3054 74898
rect 3106 74846 3118 74898
rect 75058 74846 75070 74898
rect 75122 74846 75134 74898
rect 76850 74846 76862 74898
rect 76914 74846 76926 74898
rect 3614 74786 3666 74798
rect 2034 74734 2046 74786
rect 2098 74734 2110 74786
rect 3614 74722 3666 74734
rect 4062 74786 4114 74798
rect 76066 74734 76078 74786
rect 76130 74734 76142 74786
rect 77858 74734 77870 74786
rect 77922 74734 77934 74786
rect 4062 74722 4114 74734
rect 1344 74506 78624 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 78624 74506
rect 1344 74420 78624 74454
rect 3042 74062 3054 74114
rect 3106 74062 3118 74114
rect 3614 74002 3666 74014
rect 2146 73950 2158 74002
rect 2210 73950 2222 74002
rect 3614 73938 3666 73950
rect 4398 74002 4450 74014
rect 4398 73938 4450 73950
rect 77310 74002 77362 74014
rect 77310 73938 77362 73950
rect 78094 74002 78146 74014
rect 78094 73938 78146 73950
rect 3950 73890 4002 73902
rect 3950 73826 4002 73838
rect 73390 73890 73442 73902
rect 73390 73826 73442 73838
rect 77758 73890 77810 73902
rect 77758 73826 77810 73838
rect 1344 73722 78624 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 78624 73722
rect 1344 73636 78624 73670
rect 73726 73554 73778 73566
rect 73726 73490 73778 73502
rect 69358 73442 69410 73454
rect 69358 73378 69410 73390
rect 73838 73442 73890 73454
rect 73838 73378 73890 73390
rect 70030 73330 70082 73342
rect 3042 73278 3054 73330
rect 3106 73278 3118 73330
rect 75058 73278 75070 73330
rect 75122 73278 75134 73330
rect 76850 73278 76862 73330
rect 76914 73278 76926 73330
rect 70030 73266 70082 73278
rect 3614 73218 3666 73230
rect 2034 73166 2046 73218
rect 2098 73166 2110 73218
rect 3614 73154 3666 73166
rect 69246 73218 69298 73230
rect 69246 73154 69298 73166
rect 72494 73218 72546 73230
rect 76066 73166 76078 73218
rect 76130 73166 76142 73218
rect 77858 73166 77870 73218
rect 77922 73166 77934 73218
rect 72494 73154 72546 73166
rect 69134 73106 69186 73118
rect 69134 73042 69186 73054
rect 73614 73106 73666 73118
rect 73614 73042 73666 73054
rect 1344 72938 78624 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 78624 72938
rect 1344 72852 78624 72886
rect 74062 72658 74114 72670
rect 74062 72594 74114 72606
rect 74174 72658 74226 72670
rect 74174 72594 74226 72606
rect 74622 72658 74674 72670
rect 74622 72594 74674 72606
rect 72158 72546 72210 72558
rect 75070 72546 75122 72558
rect 3042 72494 3054 72546
rect 3106 72494 3118 72546
rect 73042 72494 73054 72546
rect 73106 72494 73118 72546
rect 72158 72482 72210 72494
rect 75070 72482 75122 72494
rect 69358 72434 69410 72446
rect 2146 72382 2158 72434
rect 2210 72382 2222 72434
rect 69358 72370 69410 72382
rect 69470 72434 69522 72446
rect 69470 72370 69522 72382
rect 71822 72434 71874 72446
rect 71822 72370 71874 72382
rect 73278 72434 73330 72446
rect 73278 72370 73330 72382
rect 3502 72322 3554 72334
rect 3502 72258 3554 72270
rect 68686 72322 68738 72334
rect 68686 72258 68738 72270
rect 69582 72322 69634 72334
rect 69582 72258 69634 72270
rect 73950 72322 74002 72334
rect 73950 72258 74002 72270
rect 1344 72154 78624 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 78624 72154
rect 1344 72068 78624 72102
rect 72494 71986 72546 71998
rect 72494 71922 72546 71934
rect 73390 71986 73442 71998
rect 73390 71922 73442 71934
rect 74062 71986 74114 71998
rect 74062 71922 74114 71934
rect 71150 71874 71202 71886
rect 71150 71810 71202 71822
rect 70702 71762 70754 71774
rect 3042 71710 3054 71762
rect 3106 71710 3118 71762
rect 70702 71698 70754 71710
rect 71486 71762 71538 71774
rect 72258 71710 72270 71762
rect 72322 71710 72334 71762
rect 75058 71710 75070 71762
rect 75122 71710 75134 71762
rect 76850 71710 76862 71762
rect 76914 71710 76926 71762
rect 71486 71698 71538 71710
rect 3614 71650 3666 71662
rect 2034 71598 2046 71650
rect 2098 71598 2110 71650
rect 3614 71586 3666 71598
rect 73502 71650 73554 71662
rect 73502 71586 73554 71598
rect 74174 71650 74226 71662
rect 76066 71598 76078 71650
rect 76130 71598 76142 71650
rect 77858 71598 77870 71650
rect 77922 71598 77934 71650
rect 74174 71586 74226 71598
rect 1344 71370 78624 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 78624 71370
rect 1344 71284 78624 71318
rect 3042 70926 3054 70978
rect 3106 70926 3118 70978
rect 71698 70926 71710 70978
rect 71762 70926 71774 70978
rect 70590 70866 70642 70878
rect 2146 70814 2158 70866
rect 2210 70814 2222 70866
rect 70590 70802 70642 70814
rect 70926 70866 70978 70878
rect 70926 70802 70978 70814
rect 71934 70866 71986 70878
rect 71934 70802 71986 70814
rect 3502 70754 3554 70766
rect 3502 70690 3554 70702
rect 70142 70754 70194 70766
rect 70142 70690 70194 70702
rect 72382 70754 72434 70766
rect 72382 70690 72434 70702
rect 72830 70754 72882 70766
rect 72830 70690 72882 70702
rect 73726 70754 73778 70766
rect 73726 70690 73778 70702
rect 74398 70754 74450 70766
rect 74398 70690 74450 70702
rect 78206 70754 78258 70766
rect 78206 70690 78258 70702
rect 1344 70586 78624 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 78624 70586
rect 1344 70500 78624 70534
rect 71262 70418 71314 70430
rect 71262 70354 71314 70366
rect 69918 70306 69970 70318
rect 69918 70242 69970 70254
rect 69470 70194 69522 70206
rect 3042 70142 3054 70194
rect 3106 70142 3118 70194
rect 69470 70130 69522 70142
rect 70254 70194 70306 70206
rect 70254 70130 70306 70142
rect 70926 70194 70978 70206
rect 70926 70130 70978 70142
rect 71710 70194 71762 70206
rect 76850 70142 76862 70194
rect 76914 70142 76926 70194
rect 71710 70130 71762 70142
rect 3614 70082 3666 70094
rect 2034 70030 2046 70082
rect 2098 70030 2110 70082
rect 77858 70030 77870 70082
rect 77922 70030 77934 70082
rect 3614 70018 3666 70030
rect 1344 69802 78624 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 78624 69802
rect 1344 69716 78624 69750
rect 1822 69298 1874 69310
rect 1822 69234 1874 69246
rect 2718 69298 2770 69310
rect 2718 69234 2770 69246
rect 3950 69298 4002 69310
rect 3950 69234 4002 69246
rect 69358 69298 69410 69310
rect 69358 69234 69410 69246
rect 69694 69298 69746 69310
rect 69694 69234 69746 69246
rect 70254 69298 70306 69310
rect 70254 69234 70306 69246
rect 70590 69298 70642 69310
rect 70590 69234 70642 69246
rect 76526 69298 76578 69310
rect 76526 69234 76578 69246
rect 78094 69298 78146 69310
rect 78094 69234 78146 69246
rect 2158 69186 2210 69198
rect 2158 69122 2210 69134
rect 3054 69186 3106 69198
rect 3054 69122 3106 69134
rect 3502 69186 3554 69198
rect 3502 69122 3554 69134
rect 71150 69186 71202 69198
rect 71150 69122 71202 69134
rect 76190 69186 76242 69198
rect 76190 69122 76242 69134
rect 77310 69186 77362 69198
rect 77310 69122 77362 69134
rect 77758 69186 77810 69198
rect 77758 69122 77810 69134
rect 1344 69018 78624 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 78624 69018
rect 1344 68932 78624 68966
rect 2158 68738 2210 68750
rect 2158 68674 2210 68686
rect 3054 68738 3106 68750
rect 3054 68674 3106 68686
rect 67342 68738 67394 68750
rect 67342 68674 67394 68686
rect 68686 68738 68738 68750
rect 68686 68674 68738 68686
rect 76862 68738 76914 68750
rect 76862 68674 76914 68686
rect 77758 68738 77810 68750
rect 77758 68674 77810 68686
rect 2718 68626 2770 68638
rect 1922 68574 1934 68626
rect 1986 68574 1998 68626
rect 2718 68562 2770 68574
rect 3502 68626 3554 68638
rect 3502 68562 3554 68574
rect 75966 68626 76018 68638
rect 75966 68562 76018 68574
rect 77198 68626 77250 68638
rect 77970 68574 77982 68626
rect 78034 68574 78046 68626
rect 77198 68562 77250 68574
rect 66782 68514 66834 68526
rect 66782 68450 66834 68462
rect 67790 68514 67842 68526
rect 67790 68450 67842 68462
rect 69918 68514 69970 68526
rect 69918 68450 69970 68462
rect 76414 68514 76466 68526
rect 76414 68450 76466 68462
rect 67902 68402 67954 68414
rect 67902 68338 67954 68350
rect 68798 68402 68850 68414
rect 68798 68338 68850 68350
rect 1344 68234 78624 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 78624 68234
rect 1344 68148 78624 68182
rect 2718 67954 2770 67966
rect 2718 67890 2770 67902
rect 67790 67954 67842 67966
rect 67790 67890 67842 67902
rect 68574 67954 68626 67966
rect 68574 67890 68626 67902
rect 69470 67954 69522 67966
rect 69470 67890 69522 67902
rect 70030 67954 70082 67966
rect 70030 67890 70082 67902
rect 66670 67842 66722 67854
rect 66670 67778 66722 67790
rect 67118 67842 67170 67854
rect 67118 67778 67170 67790
rect 77310 67842 77362 67854
rect 77970 67790 77982 67842
rect 78034 67790 78046 67842
rect 77310 67778 77362 67790
rect 1822 67730 1874 67742
rect 1822 67666 1874 67678
rect 2158 67618 2210 67630
rect 2158 67554 2210 67566
rect 3054 67618 3106 67630
rect 3054 67554 3106 67566
rect 67230 67618 67282 67630
rect 67230 67554 67282 67566
rect 67902 67618 67954 67630
rect 67902 67554 67954 67566
rect 68462 67618 68514 67630
rect 68462 67554 68514 67566
rect 69358 67618 69410 67630
rect 69358 67554 69410 67566
rect 77758 67618 77810 67630
rect 77758 67554 77810 67566
rect 1344 67450 78624 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 78624 67450
rect 1344 67364 78624 67398
rect 2158 67170 2210 67182
rect 2158 67106 2210 67118
rect 67566 67170 67618 67182
rect 67566 67106 67618 67118
rect 68462 67170 68514 67182
rect 68462 67106 68514 67118
rect 77758 67170 77810 67182
rect 77758 67106 77810 67118
rect 65774 67058 65826 67070
rect 1922 67006 1934 67058
rect 1986 67006 1998 67058
rect 65774 66994 65826 67006
rect 65998 67058 66050 67070
rect 65998 66994 66050 67006
rect 68238 67058 68290 67070
rect 68238 66994 68290 67006
rect 68910 67058 68962 67070
rect 68910 66994 68962 67006
rect 77310 67058 77362 67070
rect 77310 66994 77362 67006
rect 78094 67058 78146 67070
rect 78094 66994 78146 67006
rect 2606 66946 2658 66958
rect 2606 66882 2658 66894
rect 65886 66946 65938 66958
rect 65886 66882 65938 66894
rect 66222 66946 66274 66958
rect 66222 66882 66274 66894
rect 67118 66946 67170 66958
rect 67118 66882 67170 66894
rect 68350 66946 68402 66958
rect 68350 66882 68402 66894
rect 68686 66946 68738 66958
rect 68686 66882 68738 66894
rect 69358 66946 69410 66958
rect 69358 66882 69410 66894
rect 66446 66834 66498 66846
rect 66446 66770 66498 66782
rect 67006 66834 67058 66846
rect 67330 66782 67342 66834
rect 67394 66831 67406 66834
rect 67890 66831 67902 66834
rect 67394 66785 67902 66831
rect 67394 66782 67406 66785
rect 67890 66782 67902 66785
rect 67954 66782 67966 66834
rect 67006 66770 67058 66782
rect 1344 66666 78624 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 78624 66666
rect 1344 66580 78624 66614
rect 63422 66498 63474 66510
rect 63422 66434 63474 66446
rect 68350 66498 68402 66510
rect 68350 66434 68402 66446
rect 66110 66386 66162 66398
rect 66110 66322 66162 66334
rect 67006 66386 67058 66398
rect 67006 66322 67058 66334
rect 68126 66386 68178 66398
rect 68126 66322 68178 66334
rect 63310 66274 63362 66286
rect 63310 66210 63362 66222
rect 63870 66274 63922 66286
rect 63870 66210 63922 66222
rect 64878 66274 64930 66286
rect 64878 66210 64930 66222
rect 66334 66274 66386 66286
rect 66334 66210 66386 66222
rect 66894 66274 66946 66286
rect 66894 66210 66946 66222
rect 67902 66274 67954 66286
rect 67902 66210 67954 66222
rect 1822 66162 1874 66174
rect 1822 66098 1874 66110
rect 62414 66162 62466 66174
rect 62414 66098 62466 66110
rect 62526 66162 62578 66174
rect 62526 66098 62578 66110
rect 65886 66162 65938 66174
rect 65886 66098 65938 66110
rect 78094 66162 78146 66174
rect 78094 66098 78146 66110
rect 2158 66050 2210 66062
rect 2158 65986 2210 65998
rect 2606 66050 2658 66062
rect 2606 65986 2658 65998
rect 61966 66050 62018 66062
rect 61966 65986 62018 65998
rect 65662 66050 65714 66062
rect 65662 65986 65714 65998
rect 65774 66050 65826 66062
rect 65774 65986 65826 65998
rect 67678 66050 67730 66062
rect 67678 65986 67730 65998
rect 67790 66050 67842 66062
rect 67790 65986 67842 65998
rect 77310 66050 77362 66062
rect 77310 65986 77362 65998
rect 77758 66050 77810 66062
rect 77758 65986 77810 65998
rect 1344 65882 78624 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 78624 65882
rect 1344 65796 78624 65830
rect 66110 65714 66162 65726
rect 66110 65650 66162 65662
rect 2158 65602 2210 65614
rect 2158 65538 2210 65550
rect 64542 65602 64594 65614
rect 64542 65538 64594 65550
rect 65886 65602 65938 65614
rect 65886 65538 65938 65550
rect 77758 65602 77810 65614
rect 77758 65538 77810 65550
rect 61854 65490 61906 65502
rect 1922 65438 1934 65490
rect 1986 65438 1998 65490
rect 61854 65426 61906 65438
rect 65662 65490 65714 65502
rect 65662 65426 65714 65438
rect 65998 65490 66050 65502
rect 65998 65426 66050 65438
rect 68014 65490 68066 65502
rect 68014 65426 68066 65438
rect 68238 65490 68290 65502
rect 68238 65426 68290 65438
rect 68686 65490 68738 65502
rect 77970 65438 77982 65490
rect 78034 65438 78046 65490
rect 68686 65426 68738 65438
rect 2606 65378 2658 65390
rect 2606 65314 2658 65326
rect 61742 65378 61794 65390
rect 61742 65314 61794 65326
rect 62302 65378 62354 65390
rect 62302 65314 62354 65326
rect 67230 65378 67282 65390
rect 67230 65314 67282 65326
rect 68126 65378 68178 65390
rect 68126 65314 68178 65326
rect 68462 65378 68514 65390
rect 68462 65314 68514 65326
rect 77310 65378 77362 65390
rect 77310 65314 77362 65326
rect 64654 65266 64706 65278
rect 64654 65202 64706 65214
rect 65438 65266 65490 65278
rect 65438 65202 65490 65214
rect 1344 65098 78624 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 78624 65098
rect 1344 65012 78624 65046
rect 65550 64818 65602 64830
rect 65550 64754 65602 64766
rect 66446 64818 66498 64830
rect 66446 64754 66498 64766
rect 67006 64818 67058 64830
rect 67006 64754 67058 64766
rect 60734 64706 60786 64718
rect 60734 64642 60786 64654
rect 61406 64706 61458 64718
rect 61406 64642 61458 64654
rect 63534 64706 63586 64718
rect 63534 64642 63586 64654
rect 64206 64706 64258 64718
rect 64206 64642 64258 64654
rect 65774 64706 65826 64718
rect 65774 64642 65826 64654
rect 67454 64706 67506 64718
rect 67454 64642 67506 64654
rect 1822 64594 1874 64606
rect 1822 64530 1874 64542
rect 66334 64594 66386 64606
rect 66334 64530 66386 64542
rect 69358 64594 69410 64606
rect 69358 64530 69410 64542
rect 76638 64594 76690 64606
rect 76638 64530 76690 64542
rect 78094 64594 78146 64606
rect 78094 64530 78146 64542
rect 2158 64482 2210 64494
rect 2158 64418 2210 64430
rect 2606 64482 2658 64494
rect 2606 64418 2658 64430
rect 61518 64482 61570 64494
rect 61518 64418 61570 64430
rect 62078 64482 62130 64494
rect 62078 64418 62130 64430
rect 63646 64482 63698 64494
rect 63646 64418 63698 64430
rect 65102 64482 65154 64494
rect 65102 64418 65154 64430
rect 65214 64482 65266 64494
rect 65214 64418 65266 64430
rect 65326 64482 65378 64494
rect 65326 64418 65378 64430
rect 67790 64482 67842 64494
rect 67790 64418 67842 64430
rect 69694 64482 69746 64494
rect 69694 64418 69746 64430
rect 77310 64482 77362 64494
rect 77310 64418 77362 64430
rect 77758 64482 77810 64494
rect 77758 64418 77810 64430
rect 1344 64314 78624 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 78624 64314
rect 1344 64228 78624 64262
rect 65886 64146 65938 64158
rect 65886 64082 65938 64094
rect 66446 64146 66498 64158
rect 66446 64082 66498 64094
rect 67678 64146 67730 64158
rect 67678 64082 67730 64094
rect 76862 64146 76914 64158
rect 76862 64082 76914 64094
rect 2158 64034 2210 64046
rect 2158 63970 2210 63982
rect 3054 64034 3106 64046
rect 3054 63970 3106 63982
rect 3502 64034 3554 64046
rect 3502 63970 3554 63982
rect 61182 64034 61234 64046
rect 61182 63970 61234 63982
rect 62190 64034 62242 64046
rect 62190 63970 62242 63982
rect 62526 64034 62578 64046
rect 62526 63970 62578 63982
rect 63422 64034 63474 64046
rect 63422 63970 63474 63982
rect 64542 64034 64594 64046
rect 64542 63970 64594 63982
rect 68686 64034 68738 64046
rect 68686 63970 68738 63982
rect 69022 64034 69074 64046
rect 69022 63970 69074 63982
rect 77758 64034 77810 64046
rect 77758 63970 77810 63982
rect 2718 63922 2770 63934
rect 1922 63870 1934 63922
rect 1986 63870 1998 63922
rect 2718 63858 2770 63870
rect 61070 63922 61122 63934
rect 61070 63858 61122 63870
rect 61630 63922 61682 63934
rect 61630 63858 61682 63870
rect 63198 63922 63250 63934
rect 63198 63858 63250 63870
rect 64430 63922 64482 63934
rect 64430 63858 64482 63870
rect 65550 63922 65602 63934
rect 67342 63922 67394 63934
rect 66658 63870 66670 63922
rect 66722 63870 66734 63922
rect 65550 63858 65602 63870
rect 67342 63858 67394 63870
rect 76414 63922 76466 63934
rect 76414 63858 76466 63870
rect 77198 63922 77250 63934
rect 77970 63870 77982 63922
rect 78034 63870 78046 63922
rect 77198 63858 77250 63870
rect 63310 63810 63362 63822
rect 63310 63746 63362 63758
rect 63646 63810 63698 63822
rect 63646 63746 63698 63758
rect 63870 63810 63922 63822
rect 63870 63746 63922 63758
rect 1344 63530 78624 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 78624 63530
rect 1344 63444 78624 63478
rect 63758 63362 63810 63374
rect 63758 63298 63810 63310
rect 2718 63250 2770 63262
rect 2718 63186 2770 63198
rect 63534 63250 63586 63262
rect 63534 63186 63586 63198
rect 64878 63250 64930 63262
rect 64878 63186 64930 63198
rect 67006 63250 67058 63262
rect 67006 63186 67058 63198
rect 61406 63138 61458 63150
rect 61406 63074 61458 63086
rect 61966 63138 62018 63150
rect 61966 63074 62018 63086
rect 63086 63138 63138 63150
rect 63086 63074 63138 63086
rect 1822 63026 1874 63038
rect 1822 62962 1874 62974
rect 59278 63026 59330 63038
rect 59278 62962 59330 62974
rect 77310 63026 77362 63038
rect 77310 62962 77362 62974
rect 78094 63026 78146 63038
rect 78094 62962 78146 62974
rect 2158 62914 2210 62926
rect 2158 62850 2210 62862
rect 3054 62914 3106 62926
rect 3054 62850 3106 62862
rect 59390 62914 59442 62926
rect 59390 62850 59442 62862
rect 59838 62914 59890 62926
rect 59838 62850 59890 62862
rect 61518 62914 61570 62926
rect 61518 62850 61570 62862
rect 63198 62914 63250 62926
rect 63198 62850 63250 62862
rect 63310 62914 63362 62926
rect 63310 62850 63362 62862
rect 65214 62914 65266 62926
rect 65214 62850 65266 62862
rect 66110 62914 66162 62926
rect 66110 62850 66162 62862
rect 77758 62914 77810 62926
rect 77758 62850 77810 62862
rect 1344 62746 78624 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 78624 62746
rect 1344 62660 78624 62694
rect 62638 62578 62690 62590
rect 62638 62514 62690 62526
rect 62862 62578 62914 62590
rect 62862 62514 62914 62526
rect 63646 62578 63698 62590
rect 63646 62514 63698 62526
rect 68798 62578 68850 62590
rect 68798 62514 68850 62526
rect 2158 62466 2210 62478
rect 2158 62402 2210 62414
rect 77758 62466 77810 62478
rect 77758 62402 77810 62414
rect 59838 62354 59890 62366
rect 63870 62354 63922 62366
rect 1922 62302 1934 62354
rect 1986 62302 1998 62354
rect 62514 62302 62526 62354
rect 62578 62302 62590 62354
rect 63970 62302 63982 62354
rect 64034 62302 64046 62354
rect 77970 62302 77982 62354
rect 78034 62302 78046 62354
rect 59838 62290 59890 62302
rect 63870 62290 63922 62302
rect 2606 62242 2658 62254
rect 2606 62178 2658 62190
rect 59726 62242 59778 62254
rect 59726 62178 59778 62190
rect 60286 62242 60338 62254
rect 60286 62178 60338 62190
rect 62750 62242 62802 62254
rect 62750 62178 62802 62190
rect 63758 62242 63810 62254
rect 63758 62178 63810 62190
rect 64318 62242 64370 62254
rect 64318 62178 64370 62190
rect 68238 62242 68290 62254
rect 68238 62178 68290 62190
rect 68350 62242 68402 62254
rect 68350 62178 68402 62190
rect 77310 62242 77362 62254
rect 77310 62178 77362 62190
rect 62190 62130 62242 62142
rect 62190 62066 62242 62078
rect 1344 61962 78624 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 78624 61962
rect 1344 61876 78624 61910
rect 62638 61794 62690 61806
rect 62638 61730 62690 61742
rect 62750 61570 62802 61582
rect 62750 61506 62802 61518
rect 64206 61570 64258 61582
rect 64206 61506 64258 61518
rect 1822 61458 1874 61470
rect 1822 61394 1874 61406
rect 2606 61458 2658 61470
rect 2606 61394 2658 61406
rect 59726 61458 59778 61470
rect 59726 61394 59778 61406
rect 60174 61458 60226 61470
rect 60174 61394 60226 61406
rect 61406 61458 61458 61470
rect 61406 61394 61458 61406
rect 62078 61458 62130 61470
rect 62078 61394 62130 61406
rect 63310 61458 63362 61470
rect 63310 61394 63362 61406
rect 63646 61458 63698 61470
rect 63646 61394 63698 61406
rect 77310 61458 77362 61470
rect 77310 61394 77362 61406
rect 78094 61458 78146 61470
rect 78094 61394 78146 61406
rect 2158 61346 2210 61358
rect 2158 61282 2210 61294
rect 60286 61346 60338 61358
rect 60286 61282 60338 61294
rect 61518 61346 61570 61358
rect 61518 61282 61570 61294
rect 77758 61346 77810 61358
rect 77758 61282 77810 61294
rect 1344 61178 78624 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 78624 61178
rect 1344 61092 78624 61126
rect 62302 61010 62354 61022
rect 62302 60946 62354 60958
rect 65326 61010 65378 61022
rect 65326 60946 65378 60958
rect 2158 60898 2210 60910
rect 2158 60834 2210 60846
rect 59726 60898 59778 60910
rect 59726 60834 59778 60846
rect 60622 60898 60674 60910
rect 60622 60834 60674 60846
rect 62526 60898 62578 60910
rect 62526 60834 62578 60846
rect 64654 60898 64706 60910
rect 64654 60834 64706 60846
rect 77758 60898 77810 60910
rect 77758 60834 77810 60846
rect 57598 60786 57650 60798
rect 1922 60734 1934 60786
rect 1986 60734 1998 60786
rect 57598 60722 57650 60734
rect 59390 60786 59442 60798
rect 59390 60722 59442 60734
rect 60846 60786 60898 60798
rect 60846 60722 60898 60734
rect 61854 60786 61906 60798
rect 61854 60722 61906 60734
rect 63086 60786 63138 60798
rect 63086 60722 63138 60734
rect 78094 60786 78146 60798
rect 78094 60722 78146 60734
rect 2606 60674 2658 60686
rect 2606 60610 2658 60622
rect 57486 60674 57538 60686
rect 57486 60610 57538 60622
rect 58046 60674 58098 60686
rect 58046 60610 58098 60622
rect 58830 60674 58882 60686
rect 58830 60610 58882 60622
rect 60734 60674 60786 60686
rect 60734 60610 60786 60622
rect 61070 60674 61122 60686
rect 61070 60610 61122 60622
rect 62078 60674 62130 60686
rect 62078 60610 62130 60622
rect 62414 60674 62466 60686
rect 62414 60610 62466 60622
rect 77310 60674 77362 60686
rect 77310 60610 77362 60622
rect 61294 60562 61346 60574
rect 61294 60498 61346 60510
rect 64542 60562 64594 60574
rect 64542 60498 64594 60510
rect 1344 60394 78624 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 78624 60394
rect 1344 60308 78624 60342
rect 60398 60114 60450 60126
rect 60398 60050 60450 60062
rect 61518 60114 61570 60126
rect 61518 60050 61570 60062
rect 62078 60114 62130 60126
rect 62078 60050 62130 60062
rect 66670 60114 66722 60126
rect 66670 60050 66722 60062
rect 67230 60114 67282 60126
rect 67230 60050 67282 60062
rect 57374 60002 57426 60014
rect 57374 59938 57426 59950
rect 57934 60002 57986 60014
rect 57934 59938 57986 59950
rect 59950 60002 60002 60014
rect 59950 59938 60002 59950
rect 60622 60002 60674 60014
rect 60622 59938 60674 59950
rect 66558 60002 66610 60014
rect 77970 59950 77982 60002
rect 78034 59950 78046 60002
rect 66558 59938 66610 59950
rect 1822 59890 1874 59902
rect 1822 59826 1874 59838
rect 57486 59890 57538 59902
rect 57486 59826 57538 59838
rect 58718 59890 58770 59902
rect 58718 59826 58770 59838
rect 60174 59890 60226 59902
rect 60174 59826 60226 59838
rect 2158 59778 2210 59790
rect 2158 59714 2210 59726
rect 2606 59778 2658 59790
rect 2606 59714 2658 59726
rect 58830 59778 58882 59790
rect 58830 59714 58882 59726
rect 59278 59778 59330 59790
rect 59278 59714 59330 59726
rect 60062 59778 60114 59790
rect 60062 59714 60114 59726
rect 61406 59778 61458 59790
rect 61406 59714 61458 59726
rect 76638 59778 76690 59790
rect 76638 59714 76690 59726
rect 77310 59778 77362 59790
rect 77310 59714 77362 59726
rect 77758 59778 77810 59790
rect 77758 59714 77810 59726
rect 1344 59610 78624 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 78624 59610
rect 1344 59524 78624 59558
rect 59838 59442 59890 59454
rect 59838 59378 59890 59390
rect 61070 59442 61122 59454
rect 61070 59378 61122 59390
rect 2158 59330 2210 59342
rect 2158 59266 2210 59278
rect 3054 59330 3106 59342
rect 3054 59266 3106 59278
rect 59614 59330 59666 59342
rect 59614 59266 59666 59278
rect 76862 59330 76914 59342
rect 76862 59266 76914 59278
rect 77758 59330 77810 59342
rect 77758 59266 77810 59278
rect 2718 59218 2770 59230
rect 1922 59166 1934 59218
rect 1986 59166 1998 59218
rect 2718 59154 2770 59166
rect 3502 59218 3554 59230
rect 3502 59154 3554 59166
rect 60286 59218 60338 59230
rect 77198 59218 77250 59230
rect 61282 59166 61294 59218
rect 61346 59166 61358 59218
rect 60286 59154 60338 59166
rect 77198 59154 77250 59166
rect 78094 59218 78146 59230
rect 78094 59154 78146 59166
rect 59726 59106 59778 59118
rect 59726 59042 59778 59054
rect 60062 59106 60114 59118
rect 60062 59042 60114 59054
rect 61854 59106 61906 59118
rect 61854 59042 61906 59054
rect 76414 59106 76466 59118
rect 76414 59042 76466 59054
rect 1344 58826 78624 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 78624 58826
rect 1344 58740 78624 58774
rect 2718 58546 2770 58558
rect 2718 58482 2770 58494
rect 59390 58546 59442 58558
rect 59390 58482 59442 58494
rect 60398 58546 60450 58558
rect 60398 58482 60450 58494
rect 56142 58434 56194 58446
rect 56142 58370 56194 58382
rect 56702 58434 56754 58446
rect 56702 58370 56754 58382
rect 58494 58434 58546 58446
rect 58494 58370 58546 58382
rect 59950 58434 60002 58446
rect 77970 58382 77982 58434
rect 78034 58382 78046 58434
rect 59950 58370 60002 58382
rect 1822 58322 1874 58334
rect 1822 58258 1874 58270
rect 57262 58322 57314 58334
rect 57262 58258 57314 58270
rect 57822 58322 57874 58334
rect 57822 58258 57874 58270
rect 77310 58322 77362 58334
rect 77310 58258 77362 58270
rect 2158 58210 2210 58222
rect 2158 58146 2210 58158
rect 3054 58210 3106 58222
rect 3054 58146 3106 58158
rect 56254 58210 56306 58222
rect 56254 58146 56306 58158
rect 57374 58210 57426 58222
rect 57374 58146 57426 58158
rect 58606 58210 58658 58222
rect 58606 58146 58658 58158
rect 59278 58210 59330 58222
rect 59278 58146 59330 58158
rect 77758 58210 77810 58222
rect 77758 58146 77810 58158
rect 1344 58042 78624 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 78624 58042
rect 1344 57956 78624 57990
rect 57598 57874 57650 57886
rect 57598 57810 57650 57822
rect 59502 57874 59554 57886
rect 59502 57810 59554 57822
rect 2158 57762 2210 57774
rect 2158 57698 2210 57710
rect 77758 57762 77810 57774
rect 77758 57698 77810 57710
rect 55134 57650 55186 57662
rect 1922 57598 1934 57650
rect 1986 57598 1998 57650
rect 55134 57586 55186 57598
rect 57822 57650 57874 57662
rect 57822 57586 57874 57598
rect 58830 57650 58882 57662
rect 58830 57586 58882 57598
rect 59278 57650 59330 57662
rect 59278 57586 59330 57598
rect 62750 57650 62802 57662
rect 62750 57586 62802 57598
rect 63198 57650 63250 57662
rect 63198 57586 63250 57598
rect 78094 57650 78146 57662
rect 78094 57586 78146 57598
rect 2606 57538 2658 57550
rect 2606 57474 2658 57486
rect 55022 57538 55074 57550
rect 55022 57474 55074 57486
rect 55582 57538 55634 57550
rect 55582 57474 55634 57486
rect 57710 57538 57762 57550
rect 57710 57474 57762 57486
rect 58046 57538 58098 57550
rect 58046 57474 58098 57486
rect 59054 57538 59106 57550
rect 59054 57474 59106 57486
rect 59390 57538 59442 57550
rect 59390 57474 59442 57486
rect 77310 57538 77362 57550
rect 77310 57474 77362 57486
rect 58270 57426 58322 57438
rect 58270 57362 58322 57374
rect 62638 57426 62690 57438
rect 62638 57362 62690 57374
rect 1344 57258 78624 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 78624 57258
rect 1344 57172 78624 57206
rect 58494 57090 58546 57102
rect 58494 57026 58546 57038
rect 59166 56978 59218 56990
rect 59166 56914 59218 56926
rect 57822 56866 57874 56878
rect 57822 56802 57874 56814
rect 58046 56866 58098 56878
rect 58146 56814 58158 56866
rect 58210 56814 58222 56866
rect 77970 56814 77982 56866
rect 78034 56814 78046 56866
rect 58046 56802 58098 56814
rect 1822 56754 1874 56766
rect 1822 56690 1874 56702
rect 56254 56754 56306 56766
rect 56254 56690 56306 56702
rect 56702 56754 56754 56766
rect 56702 56690 56754 56702
rect 2158 56642 2210 56654
rect 2158 56578 2210 56590
rect 2606 56642 2658 56654
rect 2606 56578 2658 56590
rect 56814 56642 56866 56654
rect 56814 56578 56866 56590
rect 57934 56642 57986 56654
rect 57934 56578 57986 56590
rect 59054 56642 59106 56654
rect 59054 56578 59106 56590
rect 59726 56642 59778 56654
rect 59726 56578 59778 56590
rect 77310 56642 77362 56654
rect 77310 56578 77362 56590
rect 77758 56642 77810 56654
rect 77758 56578 77810 56590
rect 1344 56474 78624 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 78624 56474
rect 1344 56388 78624 56422
rect 56590 56306 56642 56318
rect 56590 56242 56642 56254
rect 57822 56306 57874 56318
rect 57822 56242 57874 56254
rect 2158 56194 2210 56206
rect 2158 56130 2210 56142
rect 57598 56194 57650 56206
rect 57598 56130 57650 56142
rect 77758 56194 77810 56206
rect 77758 56130 77810 56142
rect 52222 56082 52274 56094
rect 1922 56030 1934 56082
rect 1986 56030 1998 56082
rect 52222 56018 52274 56030
rect 55358 56082 55410 56094
rect 55358 56018 55410 56030
rect 55582 56082 55634 56094
rect 56030 56082 56082 56094
rect 55682 56030 55694 56082
rect 55746 56030 55758 56082
rect 55582 56018 55634 56030
rect 56030 56018 56082 56030
rect 58270 56082 58322 56094
rect 58270 56018 58322 56030
rect 78094 56082 78146 56094
rect 78094 56018 78146 56030
rect 2606 55970 2658 55982
rect 2606 55906 2658 55918
rect 52110 55970 52162 55982
rect 52110 55906 52162 55918
rect 52670 55970 52722 55982
rect 52670 55906 52722 55918
rect 54686 55970 54738 55982
rect 54686 55906 54738 55918
rect 55470 55970 55522 55982
rect 55470 55906 55522 55918
rect 56702 55970 56754 55982
rect 56702 55906 56754 55918
rect 57710 55970 57762 55982
rect 57710 55906 57762 55918
rect 58046 55970 58098 55982
rect 58046 55906 58098 55918
rect 58718 55970 58770 55982
rect 58718 55906 58770 55918
rect 77310 55970 77362 55982
rect 77310 55906 77362 55918
rect 1344 55690 78624 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 78624 55690
rect 1344 55604 78624 55638
rect 57586 55470 57598 55522
rect 57650 55519 57662 55522
rect 57810 55519 57822 55522
rect 57650 55473 57822 55519
rect 57650 55470 57662 55473
rect 57810 55470 57822 55473
rect 57874 55470 57886 55522
rect 50318 55410 50370 55422
rect 50318 55346 50370 55358
rect 50878 55410 50930 55422
rect 50878 55346 50930 55358
rect 55582 55410 55634 55422
rect 55582 55346 55634 55358
rect 55134 55298 55186 55310
rect 54114 55246 54126 55298
rect 54178 55246 54190 55298
rect 55134 55234 55186 55246
rect 55806 55298 55858 55310
rect 77970 55246 77982 55298
rect 78034 55246 78046 55298
rect 55806 55234 55858 55246
rect 1822 55186 1874 55198
rect 1822 55122 1874 55134
rect 54350 55186 54402 55198
rect 54350 55122 54402 55134
rect 56926 55186 56978 55198
rect 56926 55122 56978 55134
rect 57262 55186 57314 55198
rect 57262 55122 57314 55134
rect 2158 55074 2210 55086
rect 2158 55010 2210 55022
rect 2606 55074 2658 55086
rect 2606 55010 2658 55022
rect 50430 55074 50482 55086
rect 50430 55010 50482 55022
rect 52446 55074 52498 55086
rect 52446 55010 52498 55022
rect 53566 55074 53618 55086
rect 53566 55010 53618 55022
rect 55246 55074 55298 55086
rect 55246 55010 55298 55022
rect 55358 55074 55410 55086
rect 55358 55010 55410 55022
rect 56254 55074 56306 55086
rect 56254 55010 56306 55022
rect 57710 55074 57762 55086
rect 57710 55010 57762 55022
rect 76638 55074 76690 55086
rect 76638 55010 76690 55022
rect 77310 55074 77362 55086
rect 77310 55010 77362 55022
rect 77758 55074 77810 55086
rect 77758 55010 77810 55022
rect 1344 54906 78624 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 78624 54906
rect 1344 54820 78624 54854
rect 56478 54738 56530 54750
rect 56478 54674 56530 54686
rect 57822 54738 57874 54750
rect 57822 54674 57874 54686
rect 76862 54738 76914 54750
rect 76862 54674 76914 54686
rect 2158 54626 2210 54638
rect 2158 54562 2210 54574
rect 3054 54626 3106 54638
rect 3054 54562 3106 54574
rect 51662 54626 51714 54638
rect 51662 54562 51714 54574
rect 52110 54626 52162 54638
rect 52110 54562 52162 54574
rect 52782 54626 52834 54638
rect 52782 54562 52834 54574
rect 53790 54626 53842 54638
rect 53790 54562 53842 54574
rect 55918 54626 55970 54638
rect 55918 54562 55970 54574
rect 56590 54626 56642 54638
rect 56590 54562 56642 54574
rect 77758 54626 77810 54638
rect 77758 54562 77810 54574
rect 2718 54514 2770 54526
rect 1922 54462 1934 54514
rect 1986 54462 1998 54514
rect 2718 54450 2770 54462
rect 3502 54514 3554 54526
rect 3502 54450 3554 54462
rect 52894 54514 52946 54526
rect 52894 54450 52946 54462
rect 54574 54514 54626 54526
rect 54574 54450 54626 54462
rect 54798 54514 54850 54526
rect 54798 54450 54850 54462
rect 55022 54514 55074 54526
rect 55022 54450 55074 54462
rect 57486 54514 57538 54526
rect 57486 54450 57538 54462
rect 77198 54514 77250 54526
rect 77198 54450 77250 54462
rect 78094 54514 78146 54526
rect 78094 54450 78146 54462
rect 54686 54402 54738 54414
rect 54686 54338 54738 54350
rect 76414 54402 76466 54414
rect 76414 54338 76466 54350
rect 52222 54290 52274 54302
rect 52222 54226 52274 54238
rect 53902 54290 53954 54302
rect 53902 54226 53954 54238
rect 55246 54290 55298 54302
rect 55246 54226 55298 54238
rect 55806 54290 55858 54302
rect 55806 54226 55858 54238
rect 1344 54122 78624 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 78624 54122
rect 1344 54036 78624 54070
rect 54238 53954 54290 53966
rect 57138 53902 57150 53954
rect 57202 53951 57214 53954
rect 57474 53951 57486 53954
rect 57202 53905 57486 53951
rect 57202 53902 57214 53905
rect 57474 53902 57486 53905
rect 57538 53902 57550 53954
rect 54238 53890 54290 53902
rect 2718 53842 2770 53854
rect 2718 53778 2770 53790
rect 54462 53730 54514 53742
rect 54462 53666 54514 53678
rect 54686 53730 54738 53742
rect 54686 53666 54738 53678
rect 54910 53730 54962 53742
rect 54910 53666 54962 53678
rect 55918 53730 55970 53742
rect 55918 53666 55970 53678
rect 56926 53730 56978 53742
rect 56926 53666 56978 53678
rect 57486 53730 57538 53742
rect 57486 53666 57538 53678
rect 1822 53618 1874 53630
rect 1822 53554 1874 53566
rect 2158 53618 2210 53630
rect 2158 53554 2210 53566
rect 52782 53618 52834 53630
rect 52782 53554 52834 53566
rect 53454 53618 53506 53630
rect 53454 53554 53506 53566
rect 55582 53618 55634 53630
rect 55582 53554 55634 53566
rect 78094 53618 78146 53630
rect 78094 53554 78146 53566
rect 3054 53506 3106 53518
rect 3054 53442 3106 53454
rect 52110 53506 52162 53518
rect 52110 53442 52162 53454
rect 53566 53506 53618 53518
rect 53566 53442 53618 53454
rect 54798 53506 54850 53518
rect 54798 53442 54850 53454
rect 77310 53506 77362 53518
rect 77310 53442 77362 53454
rect 77758 53506 77810 53518
rect 77758 53442 77810 53454
rect 1344 53338 78624 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 78624 53338
rect 1344 53252 78624 53286
rect 47742 53170 47794 53182
rect 47742 53106 47794 53118
rect 52670 53170 52722 53182
rect 52670 53106 52722 53118
rect 57822 53170 57874 53182
rect 57822 53106 57874 53118
rect 2158 53058 2210 53070
rect 2158 52994 2210 53006
rect 48302 53058 48354 53070
rect 48302 52994 48354 53006
rect 50318 53058 50370 53070
rect 50318 52994 50370 53006
rect 51886 53058 51938 53070
rect 51886 52994 51938 53006
rect 54350 53058 54402 53070
rect 54350 52994 54402 53006
rect 56702 53058 56754 53070
rect 56702 52994 56754 53006
rect 77758 53058 77810 53070
rect 77758 52994 77810 53006
rect 48414 52946 48466 52958
rect 52894 52946 52946 52958
rect 1922 52894 1934 52946
rect 1986 52894 1998 52946
rect 51650 52894 51662 52946
rect 51714 52894 51726 52946
rect 48414 52882 48466 52894
rect 52894 52882 52946 52894
rect 53902 52946 53954 52958
rect 53902 52882 53954 52894
rect 54574 52946 54626 52958
rect 54574 52882 54626 52894
rect 57486 52946 57538 52958
rect 77970 52894 77982 52946
rect 78034 52894 78046 52946
rect 57486 52882 57538 52894
rect 2606 52834 2658 52846
rect 2606 52770 2658 52782
rect 50206 52834 50258 52846
rect 50206 52770 50258 52782
rect 50766 52834 50818 52846
rect 50766 52770 50818 52782
rect 52782 52834 52834 52846
rect 52782 52770 52834 52782
rect 53118 52834 53170 52846
rect 53118 52770 53170 52782
rect 54126 52834 54178 52846
rect 54126 52770 54178 52782
rect 54462 52834 54514 52846
rect 54462 52770 54514 52782
rect 77310 52834 77362 52846
rect 77310 52770 77362 52782
rect 53342 52722 53394 52734
rect 53342 52658 53394 52670
rect 56590 52722 56642 52734
rect 56590 52658 56642 52670
rect 1344 52554 78624 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 78624 52554
rect 1344 52468 78624 52502
rect 52670 52386 52722 52398
rect 52670 52322 52722 52334
rect 60286 52386 60338 52398
rect 60286 52322 60338 52334
rect 46958 52274 47010 52286
rect 46958 52210 47010 52222
rect 47518 52274 47570 52286
rect 47518 52210 47570 52222
rect 48750 52274 48802 52286
rect 48750 52210 48802 52222
rect 49310 52274 49362 52286
rect 49310 52210 49362 52222
rect 51326 52274 51378 52286
rect 51326 52210 51378 52222
rect 52446 52274 52498 52286
rect 52446 52210 52498 52222
rect 59166 52274 59218 52286
rect 59166 52210 59218 52222
rect 60398 52274 60450 52286
rect 60398 52210 60450 52222
rect 61406 52274 61458 52286
rect 61406 52210 61458 52222
rect 50878 52162 50930 52174
rect 56814 52162 56866 52174
rect 56242 52110 56254 52162
rect 56306 52110 56318 52162
rect 50878 52098 50930 52110
rect 56814 52098 56866 52110
rect 57262 52162 57314 52174
rect 57262 52098 57314 52110
rect 59278 52162 59330 52174
rect 59278 52098 59330 52110
rect 59838 52162 59890 52174
rect 59838 52098 59890 52110
rect 1822 52050 1874 52062
rect 1822 51986 1874 51998
rect 2606 52050 2658 52062
rect 2606 51986 2658 51998
rect 47070 52050 47122 52062
rect 47070 51986 47122 51998
rect 52222 52050 52274 52062
rect 52222 51986 52274 51998
rect 56030 52050 56082 52062
rect 56030 51986 56082 51998
rect 78094 52050 78146 52062
rect 78094 51986 78146 51998
rect 2158 51938 2210 51950
rect 2158 51874 2210 51886
rect 48862 51938 48914 51950
rect 48862 51874 48914 51886
rect 50542 51938 50594 51950
rect 50542 51874 50594 51886
rect 51998 51938 52050 51950
rect 51998 51874 52050 51886
rect 52110 51938 52162 51950
rect 52110 51874 52162 51886
rect 77310 51938 77362 51950
rect 77310 51874 77362 51886
rect 77758 51938 77810 51950
rect 77758 51874 77810 51886
rect 1344 51770 78624 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 78624 51770
rect 1344 51684 78624 51718
rect 51886 51602 51938 51614
rect 51886 51538 51938 51550
rect 53342 51602 53394 51614
rect 53342 51538 53394 51550
rect 56142 51602 56194 51614
rect 56142 51538 56194 51550
rect 57822 51602 57874 51614
rect 57822 51538 57874 51550
rect 2158 51490 2210 51502
rect 2158 51426 2210 51438
rect 52110 51490 52162 51502
rect 52110 51426 52162 51438
rect 53678 51490 53730 51502
rect 53678 51426 53730 51438
rect 77758 51490 77810 51502
rect 77758 51426 77810 51438
rect 52334 51378 52386 51390
rect 1922 51326 1934 51378
rect 1986 51326 1998 51378
rect 52334 51314 52386 51326
rect 52558 51378 52610 51390
rect 57486 51378 57538 51390
rect 56354 51326 56366 51378
rect 56418 51326 56430 51378
rect 77970 51326 77982 51378
rect 78034 51326 78046 51378
rect 52558 51314 52610 51326
rect 57486 51314 57538 51326
rect 2606 51266 2658 51278
rect 2606 51202 2658 51214
rect 51998 51266 52050 51278
rect 51998 51202 52050 51214
rect 55582 51266 55634 51278
rect 55582 51202 55634 51214
rect 77310 51266 77362 51278
rect 77310 51202 77362 51214
rect 1344 50986 78624 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 78624 50986
rect 1344 50900 78624 50934
rect 49198 50706 49250 50718
rect 49198 50642 49250 50654
rect 49646 50706 49698 50718
rect 49646 50642 49698 50654
rect 57150 50706 57202 50718
rect 57150 50642 57202 50654
rect 68686 50706 68738 50718
rect 68686 50642 68738 50654
rect 69358 50706 69410 50718
rect 69358 50642 69410 50654
rect 70030 50706 70082 50718
rect 70030 50642 70082 50654
rect 70702 50706 70754 50718
rect 70702 50642 70754 50654
rect 77310 50706 77362 50718
rect 77310 50642 77362 50654
rect 51102 50594 51154 50606
rect 50754 50542 50766 50594
rect 50818 50542 50830 50594
rect 51102 50530 51154 50542
rect 51662 50594 51714 50606
rect 51662 50530 51714 50542
rect 51774 50594 51826 50606
rect 51774 50530 51826 50542
rect 52334 50594 52386 50606
rect 53666 50542 53678 50594
rect 53730 50542 53742 50594
rect 52334 50530 52386 50542
rect 1822 50482 1874 50494
rect 1822 50418 1874 50430
rect 3054 50482 3106 50494
rect 3054 50418 3106 50430
rect 49758 50482 49810 50494
rect 49758 50418 49810 50430
rect 50654 50482 50706 50494
rect 50654 50418 50706 50430
rect 78094 50482 78146 50494
rect 78094 50418 78146 50430
rect 2158 50370 2210 50382
rect 2158 50306 2210 50318
rect 2718 50370 2770 50382
rect 2718 50306 2770 50318
rect 50430 50370 50482 50382
rect 50430 50306 50482 50318
rect 50542 50370 50594 50382
rect 50542 50306 50594 50318
rect 53454 50370 53506 50382
rect 53454 50306 53506 50318
rect 69470 50370 69522 50382
rect 69470 50306 69522 50318
rect 70142 50370 70194 50382
rect 70142 50306 70194 50318
rect 77758 50370 77810 50382
rect 77758 50306 77810 50318
rect 1344 50202 78624 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 78624 50202
rect 1344 50116 78624 50150
rect 46622 50034 46674 50046
rect 46622 49970 46674 49982
rect 50206 50034 50258 50046
rect 50206 49970 50258 49982
rect 50990 50034 51042 50046
rect 50990 49970 51042 49982
rect 51214 50034 51266 50046
rect 51214 49970 51266 49982
rect 69806 50034 69858 50046
rect 69806 49970 69858 49982
rect 2158 49922 2210 49934
rect 2158 49858 2210 49870
rect 3054 49922 3106 49934
rect 3054 49858 3106 49870
rect 52334 49922 52386 49934
rect 52334 49858 52386 49870
rect 77758 49922 77810 49934
rect 77758 49858 77810 49870
rect 1822 49810 1874 49822
rect 1822 49746 1874 49758
rect 2718 49810 2770 49822
rect 2718 49746 2770 49758
rect 49982 49810 50034 49822
rect 49982 49746 50034 49758
rect 68910 49810 68962 49822
rect 68910 49746 68962 49758
rect 69582 49810 69634 49822
rect 69582 49746 69634 49758
rect 70254 49810 70306 49822
rect 77970 49758 77982 49810
rect 78034 49758 78046 49810
rect 70254 49746 70306 49758
rect 3502 49698 3554 49710
rect 3502 49634 3554 49646
rect 46510 49698 46562 49710
rect 46510 49634 46562 49646
rect 47070 49698 47122 49710
rect 47070 49634 47122 49646
rect 49758 49698 49810 49710
rect 49758 49634 49810 49646
rect 50094 49698 50146 49710
rect 50094 49634 50146 49646
rect 51102 49698 51154 49710
rect 51102 49634 51154 49646
rect 51438 49698 51490 49710
rect 51438 49634 51490 49646
rect 52782 49698 52834 49710
rect 52782 49634 52834 49646
rect 69694 49698 69746 49710
rect 69694 49634 69746 49646
rect 70030 49698 70082 49710
rect 70030 49634 70082 49646
rect 70702 49698 70754 49710
rect 70702 49634 70754 49646
rect 77310 49698 77362 49710
rect 77310 49634 77362 49646
rect 49534 49586 49586 49598
rect 49534 49522 49586 49534
rect 51662 49586 51714 49598
rect 51662 49522 51714 49534
rect 52222 49586 52274 49598
rect 52222 49522 52274 49534
rect 1344 49418 78624 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 78624 49418
rect 1344 49332 78624 49366
rect 48078 49250 48130 49262
rect 48078 49186 48130 49198
rect 47966 49138 48018 49150
rect 47966 49074 48018 49086
rect 48526 49138 48578 49150
rect 48526 49074 48578 49086
rect 49646 49138 49698 49150
rect 49646 49074 49698 49086
rect 68014 49138 68066 49150
rect 68014 49074 68066 49086
rect 68574 49138 68626 49150
rect 68574 49074 68626 49086
rect 69582 49138 69634 49150
rect 69582 49074 69634 49086
rect 70702 49138 70754 49150
rect 70702 49074 70754 49086
rect 49198 49026 49250 49038
rect 3042 48974 3054 49026
rect 3106 48974 3118 49026
rect 49198 48962 49250 48974
rect 49870 49026 49922 49038
rect 49870 48962 49922 48974
rect 50430 49026 50482 49038
rect 50430 48962 50482 48974
rect 69358 49026 69410 49038
rect 69358 48962 69410 48974
rect 50542 48914 50594 48926
rect 2146 48862 2158 48914
rect 2210 48862 2222 48914
rect 50542 48850 50594 48862
rect 78094 48914 78146 48926
rect 78094 48850 78146 48862
rect 3502 48802 3554 48814
rect 3502 48738 3554 48750
rect 49310 48802 49362 48814
rect 49310 48738 49362 48750
rect 49422 48802 49474 48814
rect 49422 48738 49474 48750
rect 51102 48802 51154 48814
rect 51102 48738 51154 48750
rect 68126 48802 68178 48814
rect 68126 48738 68178 48750
rect 69806 48802 69858 48814
rect 69806 48738 69858 48750
rect 69918 48802 69970 48814
rect 69918 48738 69970 48750
rect 70030 48802 70082 48814
rect 70030 48738 70082 48750
rect 76638 48802 76690 48814
rect 76638 48738 76690 48750
rect 77310 48802 77362 48814
rect 77310 48738 77362 48750
rect 77758 48802 77810 48814
rect 77758 48738 77810 48750
rect 1344 48634 78624 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 78624 48634
rect 1344 48548 78624 48582
rect 48526 48466 48578 48478
rect 48526 48402 48578 48414
rect 49758 48466 49810 48478
rect 49758 48402 49810 48414
rect 50318 48466 50370 48478
rect 50318 48402 50370 48414
rect 68910 48466 68962 48478
rect 68910 48402 68962 48414
rect 69358 48466 69410 48478
rect 69358 48402 69410 48414
rect 49870 48354 49922 48366
rect 49870 48290 49922 48302
rect 68798 48354 68850 48366
rect 68798 48290 68850 48302
rect 3042 48190 3054 48242
rect 3106 48190 3118 48242
rect 75058 48190 75070 48242
rect 75122 48190 75134 48242
rect 76962 48190 76974 48242
rect 77026 48190 77038 48242
rect 3614 48130 3666 48142
rect 2034 48078 2046 48130
rect 2098 48078 2110 48130
rect 3614 48066 3666 48078
rect 47294 48130 47346 48142
rect 47294 48066 47346 48078
rect 47854 48130 47906 48142
rect 47854 48066 47906 48078
rect 48414 48130 48466 48142
rect 48414 48066 48466 48078
rect 69918 48130 69970 48142
rect 69918 48066 69970 48078
rect 74622 48130 74674 48142
rect 76066 48078 76078 48130
rect 76130 48078 76142 48130
rect 77858 48078 77870 48130
rect 77922 48078 77934 48130
rect 74622 48066 74674 48078
rect 1344 47850 78624 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 78624 47850
rect 1344 47764 78624 47798
rect 3042 47406 3054 47458
rect 3106 47406 3118 47458
rect 47518 47346 47570 47358
rect 2146 47294 2158 47346
rect 2210 47294 2222 47346
rect 47518 47282 47570 47294
rect 48190 47346 48242 47358
rect 48190 47282 48242 47294
rect 48974 47346 49026 47358
rect 48974 47282 49026 47294
rect 3502 47234 3554 47246
rect 3502 47170 3554 47182
rect 47182 47234 47234 47246
rect 47182 47170 47234 47182
rect 48526 47234 48578 47246
rect 48526 47170 48578 47182
rect 76638 47234 76690 47246
rect 76638 47170 76690 47182
rect 1344 47066 78624 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 78624 47066
rect 1344 46980 78624 47014
rect 46510 46786 46562 46798
rect 46510 46722 46562 46734
rect 47854 46786 47906 46798
rect 47854 46722 47906 46734
rect 46846 46674 46898 46686
rect 3042 46622 3054 46674
rect 3106 46622 3118 46674
rect 47618 46622 47630 46674
rect 47682 46622 47694 46674
rect 75058 46622 75070 46674
rect 75122 46622 75134 46674
rect 77074 46622 77086 46674
rect 77138 46622 77150 46674
rect 46846 46610 46898 46622
rect 3614 46562 3666 46574
rect 2034 46510 2046 46562
rect 2098 46510 2110 46562
rect 3614 46498 3666 46510
rect 46062 46562 46114 46574
rect 46062 46498 46114 46510
rect 48302 46562 48354 46574
rect 48302 46498 48354 46510
rect 74622 46562 74674 46574
rect 76066 46510 76078 46562
rect 76130 46510 76142 46562
rect 77746 46510 77758 46562
rect 77810 46510 77822 46562
rect 74622 46498 74674 46510
rect 1344 46282 78624 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 78624 46282
rect 1344 46196 78624 46230
rect 47742 45890 47794 45902
rect 3042 45838 3054 45890
rect 3106 45838 3118 45890
rect 47742 45826 47794 45838
rect 48078 45890 48130 45902
rect 75282 45838 75294 45890
rect 75346 45838 75358 45890
rect 48078 45826 48130 45838
rect 46174 45778 46226 45790
rect 2146 45726 2158 45778
rect 2210 45726 2222 45778
rect 46174 45714 46226 45726
rect 46846 45778 46898 45790
rect 46846 45714 46898 45726
rect 47182 45778 47234 45790
rect 76178 45726 76190 45778
rect 76242 45726 76254 45778
rect 47182 45714 47234 45726
rect 3502 45666 3554 45678
rect 3502 45602 3554 45614
rect 45838 45666 45890 45678
rect 45838 45602 45890 45614
rect 74734 45666 74786 45678
rect 74734 45602 74786 45614
rect 1344 45498 78624 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 78624 45498
rect 1344 45412 78624 45446
rect 44382 45330 44434 45342
rect 44382 45266 44434 45278
rect 46510 45330 46562 45342
rect 46510 45266 46562 45278
rect 45278 45218 45330 45230
rect 45278 45154 45330 45166
rect 43934 45106 43986 45118
rect 45614 45106 45666 45118
rect 3042 45054 3054 45106
rect 3106 45054 3118 45106
rect 44594 45054 44606 45106
rect 44658 45054 44670 45106
rect 46274 45054 46286 45106
rect 46338 45054 46350 45106
rect 75058 45054 75070 45106
rect 75122 45054 75134 45106
rect 76850 45054 76862 45106
rect 76914 45054 76926 45106
rect 43934 45042 43986 45054
rect 45614 45042 45666 45054
rect 3614 44994 3666 45006
rect 2034 44942 2046 44994
rect 2098 44942 2110 44994
rect 3614 44930 3666 44942
rect 46958 44994 47010 45006
rect 46958 44930 47010 44942
rect 47406 44994 47458 45006
rect 47406 44930 47458 44942
rect 74622 44994 74674 45006
rect 76066 44942 76078 44994
rect 76130 44942 76142 44994
rect 77858 44942 77870 44994
rect 77922 44942 77934 44994
rect 74622 44930 74674 44942
rect 1344 44714 78624 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 78624 44714
rect 1344 44628 78624 44662
rect 46398 44322 46450 44334
rect 3042 44270 3054 44322
rect 3106 44270 3118 44322
rect 46398 44258 46450 44270
rect 43710 44210 43762 44222
rect 2146 44158 2158 44210
rect 2210 44158 2222 44210
rect 43710 44146 43762 44158
rect 44046 44210 44098 44222
rect 44046 44146 44098 44158
rect 44606 44210 44658 44222
rect 44606 44146 44658 44158
rect 45502 44210 45554 44222
rect 45502 44146 45554 44158
rect 45838 44210 45890 44222
rect 45838 44146 45890 44158
rect 3502 44098 3554 44110
rect 3502 44034 3554 44046
rect 46734 44098 46786 44110
rect 46734 44034 46786 44046
rect 76526 44098 76578 44110
rect 76526 44034 76578 44046
rect 1344 43930 78624 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 78624 43930
rect 1344 43844 78624 43878
rect 42926 43762 42978 43774
rect 42926 43698 42978 43710
rect 44382 43762 44434 43774
rect 44382 43698 44434 43710
rect 43262 43538 43314 43550
rect 3042 43486 3054 43538
rect 3106 43486 3118 43538
rect 44146 43486 44158 43538
rect 44210 43486 44222 43538
rect 76850 43486 76862 43538
rect 76914 43486 76926 43538
rect 43262 43474 43314 43486
rect 3614 43426 3666 43438
rect 2034 43374 2046 43426
rect 2098 43374 2110 43426
rect 3614 43362 3666 43374
rect 42478 43426 42530 43438
rect 42478 43362 42530 43374
rect 44830 43426 44882 43438
rect 44830 43362 44882 43374
rect 45278 43426 45330 43438
rect 45278 43362 45330 43374
rect 46062 43426 46114 43438
rect 46062 43362 46114 43374
rect 76414 43426 76466 43438
rect 77858 43374 77870 43426
rect 77922 43374 77934 43426
rect 76414 43362 76466 43374
rect 1344 43146 78624 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 78624 43146
rect 1344 43060 78624 43094
rect 41918 42754 41970 42766
rect 43374 42754 43426 42766
rect 3042 42702 3054 42754
rect 3106 42702 3118 42754
rect 42578 42702 42590 42754
rect 42642 42702 42654 42754
rect 41918 42690 41970 42702
rect 43374 42690 43426 42702
rect 42366 42642 42418 42654
rect 2146 42590 2158 42642
rect 2210 42590 2222 42642
rect 42366 42578 42418 42590
rect 3502 42530 3554 42542
rect 3502 42466 3554 42478
rect 43710 42530 43762 42542
rect 43710 42466 43762 42478
rect 44158 42530 44210 42542
rect 44158 42466 44210 42478
rect 1344 42362 78624 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 78624 42362
rect 1344 42276 78624 42310
rect 41694 42194 41746 42206
rect 41694 42130 41746 42142
rect 43038 42082 43090 42094
rect 43038 42018 43090 42030
rect 42030 41970 42082 41982
rect 3042 41918 3054 41970
rect 3106 41918 3118 41970
rect 42802 41918 42814 41970
rect 42866 41918 42878 41970
rect 75058 41918 75070 41970
rect 75122 41918 75134 41970
rect 76850 41918 76862 41970
rect 76914 41918 76926 41970
rect 77746 41918 77758 41970
rect 77810 41918 77822 41970
rect 42030 41906 42082 41918
rect 3614 41858 3666 41870
rect 2034 41806 2046 41858
rect 2098 41806 2110 41858
rect 3614 41794 3666 41806
rect 43486 41858 43538 41870
rect 43486 41794 43538 41806
rect 43934 41858 43986 41870
rect 43934 41794 43986 41806
rect 74622 41858 74674 41870
rect 76066 41806 76078 41858
rect 76130 41806 76142 41858
rect 74622 41794 74674 41806
rect 1344 41578 78624 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 78624 41578
rect 1344 41492 78624 41526
rect 3042 41134 3054 41186
rect 3106 41134 3118 41186
rect 42130 41134 42142 41186
rect 42194 41134 42206 41186
rect 41022 41074 41074 41086
rect 2146 41022 2158 41074
rect 2210 41022 2222 41074
rect 41022 41010 41074 41022
rect 41358 41074 41410 41086
rect 41358 41010 41410 41022
rect 42366 41074 42418 41086
rect 42366 41010 42418 41022
rect 3502 40962 3554 40974
rect 3502 40898 3554 40910
rect 40014 40962 40066 40974
rect 40014 40898 40066 40910
rect 40574 40962 40626 40974
rect 40574 40898 40626 40910
rect 42814 40962 42866 40974
rect 42814 40898 42866 40910
rect 76638 40962 76690 40974
rect 76638 40898 76690 40910
rect 1344 40794 78624 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 78624 40794
rect 1344 40708 78624 40742
rect 40238 40626 40290 40638
rect 40238 40562 40290 40574
rect 39342 40514 39394 40526
rect 39342 40450 39394 40462
rect 41918 40514 41970 40526
rect 77746 40462 77758 40514
rect 77810 40462 77822 40514
rect 41918 40450 41970 40462
rect 3614 40402 3666 40414
rect 3042 40350 3054 40402
rect 3106 40350 3118 40402
rect 3614 40338 3666 40350
rect 39678 40402 39730 40414
rect 39678 40338 39730 40350
rect 40574 40402 40626 40414
rect 40574 40338 40626 40350
rect 41582 40402 41634 40414
rect 41582 40338 41634 40350
rect 42366 40402 42418 40414
rect 42366 40338 42418 40350
rect 74622 40402 74674 40414
rect 75058 40350 75070 40402
rect 75122 40350 75134 40402
rect 75954 40350 75966 40402
rect 76018 40350 76030 40402
rect 76850 40350 76862 40402
rect 76914 40350 76926 40402
rect 74622 40338 74674 40350
rect 38894 40290 38946 40302
rect 2034 40238 2046 40290
rect 2098 40238 2110 40290
rect 38894 40226 38946 40238
rect 1344 40010 78624 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 78624 40010
rect 1344 39924 78624 39958
rect 77198 39730 77250 39742
rect 77198 39666 77250 39678
rect 2146 39566 2158 39618
rect 2210 39566 2222 39618
rect 3042 39566 3054 39618
rect 3106 39566 3118 39618
rect 75282 39566 75294 39618
rect 75346 39566 75358 39618
rect 3614 39506 3666 39518
rect 3614 39442 3666 39454
rect 38782 39506 38834 39518
rect 38782 39442 38834 39454
rect 39118 39506 39170 39518
rect 39118 39442 39170 39454
rect 39678 39506 39730 39518
rect 39678 39442 39730 39454
rect 40574 39506 40626 39518
rect 40574 39442 40626 39454
rect 40910 39506 40962 39518
rect 76178 39454 76190 39506
rect 76242 39454 76254 39506
rect 40910 39442 40962 39454
rect 38334 39394 38386 39406
rect 38334 39330 38386 39342
rect 40014 39394 40066 39406
rect 40014 39330 40066 39342
rect 41358 39394 41410 39406
rect 41358 39330 41410 39342
rect 74734 39394 74786 39406
rect 74734 39330 74786 39342
rect 1344 39226 78624 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 78624 39226
rect 1344 39140 78624 39174
rect 38334 38946 38386 38958
rect 2146 38894 2158 38946
rect 2210 38894 2222 38946
rect 38334 38882 38386 38894
rect 39790 38946 39842 38958
rect 77746 38894 77758 38946
rect 77810 38894 77822 38946
rect 39790 38882 39842 38894
rect 3614 38834 3666 38846
rect 3042 38782 3054 38834
rect 3106 38782 3118 38834
rect 3614 38770 3666 38782
rect 38670 38834 38722 38846
rect 40686 38834 40738 38846
rect 39554 38782 39566 38834
rect 39618 38782 39630 38834
rect 75058 38782 75070 38834
rect 75122 38782 75134 38834
rect 76850 38782 76862 38834
rect 76914 38782 76926 38834
rect 38670 38770 38722 38782
rect 40686 38770 40738 38782
rect 37886 38722 37938 38734
rect 37886 38658 37938 38670
rect 40238 38722 40290 38734
rect 40238 38658 40290 38670
rect 74622 38722 74674 38734
rect 76066 38670 76078 38722
rect 76130 38670 76142 38722
rect 74622 38658 74674 38670
rect 1344 38442 78624 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 78624 38442
rect 1344 38356 78624 38390
rect 76638 38162 76690 38174
rect 2034 38110 2046 38162
rect 2098 38110 2110 38162
rect 76638 38098 76690 38110
rect 3042 37998 3054 38050
rect 3106 37998 3118 38050
rect 37998 37938 38050 37950
rect 37998 37874 38050 37886
rect 38670 37938 38722 37950
rect 38670 37874 38722 37886
rect 39454 37938 39506 37950
rect 39454 37874 39506 37886
rect 3614 37826 3666 37838
rect 3614 37762 3666 37774
rect 37662 37826 37714 37838
rect 37662 37762 37714 37774
rect 39006 37826 39058 37838
rect 39006 37762 39058 37774
rect 1344 37658 78624 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 78624 37658
rect 1344 37572 78624 37606
rect 36990 37378 37042 37390
rect 2146 37326 2158 37378
rect 2210 37326 2222 37378
rect 36990 37314 37042 37326
rect 38334 37378 38386 37390
rect 77746 37326 77758 37378
rect 77810 37326 77822 37378
rect 38334 37314 38386 37326
rect 37998 37266 38050 37278
rect 3042 37214 3054 37266
rect 3106 37214 3118 37266
rect 37202 37214 37214 37266
rect 37266 37214 37278 37266
rect 75058 37214 75070 37266
rect 75122 37214 75134 37266
rect 76850 37214 76862 37266
rect 76914 37214 76926 37266
rect 37998 37202 38050 37214
rect 3614 37154 3666 37166
rect 3614 37090 3666 37102
rect 36542 37154 36594 37166
rect 36542 37090 36594 37102
rect 38782 37154 38834 37166
rect 38782 37090 38834 37102
rect 74622 37154 74674 37166
rect 76066 37102 76078 37154
rect 76130 37102 76142 37154
rect 74622 37090 74674 37102
rect 1344 36874 78624 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 78624 36874
rect 1344 36788 78624 36822
rect 38334 36594 38386 36606
rect 2034 36542 2046 36594
rect 2098 36542 2110 36594
rect 38334 36530 38386 36542
rect 76638 36594 76690 36606
rect 76638 36530 76690 36542
rect 3042 36430 3054 36482
rect 3106 36430 3118 36482
rect 35870 36370 35922 36382
rect 35870 36306 35922 36318
rect 36654 36370 36706 36382
rect 36654 36306 36706 36318
rect 37550 36370 37602 36382
rect 37550 36306 37602 36318
rect 38782 36370 38834 36382
rect 38782 36306 38834 36318
rect 3614 36258 3666 36270
rect 3614 36194 3666 36206
rect 35310 36258 35362 36270
rect 35310 36194 35362 36206
rect 36318 36258 36370 36270
rect 36318 36194 36370 36206
rect 37886 36258 37938 36270
rect 37886 36194 37938 36206
rect 1344 36090 78624 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 78624 36090
rect 1344 36004 78624 36038
rect 34638 35810 34690 35822
rect 2146 35758 2158 35810
rect 2210 35758 2222 35810
rect 34638 35746 34690 35758
rect 35534 35810 35586 35822
rect 35534 35746 35586 35758
rect 35870 35810 35922 35822
rect 35870 35746 35922 35758
rect 36990 35810 37042 35822
rect 77746 35758 77758 35810
rect 77810 35758 77822 35810
rect 36990 35746 37042 35758
rect 34974 35698 35026 35710
rect 37438 35698 37490 35710
rect 3042 35646 3054 35698
rect 3106 35646 3118 35698
rect 4834 35646 4846 35698
rect 4898 35646 4910 35698
rect 36754 35646 36766 35698
rect 36818 35646 36830 35698
rect 75058 35646 75070 35698
rect 75122 35646 75134 35698
rect 76850 35646 76862 35698
rect 76914 35646 76926 35698
rect 34974 35634 35026 35646
rect 37438 35634 37490 35646
rect 5406 35586 5458 35598
rect 3826 35534 3838 35586
rect 3890 35534 3902 35586
rect 5406 35522 5458 35534
rect 74622 35586 74674 35598
rect 76066 35534 76078 35586
rect 76130 35534 76142 35586
rect 74622 35522 74674 35534
rect 1344 35306 78624 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 78624 35306
rect 1344 35220 78624 35254
rect 3614 35026 3666 35038
rect 2034 34974 2046 35026
rect 2098 34974 2110 35026
rect 3614 34962 3666 34974
rect 77198 35026 77250 35038
rect 77198 34962 77250 34974
rect 33742 34914 33794 34926
rect 3042 34862 3054 34914
rect 3106 34862 3118 34914
rect 33742 34850 33794 34862
rect 34526 34914 34578 34926
rect 35186 34862 35198 34914
rect 35250 34862 35262 34914
rect 36082 34862 36094 34914
rect 36146 34862 36158 34914
rect 75282 34862 75294 34914
rect 75346 34862 75358 34914
rect 34526 34850 34578 34862
rect 34190 34802 34242 34814
rect 34190 34738 34242 34750
rect 36318 34802 36370 34814
rect 76178 34750 76190 34802
rect 76242 34750 76254 34802
rect 36318 34738 36370 34750
rect 4062 34690 4114 34702
rect 4062 34626 4114 34638
rect 35422 34690 35474 34702
rect 35422 34626 35474 34638
rect 36766 34690 36818 34702
rect 36766 34626 36818 34638
rect 74734 34690 74786 34702
rect 74734 34626 74786 34638
rect 1344 34522 78624 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 78624 34522
rect 1344 34436 78624 34470
rect 33630 34242 33682 34254
rect 2146 34190 2158 34242
rect 2210 34190 2222 34242
rect 33630 34178 33682 34190
rect 35086 34242 35138 34254
rect 77746 34190 77758 34242
rect 77810 34190 77822 34242
rect 35086 34178 35138 34190
rect 32958 34130 33010 34142
rect 3042 34078 3054 34130
rect 3106 34078 3118 34130
rect 32958 34066 33010 34078
rect 33966 34130 34018 34142
rect 34850 34078 34862 34130
rect 34914 34078 34926 34130
rect 75058 34078 75070 34130
rect 75122 34078 75134 34130
rect 76850 34078 76862 34130
rect 76914 34078 76926 34130
rect 33966 34066 34018 34078
rect 3614 34018 3666 34030
rect 3614 33954 3666 33966
rect 35646 34018 35698 34030
rect 35646 33954 35698 33966
rect 36094 34018 36146 34030
rect 36094 33954 36146 33966
rect 74622 34018 74674 34030
rect 76066 33966 76078 34018
rect 76130 33966 76142 34018
rect 74622 33954 74674 33966
rect 35970 33854 35982 33906
rect 36034 33903 36046 33906
rect 36194 33903 36206 33906
rect 36034 33857 36206 33903
rect 36034 33854 36046 33857
rect 36194 33854 36206 33857
rect 36258 33854 36270 33906
rect 1344 33738 78624 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 78624 33738
rect 1344 33652 78624 33686
rect 76638 33458 76690 33470
rect 2034 33406 2046 33458
rect 2098 33406 2110 33458
rect 76638 33394 76690 33406
rect 32510 33346 32562 33358
rect 34078 33346 34130 33358
rect 3042 33294 3054 33346
rect 3106 33294 3118 33346
rect 33170 33294 33182 33346
rect 33234 33294 33246 33346
rect 32510 33282 32562 33294
rect 34078 33282 34130 33294
rect 3614 33122 3666 33134
rect 3614 33058 3666 33070
rect 32958 33122 33010 33134
rect 32958 33058 33010 33070
rect 34414 33122 34466 33134
rect 34414 33058 34466 33070
rect 34862 33122 34914 33134
rect 34862 33058 34914 33070
rect 1344 32954 78624 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 78624 32954
rect 1344 32868 78624 32902
rect 34414 32786 34466 32798
rect 34414 32722 34466 32734
rect 32174 32674 32226 32686
rect 2146 32622 2158 32674
rect 2210 32622 2222 32674
rect 32174 32610 32226 32622
rect 33966 32674 34018 32686
rect 77746 32622 77758 32674
rect 77810 32622 77822 32674
rect 33966 32610 34018 32622
rect 32510 32562 32562 32574
rect 3042 32510 3054 32562
rect 3106 32510 3118 32562
rect 32510 32498 32562 32510
rect 33630 32562 33682 32574
rect 33630 32498 33682 32510
rect 74622 32562 74674 32574
rect 75058 32510 75070 32562
rect 75122 32510 75134 32562
rect 76850 32510 76862 32562
rect 76914 32510 76926 32562
rect 74622 32498 74674 32510
rect 3614 32450 3666 32462
rect 3614 32386 3666 32398
rect 31726 32450 31778 32462
rect 76066 32398 76078 32450
rect 76130 32398 76142 32450
rect 31726 32386 31778 32398
rect 1344 32170 78624 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 78624 32170
rect 1344 32084 78624 32118
rect 33406 31890 33458 31902
rect 2034 31838 2046 31890
rect 2098 31838 2110 31890
rect 33406 31826 33458 31838
rect 76638 31890 76690 31902
rect 76638 31826 76690 31838
rect 3042 31726 3054 31778
rect 3106 31726 3118 31778
rect 31166 31666 31218 31678
rect 31166 31602 31218 31614
rect 31950 31666 32002 31678
rect 31950 31602 32002 31614
rect 32622 31666 32674 31678
rect 32622 31602 32674 31614
rect 33854 31666 33906 31678
rect 33854 31602 33906 31614
rect 3614 31554 3666 31566
rect 3614 31490 3666 31502
rect 30718 31554 30770 31566
rect 30718 31490 30770 31502
rect 31614 31554 31666 31566
rect 31614 31490 31666 31502
rect 32958 31554 33010 31566
rect 32958 31490 33010 31502
rect 1344 31386 78624 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 78624 31386
rect 1344 31300 78624 31334
rect 30046 31106 30098 31118
rect 2146 31054 2158 31106
rect 2210 31054 2222 31106
rect 30046 31042 30098 31054
rect 30942 31106 30994 31118
rect 30942 31042 30994 31054
rect 32286 31106 32338 31118
rect 77746 31054 77758 31106
rect 77810 31054 77822 31106
rect 32286 31042 32338 31054
rect 31278 30994 31330 31006
rect 32734 30994 32786 31006
rect 3042 30942 3054 30994
rect 3106 30942 3118 30994
rect 4834 30942 4846 30994
rect 4898 30942 4910 30994
rect 30258 30942 30270 30994
rect 30322 30942 30334 30994
rect 32050 30942 32062 30994
rect 32114 30942 32126 30994
rect 75058 30942 75070 30994
rect 75122 30942 75134 30994
rect 76850 30942 76862 30994
rect 76914 30942 76926 30994
rect 31278 30930 31330 30942
rect 32734 30930 32786 30942
rect 5406 30882 5458 30894
rect 3826 30830 3838 30882
rect 3890 30830 3902 30882
rect 5406 30818 5458 30830
rect 74622 30882 74674 30894
rect 76066 30830 76078 30882
rect 76130 30830 76142 30882
rect 74622 30818 74674 30830
rect 1344 30602 78624 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 78624 30602
rect 1344 30516 78624 30550
rect 32062 30322 32114 30334
rect 32062 30258 32114 30270
rect 77198 30322 77250 30334
rect 77198 30258 77250 30270
rect 3614 30210 3666 30222
rect 2146 30158 2158 30210
rect 2210 30158 2222 30210
rect 3042 30158 3054 30210
rect 3106 30158 3118 30210
rect 75282 30158 75294 30210
rect 75346 30158 75358 30210
rect 3614 30146 3666 30158
rect 30382 30098 30434 30110
rect 30382 30034 30434 30046
rect 31278 30098 31330 30110
rect 31278 30034 31330 30046
rect 31614 30098 31666 30110
rect 76178 30046 76190 30098
rect 76242 30046 76254 30098
rect 31614 30034 31666 30046
rect 4062 29986 4114 29998
rect 4062 29922 4114 29934
rect 29934 29986 29986 29998
rect 29934 29922 29986 29934
rect 30718 29986 30770 29998
rect 30718 29922 30770 29934
rect 74734 29986 74786 29998
rect 74734 29922 74786 29934
rect 1344 29818 78624 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 78624 29818
rect 1344 29732 78624 29766
rect 29598 29650 29650 29662
rect 29598 29586 29650 29598
rect 28702 29538 28754 29550
rect 2146 29486 2158 29538
rect 2210 29486 2222 29538
rect 28702 29474 28754 29486
rect 30830 29538 30882 29550
rect 77746 29486 77758 29538
rect 77810 29486 77822 29538
rect 30830 29474 30882 29486
rect 29038 29426 29090 29438
rect 3042 29374 3054 29426
rect 3106 29374 3118 29426
rect 29038 29362 29090 29374
rect 29934 29426 29986 29438
rect 29934 29362 29986 29374
rect 30494 29426 30546 29438
rect 75058 29374 75070 29426
rect 75122 29374 75134 29426
rect 76850 29374 76862 29426
rect 76914 29374 76926 29426
rect 30494 29362 30546 29374
rect 3614 29314 3666 29326
rect 3614 29250 3666 29262
rect 28254 29314 28306 29326
rect 28254 29250 28306 29262
rect 31278 29314 31330 29326
rect 31278 29250 31330 29262
rect 74622 29314 74674 29326
rect 76066 29262 76078 29314
rect 76130 29262 76142 29314
rect 74622 29250 74674 29262
rect 1344 29034 78624 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 78624 29034
rect 1344 28948 78624 28982
rect 30258 28814 30270 28866
rect 30322 28863 30334 28866
rect 30930 28863 30942 28866
rect 30322 28817 30942 28863
rect 30322 28814 30334 28817
rect 30930 28814 30942 28817
rect 30994 28814 31006 28866
rect 76638 28754 76690 28766
rect 2034 28702 2046 28754
rect 2098 28702 2110 28754
rect 76638 28690 76690 28702
rect 3614 28642 3666 28654
rect 3042 28590 3054 28642
rect 3106 28590 3118 28642
rect 3614 28578 3666 28590
rect 27806 28642 27858 28654
rect 27806 28578 27858 28590
rect 30382 28642 30434 28654
rect 30382 28578 30434 28590
rect 30830 28642 30882 28654
rect 30830 28578 30882 28590
rect 28254 28530 28306 28542
rect 28254 28466 28306 28478
rect 28590 28530 28642 28542
rect 28590 28466 28642 28478
rect 29598 28530 29650 28542
rect 29598 28466 29650 28478
rect 29934 28418 29986 28430
rect 29934 28354 29986 28366
rect 1344 28250 78624 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 78624 28250
rect 1344 28164 78624 28198
rect 27582 27970 27634 27982
rect 2146 27918 2158 27970
rect 2210 27918 2222 27970
rect 27582 27906 27634 27918
rect 28926 27970 28978 27982
rect 77746 27918 77758 27970
rect 77810 27918 77822 27970
rect 28926 27906 28978 27918
rect 27134 27858 27186 27870
rect 3042 27806 3054 27858
rect 3106 27806 3118 27858
rect 27134 27794 27186 27806
rect 27918 27858 27970 27870
rect 27918 27794 27970 27806
rect 28590 27858 28642 27870
rect 28590 27794 28642 27806
rect 29822 27858 29874 27870
rect 75058 27806 75070 27858
rect 75122 27806 75134 27858
rect 76850 27806 76862 27858
rect 76914 27806 76926 27858
rect 29822 27794 29874 27806
rect 3614 27746 3666 27758
rect 3614 27682 3666 27694
rect 29374 27746 29426 27758
rect 29374 27682 29426 27694
rect 74622 27746 74674 27758
rect 76066 27694 76078 27746
rect 76130 27694 76142 27746
rect 74622 27682 74674 27694
rect 1344 27466 78624 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 78624 27466
rect 1344 27380 78624 27414
rect 76638 27186 76690 27198
rect 2034 27134 2046 27186
rect 2098 27134 2110 27186
rect 76638 27122 76690 27134
rect 3614 27074 3666 27086
rect 3042 27022 3054 27074
rect 3106 27022 3118 27074
rect 3614 27010 3666 27022
rect 26462 26962 26514 26974
rect 26462 26898 26514 26910
rect 27246 26962 27298 26974
rect 27246 26898 27298 26910
rect 28030 26962 28082 26974
rect 28030 26898 28082 26910
rect 28814 26962 28866 26974
rect 28814 26898 28866 26910
rect 26910 26850 26962 26862
rect 26910 26786 26962 26798
rect 28366 26850 28418 26862
rect 28366 26786 28418 26798
rect 1344 26682 78624 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 78624 26682
rect 1344 26596 78624 26630
rect 26238 26402 26290 26414
rect 2146 26350 2158 26402
rect 2210 26350 2222 26402
rect 26238 26338 26290 26350
rect 27694 26402 27746 26414
rect 77746 26350 77758 26402
rect 77810 26350 77822 26402
rect 27694 26338 27746 26350
rect 27358 26290 27410 26302
rect 2930 26238 2942 26290
rect 2994 26238 3006 26290
rect 4834 26238 4846 26290
rect 4898 26238 4910 26290
rect 26450 26238 26462 26290
rect 26514 26238 26526 26290
rect 75058 26238 75070 26290
rect 75122 26238 75134 26290
rect 76850 26238 76862 26290
rect 76914 26238 76926 26290
rect 27358 26226 27410 26238
rect 5406 26178 5458 26190
rect 3826 26126 3838 26178
rect 3890 26126 3902 26178
rect 5406 26114 5458 26126
rect 25790 26178 25842 26190
rect 25790 26114 25842 26126
rect 74622 26178 74674 26190
rect 76066 26126 76078 26178
rect 76130 26126 76142 26178
rect 74622 26114 74674 26126
rect 1344 25898 78624 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 78624 25898
rect 1344 25812 78624 25846
rect 77198 25618 77250 25630
rect 2034 25566 2046 25618
rect 2098 25566 2110 25618
rect 77198 25554 77250 25566
rect 25566 25506 25618 25518
rect 3042 25454 3054 25506
rect 3106 25454 3118 25506
rect 25566 25442 25618 25454
rect 27582 25506 27634 25518
rect 75282 25454 75294 25506
rect 75346 25454 75358 25506
rect 27582 25442 27634 25454
rect 4062 25394 4114 25406
rect 4062 25330 4114 25342
rect 24334 25394 24386 25406
rect 24334 25330 24386 25342
rect 24670 25394 24722 25406
rect 24670 25330 24722 25342
rect 25230 25394 25282 25406
rect 25230 25330 25282 25342
rect 26350 25394 26402 25406
rect 26350 25330 26402 25342
rect 27134 25394 27186 25406
rect 76178 25342 76190 25394
rect 76242 25342 76254 25394
rect 27134 25330 27186 25342
rect 3614 25282 3666 25294
rect 3614 25218 3666 25230
rect 26686 25282 26738 25294
rect 26686 25218 26738 25230
rect 74734 25282 74786 25294
rect 74734 25218 74786 25230
rect 1344 25114 78624 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 78624 25114
rect 1344 25028 78624 25062
rect 24110 24834 24162 24846
rect 2146 24782 2158 24834
rect 2210 24782 2222 24834
rect 24110 24770 24162 24782
rect 26126 24834 26178 24846
rect 77746 24782 77758 24834
rect 77810 24782 77822 24834
rect 26126 24770 26178 24782
rect 24446 24722 24498 24734
rect 3042 24670 3054 24722
rect 3106 24670 3118 24722
rect 25890 24670 25902 24722
rect 25954 24670 25966 24722
rect 75058 24670 75070 24722
rect 75122 24670 75134 24722
rect 76850 24670 76862 24722
rect 76914 24670 76926 24722
rect 24446 24658 24498 24670
rect 3614 24610 3666 24622
rect 3614 24546 3666 24558
rect 24894 24610 24946 24622
rect 24894 24546 24946 24558
rect 26574 24610 26626 24622
rect 26574 24546 26626 24558
rect 27022 24610 27074 24622
rect 27022 24546 27074 24558
rect 74622 24610 74674 24622
rect 76066 24558 76078 24610
rect 76130 24558 76142 24610
rect 74622 24546 74674 24558
rect 26338 24446 26350 24498
rect 26402 24495 26414 24498
rect 26562 24495 26574 24498
rect 26402 24449 26574 24495
rect 26402 24446 26414 24449
rect 26562 24446 26574 24449
rect 26626 24446 26638 24498
rect 1344 24330 78624 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 78624 24330
rect 1344 24244 78624 24278
rect 76638 24050 76690 24062
rect 2034 23998 2046 24050
rect 2098 23998 2110 24050
rect 76638 23986 76690 23998
rect 3042 23886 3054 23938
rect 3106 23886 3118 23938
rect 25554 23886 25566 23938
rect 25618 23886 25630 23938
rect 23998 23826 24050 23838
rect 23998 23762 24050 23774
rect 26350 23826 26402 23838
rect 26350 23762 26402 23774
rect 26686 23826 26738 23838
rect 26686 23762 26738 23774
rect 3614 23714 3666 23726
rect 3614 23650 3666 23662
rect 23102 23714 23154 23726
rect 23102 23650 23154 23662
rect 23662 23714 23714 23726
rect 23662 23650 23714 23662
rect 24670 23714 24722 23726
rect 24670 23650 24722 23662
rect 25790 23714 25842 23726
rect 25790 23650 25842 23662
rect 1344 23546 78624 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 78624 23546
rect 1344 23460 78624 23494
rect 26014 23378 26066 23390
rect 26014 23314 26066 23326
rect 22430 23266 22482 23278
rect 2146 23214 2158 23266
rect 2210 23214 2222 23266
rect 22430 23202 22482 23214
rect 23886 23266 23938 23278
rect 77746 23214 77758 23266
rect 77810 23214 77822 23266
rect 23886 23202 23938 23214
rect 22766 23154 22818 23166
rect 24782 23154 24834 23166
rect 3042 23102 3054 23154
rect 3106 23102 3118 23154
rect 23650 23102 23662 23154
rect 23714 23102 23726 23154
rect 75058 23102 75070 23154
rect 75122 23102 75134 23154
rect 76850 23102 76862 23154
rect 76914 23102 76926 23154
rect 22766 23090 22818 23102
rect 24782 23090 24834 23102
rect 3614 23042 3666 23054
rect 3614 22978 3666 22990
rect 24334 23042 24386 23054
rect 24334 22978 24386 22990
rect 25566 23042 25618 23054
rect 25566 22978 25618 22990
rect 74622 23042 74674 23054
rect 76066 22990 76078 23042
rect 76130 22990 76142 23042
rect 74622 22978 74674 22990
rect 1344 22762 78624 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 78624 22762
rect 1344 22676 78624 22710
rect 76638 22482 76690 22494
rect 2034 22430 2046 22482
rect 2098 22430 2110 22482
rect 76638 22418 76690 22430
rect 3042 22318 3054 22370
rect 3106 22318 3118 22370
rect 3614 22258 3666 22270
rect 3614 22194 3666 22206
rect 22094 22258 22146 22270
rect 22094 22194 22146 22206
rect 22430 22258 22482 22270
rect 22430 22194 22482 22206
rect 22990 22258 23042 22270
rect 22990 22194 23042 22206
rect 21646 22146 21698 22158
rect 21646 22082 21698 22094
rect 23326 22146 23378 22158
rect 23326 22082 23378 22094
rect 1344 21978 78624 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 78624 21978
rect 1344 21892 78624 21926
rect 21646 21698 21698 21710
rect 2146 21646 2158 21698
rect 2210 21646 2222 21698
rect 21646 21634 21698 21646
rect 23998 21698 24050 21710
rect 77746 21646 77758 21698
rect 77810 21646 77822 21698
rect 23998 21634 24050 21646
rect 23662 21586 23714 21598
rect 2930 21534 2942 21586
rect 2994 21534 3006 21586
rect 4834 21534 4846 21586
rect 4898 21534 4910 21586
rect 21858 21534 21870 21586
rect 21922 21534 21934 21586
rect 75058 21534 75070 21586
rect 75122 21534 75134 21586
rect 76850 21534 76862 21586
rect 76914 21534 76926 21586
rect 23662 21522 23714 21534
rect 5406 21474 5458 21486
rect 3826 21422 3838 21474
rect 3890 21422 3902 21474
rect 5406 21410 5458 21422
rect 22654 21474 22706 21486
rect 22654 21410 22706 21422
rect 23102 21474 23154 21486
rect 23102 21410 23154 21422
rect 74622 21474 74674 21486
rect 76066 21422 76078 21474
rect 76130 21422 76142 21474
rect 74622 21410 74674 21422
rect 1344 21194 78624 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 78624 21194
rect 1344 21108 78624 21142
rect 77198 20914 77250 20926
rect 2034 20862 2046 20914
rect 2098 20862 2110 20914
rect 77198 20850 77250 20862
rect 3042 20750 3054 20802
rect 3106 20750 3118 20802
rect 75282 20750 75294 20802
rect 75346 20750 75358 20802
rect 4062 20690 4114 20702
rect 4062 20626 4114 20638
rect 21646 20690 21698 20702
rect 21646 20626 21698 20638
rect 21982 20690 22034 20702
rect 21982 20626 22034 20638
rect 23214 20690 23266 20702
rect 76178 20638 76190 20690
rect 76242 20638 76254 20690
rect 23214 20626 23266 20638
rect 3614 20578 3666 20590
rect 3614 20514 3666 20526
rect 20638 20578 20690 20590
rect 20638 20514 20690 20526
rect 22430 20578 22482 20590
rect 22430 20514 22482 20526
rect 23550 20578 23602 20590
rect 23550 20514 23602 20526
rect 74734 20578 74786 20590
rect 74734 20514 74786 20526
rect 1344 20410 78624 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 78624 20410
rect 1344 20324 78624 20358
rect 19966 20242 20018 20254
rect 19966 20178 20018 20190
rect 21198 20130 21250 20142
rect 2146 20078 2158 20130
rect 2210 20078 2222 20130
rect 77746 20078 77758 20130
rect 77810 20078 77822 20130
rect 21198 20066 21250 20078
rect 19518 20018 19570 20030
rect 3042 19966 3054 20018
rect 3106 19966 3118 20018
rect 19518 19954 19570 19966
rect 20302 20018 20354 20030
rect 20302 19954 20354 19966
rect 20862 20018 20914 20030
rect 75058 19966 75070 20018
rect 75122 19966 75134 20018
rect 76850 19966 76862 20018
rect 76914 19966 76926 20018
rect 20862 19954 20914 19966
rect 3614 19906 3666 19918
rect 3614 19842 3666 19854
rect 21758 19906 21810 19918
rect 21758 19842 21810 19854
rect 22206 19906 22258 19918
rect 22206 19842 22258 19854
rect 22878 19906 22930 19918
rect 22878 19842 22930 19854
rect 74622 19906 74674 19918
rect 76066 19854 76078 19906
rect 76130 19854 76142 19906
rect 74622 19842 74674 19854
rect 1344 19626 78624 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 78624 19626
rect 1344 19540 78624 19574
rect 76638 19346 76690 19358
rect 2034 19294 2046 19346
rect 2098 19294 2110 19346
rect 76638 19282 76690 19294
rect 3042 19182 3054 19234
rect 3106 19182 3118 19234
rect 20514 19182 20526 19234
rect 20578 19182 20590 19234
rect 18958 19122 19010 19134
rect 18958 19058 19010 19070
rect 19518 19122 19570 19134
rect 19518 19058 19570 19070
rect 19854 19122 19906 19134
rect 19854 19058 19906 19070
rect 21646 19122 21698 19134
rect 21646 19058 21698 19070
rect 21982 19122 22034 19134
rect 21982 19058 22034 19070
rect 3614 19010 3666 19022
rect 3614 18946 3666 18958
rect 18174 19010 18226 19022
rect 18174 18946 18226 18958
rect 18622 19010 18674 19022
rect 18622 18946 18674 18958
rect 20750 19010 20802 19022
rect 20750 18946 20802 18958
rect 1344 18842 78624 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 78624 18842
rect 1344 18756 78624 18790
rect 21534 18674 21586 18686
rect 56242 18622 56254 18674
rect 56306 18622 56318 18674
rect 21534 18610 21586 18622
rect 18622 18562 18674 18574
rect 2146 18510 2158 18562
rect 2210 18510 2222 18562
rect 18622 18498 18674 18510
rect 21086 18562 21138 18574
rect 21086 18498 21138 18510
rect 55582 18562 55634 18574
rect 55582 18498 55634 18510
rect 18958 18450 19010 18462
rect 3042 18398 3054 18450
rect 3106 18398 3118 18450
rect 18958 18386 19010 18398
rect 20750 18450 20802 18462
rect 20750 18386 20802 18398
rect 55806 18450 55858 18462
rect 55806 18386 55858 18398
rect 56030 18450 56082 18462
rect 56030 18386 56082 18398
rect 56254 18450 56306 18462
rect 75058 18398 75070 18450
rect 75122 18398 75134 18450
rect 76850 18398 76862 18450
rect 76914 18398 76926 18450
rect 77746 18398 77758 18450
rect 77810 18398 77822 18450
rect 56254 18386 56306 18398
rect 3614 18338 3666 18350
rect 3614 18274 3666 18286
rect 18174 18338 18226 18350
rect 18174 18274 18226 18286
rect 19630 18338 19682 18350
rect 19630 18274 19682 18286
rect 20078 18338 20130 18350
rect 20078 18274 20130 18286
rect 54574 18338 54626 18350
rect 54574 18274 54626 18286
rect 55022 18338 55074 18350
rect 55022 18274 55074 18286
rect 74622 18338 74674 18350
rect 76066 18286 76078 18338
rect 76130 18286 76142 18338
rect 74622 18274 74674 18286
rect 1344 18058 78624 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 78624 18058
rect 1344 17972 78624 18006
rect 20526 17890 20578 17902
rect 20526 17826 20578 17838
rect 20750 17890 20802 17902
rect 20750 17826 20802 17838
rect 56142 17890 56194 17902
rect 56142 17826 56194 17838
rect 21982 17778 22034 17790
rect 55582 17778 55634 17790
rect 2034 17726 2046 17778
rect 2098 17726 2110 17778
rect 26114 17726 26126 17778
rect 26178 17726 26190 17778
rect 21982 17714 22034 17726
rect 55582 17714 55634 17726
rect 20302 17666 20354 17678
rect 3042 17614 3054 17666
rect 3106 17614 3118 17666
rect 20066 17614 20078 17666
rect 20130 17614 20142 17666
rect 20302 17602 20354 17614
rect 76638 17666 76690 17678
rect 76638 17602 76690 17614
rect 18062 17554 18114 17566
rect 18062 17490 18114 17502
rect 18622 17554 18674 17566
rect 18622 17490 18674 17502
rect 18958 17554 19010 17566
rect 18958 17490 19010 17502
rect 20862 17554 20914 17566
rect 20862 17490 20914 17502
rect 21534 17554 21586 17566
rect 21534 17490 21586 17502
rect 25790 17554 25842 17566
rect 25790 17490 25842 17502
rect 27022 17554 27074 17566
rect 27022 17490 27074 17502
rect 54798 17554 54850 17566
rect 54798 17490 54850 17502
rect 55470 17554 55522 17566
rect 55470 17490 55522 17502
rect 56030 17554 56082 17566
rect 56030 17490 56082 17502
rect 3614 17442 3666 17454
rect 3614 17378 3666 17390
rect 16382 17442 16434 17454
rect 16382 17378 16434 17390
rect 17166 17442 17218 17454
rect 17166 17378 17218 17390
rect 17726 17442 17778 17454
rect 17726 17378 17778 17390
rect 19406 17442 19458 17454
rect 19406 17378 19458 17390
rect 26014 17442 26066 17454
rect 26014 17378 26066 17390
rect 26574 17442 26626 17454
rect 26574 17378 26626 17390
rect 53566 17442 53618 17454
rect 53566 17378 53618 17390
rect 54014 17442 54066 17454
rect 54014 17378 54066 17390
rect 55022 17442 55074 17454
rect 55022 17378 55074 17390
rect 55246 17442 55298 17454
rect 55246 17378 55298 17390
rect 56590 17442 56642 17454
rect 56590 17378 56642 17390
rect 1344 17274 78624 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 78624 17274
rect 1344 17188 78624 17222
rect 19854 17106 19906 17118
rect 19854 17042 19906 17054
rect 20302 17106 20354 17118
rect 20302 17042 20354 17054
rect 20750 17106 20802 17118
rect 20750 17042 20802 17054
rect 22990 17106 23042 17118
rect 22990 17042 23042 17054
rect 74622 17106 74674 17118
rect 74622 17042 74674 17054
rect 15710 16994 15762 17006
rect 2146 16942 2158 16994
rect 2210 16942 2222 16994
rect 15710 16930 15762 16942
rect 16606 16994 16658 17006
rect 16606 16930 16658 16942
rect 18622 16994 18674 17006
rect 26014 16994 26066 17006
rect 25778 16942 25790 16994
rect 25842 16942 25854 16994
rect 77746 16942 77758 16994
rect 77810 16942 77822 16994
rect 18622 16930 18674 16942
rect 26014 16930 26066 16942
rect 5406 16882 5458 16894
rect 16942 16882 16994 16894
rect 3042 16830 3054 16882
rect 3106 16830 3118 16882
rect 4834 16830 4846 16882
rect 4898 16830 4910 16882
rect 15922 16830 15934 16882
rect 15986 16830 15998 16882
rect 5406 16818 5458 16830
rect 16942 16818 16994 16830
rect 18286 16882 18338 16894
rect 18286 16818 18338 16830
rect 19518 16882 19570 16894
rect 19518 16818 19570 16830
rect 21534 16882 21586 16894
rect 21534 16818 21586 16830
rect 21870 16882 21922 16894
rect 21870 16818 21922 16830
rect 22990 16882 23042 16894
rect 22990 16818 23042 16830
rect 24446 16882 24498 16894
rect 24446 16818 24498 16830
rect 24894 16882 24946 16894
rect 24894 16818 24946 16830
rect 25678 16882 25730 16894
rect 26686 16882 26738 16894
rect 26226 16830 26238 16882
rect 26290 16830 26302 16882
rect 25678 16818 25730 16830
rect 26686 16818 26738 16830
rect 54462 16882 54514 16894
rect 75058 16830 75070 16882
rect 75122 16830 75134 16882
rect 75954 16830 75966 16882
rect 76018 16830 76030 16882
rect 76850 16830 76862 16882
rect 76914 16830 76926 16882
rect 54462 16818 54514 16830
rect 17726 16770 17778 16782
rect 3826 16718 3838 16770
rect 3890 16718 3902 16770
rect 17726 16706 17778 16718
rect 22318 16770 22370 16782
rect 22318 16706 22370 16718
rect 23326 16770 23378 16782
rect 23326 16706 23378 16718
rect 23550 16770 23602 16782
rect 23550 16706 23602 16718
rect 23102 16658 23154 16670
rect 23102 16594 23154 16606
rect 1344 16490 78624 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 78624 16490
rect 1344 16404 78624 16438
rect 18510 16322 18562 16334
rect 16930 16270 16942 16322
rect 16994 16319 17006 16322
rect 17714 16319 17726 16322
rect 16994 16273 17726 16319
rect 16994 16270 17006 16273
rect 17714 16270 17726 16273
rect 17778 16270 17790 16322
rect 18510 16258 18562 16270
rect 22878 16322 22930 16334
rect 23202 16270 23214 16322
rect 23266 16270 23278 16322
rect 22878 16258 22930 16270
rect 3614 16210 3666 16222
rect 2034 16158 2046 16210
rect 2098 16158 2110 16210
rect 3614 16146 3666 16158
rect 16830 16210 16882 16222
rect 16830 16146 16882 16158
rect 18958 16210 19010 16222
rect 18958 16146 19010 16158
rect 77198 16210 77250 16222
rect 77198 16146 77250 16158
rect 18734 16098 18786 16110
rect 3042 16046 3054 16098
rect 3106 16046 3118 16098
rect 18274 16046 18286 16098
rect 18338 16046 18350 16098
rect 18734 16034 18786 16046
rect 19070 16098 19122 16110
rect 19070 16034 19122 16046
rect 22654 16098 22706 16110
rect 75282 16046 75294 16098
rect 75346 16046 75358 16098
rect 22654 16034 22706 16046
rect 15710 15986 15762 15998
rect 15710 15922 15762 15934
rect 16046 15986 16098 15998
rect 16046 15922 16098 15934
rect 19630 15986 19682 15998
rect 76178 15934 76190 15986
rect 76242 15934 76254 15986
rect 19630 15922 19682 15934
rect 4062 15874 4114 15886
rect 4062 15810 4114 15822
rect 17278 15874 17330 15886
rect 17278 15810 17330 15822
rect 17726 15874 17778 15886
rect 17726 15810 17778 15822
rect 19966 15874 20018 15886
rect 19966 15810 20018 15822
rect 23886 15874 23938 15886
rect 23886 15810 23938 15822
rect 74734 15874 74786 15886
rect 74734 15810 74786 15822
rect 1344 15706 78624 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 78624 15706
rect 1344 15620 78624 15654
rect 19294 15538 19346 15550
rect 19294 15474 19346 15486
rect 14702 15426 14754 15438
rect 2146 15374 2158 15426
rect 2210 15374 2222 15426
rect 14702 15362 14754 15374
rect 55918 15426 55970 15438
rect 77746 15374 77758 15426
rect 77810 15374 77822 15426
rect 55918 15362 55970 15374
rect 15038 15314 15090 15326
rect 3042 15262 3054 15314
rect 3106 15262 3118 15314
rect 15038 15250 15090 15262
rect 55022 15314 55074 15326
rect 55022 15250 55074 15262
rect 55582 15314 55634 15326
rect 75058 15262 75070 15314
rect 75122 15262 75134 15314
rect 76850 15262 76862 15314
rect 76914 15262 76926 15314
rect 55582 15250 55634 15262
rect 3614 15202 3666 15214
rect 3614 15138 3666 15150
rect 15486 15202 15538 15214
rect 15486 15138 15538 15150
rect 16270 15202 16322 15214
rect 16270 15138 16322 15150
rect 17054 15202 17106 15214
rect 17054 15138 17106 15150
rect 17726 15202 17778 15214
rect 17726 15138 17778 15150
rect 18174 15202 18226 15214
rect 18174 15138 18226 15150
rect 74622 15202 74674 15214
rect 76066 15150 76078 15202
rect 76130 15150 76142 15202
rect 74622 15138 74674 15150
rect 1344 14922 78624 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 78624 14922
rect 1344 14836 78624 14870
rect 54798 14754 54850 14766
rect 54798 14690 54850 14702
rect 53902 14642 53954 14654
rect 2034 14590 2046 14642
rect 2098 14590 2110 14642
rect 53902 14578 53954 14590
rect 76638 14642 76690 14654
rect 76638 14578 76690 14590
rect 55022 14530 55074 14542
rect 56590 14530 56642 14542
rect 3042 14478 3054 14530
rect 3106 14478 3118 14530
rect 55234 14478 55246 14530
rect 55298 14478 55310 14530
rect 55906 14478 55918 14530
rect 55970 14478 55982 14530
rect 55022 14466 55074 14478
rect 56590 14466 56642 14478
rect 14366 14418 14418 14430
rect 14366 14354 14418 14366
rect 14814 14418 14866 14430
rect 14814 14354 14866 14366
rect 53454 14418 53506 14430
rect 53454 14354 53506 14366
rect 56142 14418 56194 14430
rect 56142 14354 56194 14366
rect 3614 14306 3666 14318
rect 3614 14242 3666 14254
rect 14030 14306 14082 14318
rect 14030 14242 14082 14254
rect 55134 14306 55186 14318
rect 55134 14242 55186 14254
rect 1344 14138 78624 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 78624 14138
rect 1344 14052 78624 14086
rect 12462 13858 12514 13870
rect 2146 13806 2158 13858
rect 2210 13806 2222 13858
rect 12462 13794 12514 13806
rect 13358 13858 13410 13870
rect 13358 13794 13410 13806
rect 55582 13858 55634 13870
rect 55582 13794 55634 13806
rect 57822 13858 57874 13870
rect 77746 13806 77758 13858
rect 77810 13806 77822 13858
rect 57822 13794 57874 13806
rect 12014 13746 12066 13758
rect 3042 13694 3054 13746
rect 3106 13694 3118 13746
rect 12014 13682 12066 13694
rect 12798 13746 12850 13758
rect 12798 13682 12850 13694
rect 13694 13746 13746 13758
rect 13694 13682 13746 13694
rect 55246 13746 55298 13758
rect 55246 13682 55298 13694
rect 56702 13746 56754 13758
rect 56702 13682 56754 13694
rect 57486 13746 57538 13758
rect 57486 13682 57538 13694
rect 74622 13746 74674 13758
rect 75058 13694 75070 13746
rect 75122 13694 75134 13746
rect 76850 13694 76862 13746
rect 76914 13694 76926 13746
rect 74622 13682 74674 13694
rect 3614 13634 3666 13646
rect 3614 13570 3666 13582
rect 14142 13634 14194 13646
rect 14142 13570 14194 13582
rect 54350 13634 54402 13646
rect 76066 13582 76078 13634
rect 76130 13582 76142 13634
rect 54350 13570 54402 13582
rect 1344 13354 78624 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 78624 13354
rect 1344 13268 78624 13302
rect 54910 13074 54962 13086
rect 2034 13022 2046 13074
rect 2098 13022 2110 13074
rect 54910 13010 54962 13022
rect 76638 13074 76690 13086
rect 76638 13010 76690 13022
rect 3042 12910 3054 12962
rect 3106 12910 3118 12962
rect 3614 12738 3666 12750
rect 3614 12674 3666 12686
rect 12014 12738 12066 12750
rect 12014 12674 12066 12686
rect 13022 12738 13074 12750
rect 13022 12674 13074 12686
rect 1344 12570 78624 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 78624 12570
rect 1344 12484 78624 12518
rect 11342 12290 11394 12302
rect 2146 12238 2158 12290
rect 2210 12238 2222 12290
rect 11342 12226 11394 12238
rect 12238 12290 12290 12302
rect 12238 12226 12290 12238
rect 13582 12290 13634 12302
rect 77746 12238 77758 12290
rect 77810 12238 77822 12290
rect 13582 12226 13634 12238
rect 11678 12178 11730 12190
rect 3042 12126 3054 12178
rect 3106 12126 3118 12178
rect 4834 12126 4846 12178
rect 4898 12126 4910 12178
rect 11678 12114 11730 12126
rect 12574 12178 12626 12190
rect 12574 12114 12626 12126
rect 13246 12178 13298 12190
rect 13246 12114 13298 12126
rect 14030 12178 14082 12190
rect 75058 12126 75070 12178
rect 75122 12126 75134 12178
rect 76850 12126 76862 12178
rect 76914 12126 76926 12178
rect 14030 12114 14082 12126
rect 74622 12066 74674 12078
rect 3826 12014 3838 12066
rect 3890 12014 3902 12066
rect 76066 12014 76078 12066
rect 76130 12014 76142 12066
rect 74622 12002 74674 12014
rect 1344 11786 78624 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 78624 11786
rect 1344 11700 78624 11734
rect 3614 11506 3666 11518
rect 2034 11454 2046 11506
rect 2098 11454 2110 11506
rect 3614 11442 3666 11454
rect 4062 11506 4114 11518
rect 4062 11442 4114 11454
rect 77198 11506 77250 11518
rect 77198 11442 77250 11454
rect 3042 11342 3054 11394
rect 3106 11342 3118 11394
rect 75282 11342 75294 11394
rect 75346 11342 75358 11394
rect 10782 11282 10834 11294
rect 10782 11218 10834 11230
rect 11118 11282 11170 11294
rect 11118 11218 11170 11230
rect 11678 11282 11730 11294
rect 11678 11218 11730 11230
rect 12574 11282 12626 11294
rect 12574 11218 12626 11230
rect 12910 11282 12962 11294
rect 76178 11230 76190 11282
rect 76242 11230 76254 11282
rect 12910 11218 12962 11230
rect 12014 11170 12066 11182
rect 12014 11106 12066 11118
rect 74734 11170 74786 11182
rect 74734 11106 74786 11118
rect 1344 11002 78624 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 78624 11002
rect 1344 10916 78624 10950
rect 10110 10722 10162 10734
rect 2146 10670 2158 10722
rect 2210 10670 2222 10722
rect 10110 10658 10162 10670
rect 11454 10722 11506 10734
rect 77746 10670 77758 10722
rect 77810 10670 77822 10722
rect 11454 10658 11506 10670
rect 10446 10610 10498 10622
rect 3042 10558 3054 10610
rect 3106 10558 3118 10610
rect 10446 10546 10498 10558
rect 11118 10610 11170 10622
rect 75058 10558 75070 10610
rect 75122 10558 75134 10610
rect 76850 10558 76862 10610
rect 76914 10558 76926 10610
rect 11118 10546 11170 10558
rect 12238 10498 12290 10510
rect 12238 10434 12290 10446
rect 74622 10498 74674 10510
rect 76066 10446 76078 10498
rect 76130 10446 76142 10498
rect 74622 10434 74674 10446
rect 1344 10218 78624 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 78624 10218
rect 1344 10132 78624 10166
rect 76638 9938 76690 9950
rect 2034 9886 2046 9938
rect 2098 9886 2110 9938
rect 76638 9874 76690 9886
rect 3042 9774 3054 9826
rect 3106 9774 3118 9826
rect 9650 9774 9662 9826
rect 9714 9774 9726 9826
rect 9438 9714 9490 9726
rect 9438 9650 9490 9662
rect 10558 9714 10610 9726
rect 10558 9650 10610 9662
rect 10894 9602 10946 9614
rect 10894 9538 10946 9550
rect 1344 9434 78624 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 78624 9434
rect 1344 9348 78624 9382
rect 8654 9154 8706 9166
rect 2146 9102 2158 9154
rect 2210 9102 2222 9154
rect 8654 9090 8706 9102
rect 10222 9154 10274 9166
rect 77746 9102 77758 9154
rect 77810 9102 77822 9154
rect 10222 9090 10274 9102
rect 8990 9042 9042 9054
rect 3042 8990 3054 9042
rect 3106 8990 3118 9042
rect 8990 8978 9042 8990
rect 9886 9042 9938 9054
rect 9886 8978 9938 8990
rect 74622 9042 74674 9054
rect 75058 8990 75070 9042
rect 75122 8990 75134 9042
rect 76850 8990 76862 9042
rect 76914 8990 76926 9042
rect 74622 8978 74674 8990
rect 76066 8878 76078 8930
rect 76130 8878 76142 8930
rect 1344 8650 78624 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 78624 8650
rect 1344 8564 78624 8598
rect 76638 8370 76690 8382
rect 2034 8318 2046 8370
rect 2098 8318 2110 8370
rect 76638 8306 76690 8318
rect 3042 8206 3054 8258
rect 3106 8206 3118 8258
rect 7982 8146 8034 8158
rect 7982 8082 8034 8094
rect 8318 8146 8370 8158
rect 8318 8082 8370 8094
rect 9102 8146 9154 8158
rect 9102 8082 9154 8094
rect 9438 8034 9490 8046
rect 9438 7970 9490 7982
rect 1344 7866 78624 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 78624 7866
rect 1344 7780 78624 7814
rect 6526 7586 6578 7598
rect 2146 7534 2158 7586
rect 2210 7534 2222 7586
rect 6526 7522 6578 7534
rect 7422 7586 7474 7598
rect 7422 7522 7474 7534
rect 8766 7586 8818 7598
rect 77746 7534 77758 7586
rect 77810 7534 77822 7586
rect 8766 7522 8818 7534
rect 6862 7474 6914 7486
rect 8430 7474 8482 7486
rect 3042 7422 3054 7474
rect 3106 7422 3118 7474
rect 4834 7422 4846 7474
rect 4898 7422 4910 7474
rect 7634 7422 7646 7474
rect 7698 7422 7710 7474
rect 75058 7422 75070 7474
rect 75122 7422 75134 7474
rect 76850 7422 76862 7474
rect 76914 7422 76926 7474
rect 6862 7410 6914 7422
rect 8430 7410 8482 7422
rect 74622 7362 74674 7374
rect 3826 7310 3838 7362
rect 3890 7310 3902 7362
rect 76066 7310 76078 7362
rect 76130 7310 76142 7362
rect 74622 7298 74674 7310
rect 1344 7082 78624 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 78624 7082
rect 1344 6996 78624 7030
rect 77198 6802 77250 6814
rect 77198 6738 77250 6750
rect 7758 6690 7810 6702
rect 2146 6638 2158 6690
rect 2210 6638 2222 6690
rect 3042 6638 3054 6690
rect 3106 6638 3118 6690
rect 75282 6638 75294 6690
rect 75346 6638 75358 6690
rect 7758 6626 7810 6638
rect 5966 6578 6018 6590
rect 5966 6514 6018 6526
rect 6302 6578 6354 6590
rect 6302 6514 6354 6526
rect 6862 6578 6914 6590
rect 6862 6514 6914 6526
rect 8094 6578 8146 6590
rect 76178 6526 76190 6578
rect 76242 6526 76254 6578
rect 8094 6514 8146 6526
rect 7198 6466 7250 6478
rect 7198 6402 7250 6414
rect 74734 6466 74786 6478
rect 74734 6402 74786 6414
rect 1344 6298 78624 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 78624 6298
rect 1344 6212 78624 6246
rect 54238 6130 54290 6142
rect 54238 6066 54290 6078
rect 55022 6130 55074 6142
rect 55022 6066 55074 6078
rect 57374 6130 57426 6142
rect 57374 6066 57426 6078
rect 58158 6130 58210 6142
rect 58158 6066 58210 6078
rect 58718 6130 58770 6142
rect 58718 6066 58770 6078
rect 59166 6130 59218 6142
rect 59166 6066 59218 6078
rect 60286 6130 60338 6142
rect 60286 6066 60338 6078
rect 60734 6130 60786 6142
rect 60734 6066 60786 6078
rect 61182 6130 61234 6142
rect 61182 6066 61234 6078
rect 61630 6130 61682 6142
rect 61630 6066 61682 6078
rect 62078 6130 62130 6142
rect 62078 6066 62130 6078
rect 64206 6130 64258 6142
rect 64206 6066 64258 6078
rect 65326 6130 65378 6142
rect 65326 6066 65378 6078
rect 65774 6130 65826 6142
rect 65774 6066 65826 6078
rect 66222 6130 66274 6142
rect 66222 6066 66274 6078
rect 66782 6130 66834 6142
rect 66782 6066 66834 6078
rect 67678 6130 67730 6142
rect 67678 6066 67730 6078
rect 69022 6130 69074 6142
rect 69022 6066 69074 6078
rect 69470 6130 69522 6142
rect 69470 6066 69522 6078
rect 5294 6018 5346 6030
rect 2146 5966 2158 6018
rect 2210 5966 2222 6018
rect 5294 5954 5346 5966
rect 6750 6018 6802 6030
rect 77746 5966 77758 6018
rect 77810 5966 77822 6018
rect 6750 5954 6802 5966
rect 5630 5906 5682 5918
rect 3042 5854 3054 5906
rect 3106 5854 3118 5906
rect 5630 5842 5682 5854
rect 6414 5906 6466 5918
rect 75058 5854 75070 5906
rect 75122 5854 75134 5906
rect 76850 5854 76862 5906
rect 76914 5854 76926 5906
rect 6414 5842 6466 5854
rect 56366 5794 56418 5806
rect 56366 5730 56418 5742
rect 67230 5794 67282 5806
rect 67230 5730 67282 5742
rect 68126 5794 68178 5806
rect 68126 5730 68178 5742
rect 74622 5794 74674 5806
rect 76066 5742 76078 5794
rect 76130 5742 76142 5794
rect 74622 5730 74674 5742
rect 66210 5630 66222 5682
rect 66274 5679 66286 5682
rect 66546 5679 66558 5682
rect 66274 5633 66558 5679
rect 66274 5630 66286 5633
rect 66546 5630 66558 5633
rect 66610 5630 66622 5682
rect 1344 5514 78624 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 78624 5514
rect 1344 5428 78624 5462
rect 49310 5234 49362 5246
rect 2034 5182 2046 5234
rect 2098 5182 2110 5234
rect 49310 5170 49362 5182
rect 49982 5234 50034 5246
rect 49982 5170 50034 5182
rect 50318 5234 50370 5246
rect 50318 5170 50370 5182
rect 51102 5234 51154 5246
rect 51102 5170 51154 5182
rect 51774 5234 51826 5246
rect 51774 5170 51826 5182
rect 52334 5234 52386 5246
rect 52334 5170 52386 5182
rect 52782 5234 52834 5246
rect 74398 5234 74450 5246
rect 54114 5182 54126 5234
rect 54178 5182 54190 5234
rect 55906 5182 55918 5234
rect 55970 5182 55982 5234
rect 57474 5182 57486 5234
rect 57538 5182 57550 5234
rect 59490 5182 59502 5234
rect 59554 5182 59566 5234
rect 62066 5182 62078 5234
rect 62130 5182 62142 5234
rect 63522 5182 63534 5234
rect 63586 5182 63598 5234
rect 65538 5182 65550 5234
rect 65602 5182 65614 5234
rect 68002 5182 68014 5234
rect 68066 5182 68078 5234
rect 70018 5182 70030 5234
rect 70082 5182 70094 5234
rect 52782 5170 52834 5182
rect 74398 5170 74450 5182
rect 76638 5234 76690 5246
rect 76638 5170 76690 5182
rect 3042 5070 3054 5122
rect 3106 5070 3118 5122
rect 53442 5070 53454 5122
rect 53506 5070 53518 5122
rect 55234 5070 55246 5122
rect 55298 5070 55310 5122
rect 58482 5070 58494 5122
rect 58546 5070 58558 5122
rect 60274 5070 60286 5122
rect 60338 5070 60350 5122
rect 61394 5070 61406 5122
rect 61458 5070 61470 5122
rect 64306 5070 64318 5122
rect 64370 5070 64382 5122
rect 66322 5070 66334 5122
rect 66386 5070 66398 5122
rect 67330 5070 67342 5122
rect 67394 5070 67406 5122
rect 69346 5070 69358 5122
rect 69410 5070 69422 5122
rect 4622 5010 4674 5022
rect 4622 4946 4674 4958
rect 4958 5010 5010 5022
rect 4958 4946 5010 4958
rect 5742 5010 5794 5022
rect 5742 4946 5794 4958
rect 72046 5010 72098 5022
rect 72046 4946 72098 4958
rect 72382 5010 72434 5022
rect 72382 4946 72434 4958
rect 6078 4898 6130 4910
rect 6078 4834 6130 4846
rect 10334 4898 10386 4910
rect 10334 4834 10386 4846
rect 12126 4898 12178 4910
rect 12126 4834 12178 4846
rect 14254 4898 14306 4910
rect 14254 4834 14306 4846
rect 16046 4898 16098 4910
rect 16046 4834 16098 4846
rect 18174 4898 18226 4910
rect 18174 4834 18226 4846
rect 20862 4898 20914 4910
rect 20862 4834 20914 4846
rect 24782 4898 24834 4910
rect 24782 4834 24834 4846
rect 26014 4898 26066 4910
rect 26014 4834 26066 4846
rect 29934 4898 29986 4910
rect 29934 4834 29986 4846
rect 30830 4898 30882 4910
rect 30830 4834 30882 4846
rect 32734 4898 32786 4910
rect 32734 4834 32786 4846
rect 35646 4898 35698 4910
rect 35646 4834 35698 4846
rect 37774 4898 37826 4910
rect 37774 4834 37826 4846
rect 47630 4898 47682 4910
rect 47630 4834 47682 4846
rect 71038 4898 71090 4910
rect 71038 4834 71090 4846
rect 71598 4898 71650 4910
rect 71598 4834 71650 4846
rect 72830 4898 72882 4910
rect 72830 4834 72882 4846
rect 73390 4898 73442 4910
rect 73390 4834 73442 4846
rect 74062 4898 74114 4910
rect 74062 4834 74114 4846
rect 74958 4898 75010 4910
rect 74958 4834 75010 4846
rect 1344 4730 78624 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 78624 4730
rect 1344 4644 78624 4678
rect 5854 4562 5906 4574
rect 5854 4498 5906 4510
rect 6862 4562 6914 4574
rect 6862 4498 6914 4510
rect 9774 4562 9826 4574
rect 9774 4498 9826 4510
rect 11902 4562 11954 4574
rect 11902 4498 11954 4510
rect 13918 4562 13970 4574
rect 13918 4498 13970 4510
rect 15934 4562 15986 4574
rect 15934 4498 15986 4510
rect 18062 4562 18114 4574
rect 18062 4498 18114 4510
rect 20638 4562 20690 4574
rect 20638 4498 20690 4510
rect 21982 4562 22034 4574
rect 21982 4498 22034 4510
rect 24670 4562 24722 4574
rect 24670 4498 24722 4510
rect 26686 4562 26738 4574
rect 26686 4498 26738 4510
rect 29374 4562 29426 4574
rect 29374 4498 29426 4510
rect 30718 4562 30770 4574
rect 30718 4498 30770 4510
rect 32734 4562 32786 4574
rect 32734 4498 32786 4510
rect 35422 4562 35474 4574
rect 35422 4498 35474 4510
rect 37438 4562 37490 4574
rect 37438 4498 37490 4510
rect 39454 4562 39506 4574
rect 39454 4498 39506 4510
rect 41918 4562 41970 4574
rect 41918 4498 41970 4510
rect 44158 4562 44210 4574
rect 44158 4498 44210 4510
rect 46846 4562 46898 4574
rect 46846 4498 46898 4510
rect 48190 4562 48242 4574
rect 48190 4498 48242 4510
rect 71150 4562 71202 4574
rect 71150 4498 71202 4510
rect 71710 4562 71762 4574
rect 71710 4498 71762 4510
rect 73726 4562 73778 4574
rect 73726 4498 73778 4510
rect 74286 4562 74338 4574
rect 74286 4498 74338 4510
rect 75182 4562 75234 4574
rect 75182 4498 75234 4510
rect 47854 4450 47906 4462
rect 47854 4386 47906 4398
rect 5518 4338 5570 4350
rect 11566 4338 11618 4350
rect 7074 4286 7086 4338
rect 7138 4286 7150 4338
rect 9986 4286 9998 4338
rect 10050 4286 10062 4338
rect 5518 4274 5570 4286
rect 11566 4274 11618 4286
rect 13582 4338 13634 4350
rect 13582 4274 13634 4286
rect 15150 4338 15202 4350
rect 15150 4274 15202 4286
rect 15598 4338 15650 4350
rect 15598 4274 15650 4286
rect 17054 4338 17106 4350
rect 17054 4274 17106 4286
rect 17726 4338 17778 4350
rect 17726 4274 17778 4286
rect 19854 4338 19906 4350
rect 19854 4274 19906 4286
rect 20302 4338 20354 4350
rect 20302 4274 20354 4286
rect 21198 4338 21250 4350
rect 21198 4274 21250 4286
rect 21646 4338 21698 4350
rect 21646 4274 21698 4286
rect 23886 4338 23938 4350
rect 23886 4274 23938 4286
rect 24334 4338 24386 4350
rect 24334 4274 24386 4286
rect 25902 4338 25954 4350
rect 25902 4274 25954 4286
rect 26350 4338 26402 4350
rect 26350 4274 26402 4286
rect 29038 4338 29090 4350
rect 29038 4274 29090 4286
rect 30382 4338 30434 4350
rect 30382 4274 30434 4286
rect 32398 4338 32450 4350
rect 32398 4274 32450 4286
rect 35086 4338 35138 4350
rect 35086 4274 35138 4286
rect 37102 4338 37154 4350
rect 37102 4274 37154 4286
rect 38670 4338 38722 4350
rect 38670 4274 38722 4286
rect 39118 4338 39170 4350
rect 39118 4274 39170 4286
rect 41582 4338 41634 4350
rect 41582 4274 41634 4286
rect 43822 4338 43874 4350
rect 43822 4274 43874 4286
rect 46510 4338 46562 4350
rect 56590 4338 56642 4350
rect 64542 4338 64594 4350
rect 70814 4338 70866 4350
rect 49522 4286 49534 4338
rect 49586 4286 49598 4338
rect 51314 4286 51326 4338
rect 51378 4286 51390 4338
rect 53106 4286 53118 4338
rect 53170 4286 53182 4338
rect 55906 4286 55918 4338
rect 55970 4286 55982 4338
rect 57586 4286 57598 4338
rect 57650 4286 57662 4338
rect 59266 4286 59278 4338
rect 59330 4286 59342 4338
rect 61058 4286 61070 4338
rect 61122 4286 61134 4338
rect 63858 4286 63870 4338
rect 63922 4286 63934 4338
rect 65650 4286 65662 4338
rect 65714 4286 65726 4338
rect 67442 4286 67454 4338
rect 67506 4286 67518 4338
rect 69122 4286 69134 4338
rect 69186 4286 69198 4338
rect 46510 4274 46562 4286
rect 56590 4274 56642 4286
rect 64542 4274 64594 4286
rect 70814 4274 70866 4286
rect 72046 4338 72098 4350
rect 72046 4274 72098 4286
rect 72494 4338 72546 4350
rect 72494 4274 72546 4286
rect 73390 4338 73442 4350
rect 74498 4286 74510 4338
rect 74562 4286 74574 4338
rect 75394 4286 75406 4338
rect 75458 4286 75470 4338
rect 73390 4274 73442 4286
rect 5070 4226 5122 4238
rect 5070 4162 5122 4174
rect 6414 4226 6466 4238
rect 6414 4162 6466 4174
rect 7646 4226 7698 4238
rect 7646 4162 7698 4174
rect 8094 4226 8146 4238
rect 8094 4162 8146 4174
rect 8654 4226 8706 4238
rect 8654 4162 8706 4174
rect 8990 4226 9042 4238
rect 8990 4162 9042 4174
rect 10670 4226 10722 4238
rect 10670 4162 10722 4174
rect 11118 4226 11170 4238
rect 11118 4162 11170 4174
rect 12686 4226 12738 4238
rect 12686 4162 12738 4174
rect 13134 4226 13186 4238
rect 13134 4162 13186 4174
rect 14702 4226 14754 4238
rect 14702 4162 14754 4174
rect 16606 4226 16658 4238
rect 16606 4162 16658 4174
rect 18846 4226 18898 4238
rect 18846 4162 18898 4174
rect 19406 4226 19458 4238
rect 19406 4162 19458 4174
rect 22430 4226 22482 4238
rect 22430 4162 22482 4174
rect 22878 4226 22930 4238
rect 22878 4162 22930 4174
rect 23438 4226 23490 4238
rect 23438 4162 23490 4174
rect 27134 4226 27186 4238
rect 27134 4162 27186 4174
rect 27582 4226 27634 4238
rect 27582 4162 27634 4174
rect 28142 4226 28194 4238
rect 28142 4162 28194 4174
rect 28590 4226 28642 4238
rect 28590 4162 28642 4174
rect 29934 4226 29986 4238
rect 29934 4162 29986 4174
rect 31502 4226 31554 4238
rect 31502 4162 31554 4174
rect 31950 4226 32002 4238
rect 31950 4162 32002 4174
rect 33630 4226 33682 4238
rect 33630 4162 33682 4174
rect 34190 4226 34242 4238
rect 34190 4162 34242 4174
rect 34638 4226 34690 4238
rect 34638 4162 34690 4174
rect 36206 4226 36258 4238
rect 36206 4162 36258 4174
rect 36654 4226 36706 4238
rect 36654 4162 36706 4174
rect 38222 4226 38274 4238
rect 38222 4162 38274 4174
rect 39902 4226 39954 4238
rect 39902 4162 39954 4174
rect 40350 4226 40402 4238
rect 40350 4162 40402 4174
rect 40910 4226 40962 4238
rect 40910 4162 40962 4174
rect 42478 4226 42530 4238
rect 42478 4162 42530 4174
rect 42926 4226 42978 4238
rect 42926 4162 42978 4174
rect 43374 4226 43426 4238
rect 43374 4162 43426 4174
rect 44718 4226 44770 4238
rect 44718 4162 44770 4174
rect 45614 4226 45666 4238
rect 45614 4162 45666 4174
rect 46062 4226 46114 4238
rect 46062 4162 46114 4174
rect 47294 4226 47346 4238
rect 47294 4162 47346 4174
rect 48638 4226 48690 4238
rect 50194 4174 50206 4226
rect 50258 4174 50270 4226
rect 52098 4174 52110 4226
rect 52162 4174 52174 4226
rect 53778 4174 53790 4226
rect 53842 4174 53854 4226
rect 55122 4174 55134 4226
rect 55186 4174 55198 4226
rect 58146 4174 58158 4226
rect 58210 4174 58222 4226
rect 59938 4174 59950 4226
rect 60002 4174 60014 4226
rect 61842 4174 61854 4226
rect 61906 4174 61918 4226
rect 63074 4174 63086 4226
rect 63138 4174 63150 4226
rect 66098 4174 66110 4226
rect 66162 4174 66174 4226
rect 67890 4174 67902 4226
rect 67954 4174 67966 4226
rect 69682 4174 69694 4226
rect 69746 4174 69758 4226
rect 48638 4162 48690 4174
rect 1344 3946 78624 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 78624 3946
rect 1344 3860 78624 3894
rect 73166 3666 73218 3678
rect 53442 3614 53454 3666
rect 53506 3614 53518 3666
rect 55234 3614 55246 3666
rect 55298 3614 55310 3666
rect 57362 3614 57374 3666
rect 57426 3614 57438 3666
rect 61282 3614 61294 3666
rect 61346 3614 61358 3666
rect 65202 3614 65214 3666
rect 65266 3614 65278 3666
rect 66994 3614 67006 3666
rect 67058 3614 67070 3666
rect 73166 3602 73218 3614
rect 17950 3554 18002 3566
rect 19406 3554 19458 3566
rect 5954 3502 5966 3554
rect 6018 3502 6030 3554
rect 12562 3502 12574 3554
rect 12626 3502 12638 3554
rect 14690 3502 14702 3554
rect 14754 3502 14766 3554
rect 15586 3502 15598 3554
rect 15650 3502 15662 3554
rect 16594 3502 16606 3554
rect 16658 3502 16670 3554
rect 18610 3502 18622 3554
rect 18674 3502 18686 3554
rect 17950 3490 18002 3502
rect 19406 3490 19458 3502
rect 20638 3554 20690 3566
rect 22766 3554 22818 3566
rect 24558 3554 24610 3566
rect 21634 3502 21646 3554
rect 21698 3502 21710 3554
rect 23426 3502 23438 3554
rect 23490 3502 23502 3554
rect 20638 3490 20690 3502
rect 22766 3490 22818 3502
rect 24558 3490 24610 3502
rect 25790 3554 25842 3566
rect 25790 3490 25842 3502
rect 26686 3554 26738 3566
rect 39342 3554 39394 3566
rect 27458 3502 27470 3554
rect 27522 3502 27534 3554
rect 29586 3502 29598 3554
rect 29650 3502 29662 3554
rect 36194 3502 36206 3554
rect 36258 3502 36270 3554
rect 38210 3502 38222 3554
rect 38274 3502 38286 3554
rect 26686 3490 26738 3502
rect 39342 3490 39394 3502
rect 40238 3554 40290 3566
rect 40238 3490 40290 3502
rect 42702 3554 42754 3566
rect 42702 3490 42754 3502
rect 43598 3554 43650 3566
rect 43598 3490 43650 3502
rect 44942 3554 44994 3566
rect 44942 3490 44994 3502
rect 45838 3554 45890 3566
rect 45838 3490 45890 3502
rect 47070 3554 47122 3566
rect 47070 3490 47122 3502
rect 47966 3554 48018 3566
rect 50082 3502 50094 3554
rect 50146 3502 50158 3554
rect 50866 3502 50878 3554
rect 50930 3502 50942 3554
rect 52770 3502 52782 3554
rect 52834 3502 52846 3554
rect 54674 3502 54686 3554
rect 54738 3502 54750 3554
rect 56690 3502 56702 3554
rect 56754 3502 56766 3554
rect 58482 3502 58494 3554
rect 58546 3502 58558 3554
rect 60610 3502 60622 3554
rect 60674 3502 60686 3554
rect 62402 3502 62414 3554
rect 62466 3502 62478 3554
rect 64530 3502 64542 3554
rect 64594 3502 64606 3554
rect 66546 3502 66558 3554
rect 66610 3502 66622 3554
rect 68450 3502 68462 3554
rect 68514 3502 68526 3554
rect 70578 3502 70590 3554
rect 70642 3502 70654 3554
rect 71250 3502 71262 3554
rect 71314 3502 71326 3554
rect 74274 3502 74286 3554
rect 74338 3502 74350 3554
rect 47966 3490 48018 3502
rect 5070 3442 5122 3454
rect 5070 3378 5122 3390
rect 6190 3442 6242 3454
rect 6190 3378 6242 3390
rect 6750 3442 6802 3454
rect 6750 3378 6802 3390
rect 7086 3442 7138 3454
rect 7086 3378 7138 3390
rect 7646 3442 7698 3454
rect 7646 3378 7698 3390
rect 7982 3442 8034 3454
rect 7982 3378 8034 3390
rect 8542 3442 8594 3454
rect 8542 3378 8594 3390
rect 10110 3442 10162 3454
rect 10110 3378 10162 3390
rect 10670 3442 10722 3454
rect 10670 3378 10722 3390
rect 11902 3442 11954 3454
rect 11902 3378 11954 3390
rect 14030 3442 14082 3454
rect 14030 3378 14082 3390
rect 28142 3442 28194 3454
rect 28142 3378 28194 3390
rect 30606 3442 30658 3454
rect 30606 3378 30658 3390
rect 31502 3442 31554 3454
rect 31502 3378 31554 3390
rect 32398 3442 32450 3454
rect 32398 3378 32450 3390
rect 33630 3442 33682 3454
rect 33630 3378 33682 3390
rect 34190 3442 34242 3454
rect 34190 3378 34242 3390
rect 35422 3442 35474 3454
rect 35422 3378 35474 3390
rect 37550 3442 37602 3454
rect 37550 3378 37602 3390
rect 41358 3442 41410 3454
rect 41358 3378 41410 3390
rect 41806 3442 41858 3454
rect 72718 3442 72770 3454
rect 49186 3390 49198 3442
rect 49250 3390 49262 3442
rect 51538 3390 51550 3442
rect 51602 3390 51614 3442
rect 59378 3390 59390 3442
rect 59442 3390 59454 3442
rect 63298 3390 63310 3442
rect 63362 3390 63374 3442
rect 69346 3390 69358 3442
rect 69410 3390 69422 3442
rect 74946 3390 74958 3442
rect 75010 3390 75022 3442
rect 41806 3378 41858 3390
rect 72718 3378 72770 3390
rect 8878 3330 8930 3342
rect 8878 3266 8930 3278
rect 9774 3330 9826 3342
rect 9774 3266 9826 3278
rect 11006 3330 11058 3342
rect 11006 3266 11058 3278
rect 11566 3330 11618 3342
rect 11566 3266 11618 3278
rect 12798 3330 12850 3342
rect 12798 3266 12850 3278
rect 13694 3330 13746 3342
rect 13694 3266 13746 3278
rect 14926 3330 14978 3342
rect 14926 3266 14978 3278
rect 15822 3330 15874 3342
rect 15822 3266 15874 3278
rect 16382 3330 16434 3342
rect 16382 3266 16434 3278
rect 17614 3330 17666 3342
rect 17614 3266 17666 3278
rect 18846 3330 18898 3342
rect 18846 3266 18898 3278
rect 19742 3330 19794 3342
rect 19742 3266 19794 3278
rect 20302 3330 20354 3342
rect 20302 3266 20354 3278
rect 21870 3330 21922 3342
rect 21870 3266 21922 3278
rect 22430 3330 22482 3342
rect 22430 3266 22482 3278
rect 23662 3330 23714 3342
rect 23662 3266 23714 3278
rect 24222 3330 24274 3342
rect 24222 3266 24274 3278
rect 25454 3330 25506 3342
rect 25454 3266 25506 3278
rect 26350 3330 26402 3342
rect 26350 3266 26402 3278
rect 27246 3330 27298 3342
rect 27246 3266 27298 3278
rect 28478 3330 28530 3342
rect 28478 3266 28530 3278
rect 29374 3330 29426 3342
rect 29374 3266 29426 3278
rect 30270 3330 30322 3342
rect 30270 3266 30322 3278
rect 31166 3330 31218 3342
rect 31166 3266 31218 3278
rect 32062 3330 32114 3342
rect 32062 3266 32114 3278
rect 33294 3330 33346 3342
rect 33294 3266 33346 3278
rect 34526 3330 34578 3342
rect 34526 3266 34578 3278
rect 35086 3330 35138 3342
rect 35086 3266 35138 3278
rect 35982 3330 36034 3342
rect 35982 3266 36034 3278
rect 37214 3330 37266 3342
rect 37214 3266 37266 3278
rect 38446 3330 38498 3342
rect 38446 3266 38498 3278
rect 39006 3330 39058 3342
rect 39006 3266 39058 3278
rect 39902 3330 39954 3342
rect 39902 3266 39954 3278
rect 42142 3330 42194 3342
rect 42142 3266 42194 3278
rect 43038 3330 43090 3342
rect 43038 3266 43090 3278
rect 43934 3330 43986 3342
rect 43934 3266 43986 3278
rect 45278 3330 45330 3342
rect 45278 3266 45330 3278
rect 46174 3330 46226 3342
rect 46174 3266 46226 3278
rect 46734 3330 46786 3342
rect 46734 3266 46786 3278
rect 47630 3330 47682 3342
rect 47630 3266 47682 3278
rect 72382 3330 72434 3342
rect 72382 3266 72434 3278
rect 1344 3162 78624 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 78624 3162
rect 1344 3076 78624 3110
<< via1 >>
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 3054 74846 3106 74898
rect 75070 74846 75122 74898
rect 76862 74846 76914 74898
rect 2046 74734 2098 74786
rect 3614 74734 3666 74786
rect 4062 74734 4114 74786
rect 76078 74734 76130 74786
rect 77870 74734 77922 74786
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 3054 74062 3106 74114
rect 2158 73950 2210 74002
rect 3614 73950 3666 74002
rect 4398 73950 4450 74002
rect 77310 73950 77362 74002
rect 78094 73950 78146 74002
rect 3950 73838 4002 73890
rect 73390 73838 73442 73890
rect 77758 73838 77810 73890
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 73726 73502 73778 73554
rect 69358 73390 69410 73442
rect 73838 73390 73890 73442
rect 3054 73278 3106 73330
rect 70030 73278 70082 73330
rect 75070 73278 75122 73330
rect 76862 73278 76914 73330
rect 2046 73166 2098 73218
rect 3614 73166 3666 73218
rect 69246 73166 69298 73218
rect 72494 73166 72546 73218
rect 76078 73166 76130 73218
rect 77870 73166 77922 73218
rect 69134 73054 69186 73106
rect 73614 73054 73666 73106
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 74062 72606 74114 72658
rect 74174 72606 74226 72658
rect 74622 72606 74674 72658
rect 3054 72494 3106 72546
rect 72158 72494 72210 72546
rect 73054 72494 73106 72546
rect 75070 72494 75122 72546
rect 2158 72382 2210 72434
rect 69358 72382 69410 72434
rect 69470 72382 69522 72434
rect 71822 72382 71874 72434
rect 73278 72382 73330 72434
rect 3502 72270 3554 72322
rect 68686 72270 68738 72322
rect 69582 72270 69634 72322
rect 73950 72270 74002 72322
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 72494 71934 72546 71986
rect 73390 71934 73442 71986
rect 74062 71934 74114 71986
rect 71150 71822 71202 71874
rect 3054 71710 3106 71762
rect 70702 71710 70754 71762
rect 71486 71710 71538 71762
rect 72270 71710 72322 71762
rect 75070 71710 75122 71762
rect 76862 71710 76914 71762
rect 2046 71598 2098 71650
rect 3614 71598 3666 71650
rect 73502 71598 73554 71650
rect 74174 71598 74226 71650
rect 76078 71598 76130 71650
rect 77870 71598 77922 71650
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 3054 70926 3106 70978
rect 71710 70926 71762 70978
rect 2158 70814 2210 70866
rect 70590 70814 70642 70866
rect 70926 70814 70978 70866
rect 71934 70814 71986 70866
rect 3502 70702 3554 70754
rect 70142 70702 70194 70754
rect 72382 70702 72434 70754
rect 72830 70702 72882 70754
rect 73726 70702 73778 70754
rect 74398 70702 74450 70754
rect 78206 70702 78258 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 71262 70366 71314 70418
rect 69918 70254 69970 70306
rect 3054 70142 3106 70194
rect 69470 70142 69522 70194
rect 70254 70142 70306 70194
rect 70926 70142 70978 70194
rect 71710 70142 71762 70194
rect 76862 70142 76914 70194
rect 2046 70030 2098 70082
rect 3614 70030 3666 70082
rect 77870 70030 77922 70082
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 1822 69246 1874 69298
rect 2718 69246 2770 69298
rect 3950 69246 4002 69298
rect 69358 69246 69410 69298
rect 69694 69246 69746 69298
rect 70254 69246 70306 69298
rect 70590 69246 70642 69298
rect 76526 69246 76578 69298
rect 78094 69246 78146 69298
rect 2158 69134 2210 69186
rect 3054 69134 3106 69186
rect 3502 69134 3554 69186
rect 71150 69134 71202 69186
rect 76190 69134 76242 69186
rect 77310 69134 77362 69186
rect 77758 69134 77810 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 2158 68686 2210 68738
rect 3054 68686 3106 68738
rect 67342 68686 67394 68738
rect 68686 68686 68738 68738
rect 76862 68686 76914 68738
rect 77758 68686 77810 68738
rect 1934 68574 1986 68626
rect 2718 68574 2770 68626
rect 3502 68574 3554 68626
rect 75966 68574 76018 68626
rect 77198 68574 77250 68626
rect 77982 68574 78034 68626
rect 66782 68462 66834 68514
rect 67790 68462 67842 68514
rect 69918 68462 69970 68514
rect 76414 68462 76466 68514
rect 67902 68350 67954 68402
rect 68798 68350 68850 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 2718 67902 2770 67954
rect 67790 67902 67842 67954
rect 68574 67902 68626 67954
rect 69470 67902 69522 67954
rect 70030 67902 70082 67954
rect 66670 67790 66722 67842
rect 67118 67790 67170 67842
rect 77310 67790 77362 67842
rect 77982 67790 78034 67842
rect 1822 67678 1874 67730
rect 2158 67566 2210 67618
rect 3054 67566 3106 67618
rect 67230 67566 67282 67618
rect 67902 67566 67954 67618
rect 68462 67566 68514 67618
rect 69358 67566 69410 67618
rect 77758 67566 77810 67618
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 2158 67118 2210 67170
rect 67566 67118 67618 67170
rect 68462 67118 68514 67170
rect 77758 67118 77810 67170
rect 1934 67006 1986 67058
rect 65774 67006 65826 67058
rect 65998 67006 66050 67058
rect 68238 67006 68290 67058
rect 68910 67006 68962 67058
rect 77310 67006 77362 67058
rect 78094 67006 78146 67058
rect 2606 66894 2658 66946
rect 65886 66894 65938 66946
rect 66222 66894 66274 66946
rect 67118 66894 67170 66946
rect 68350 66894 68402 66946
rect 68686 66894 68738 66946
rect 69358 66894 69410 66946
rect 66446 66782 66498 66834
rect 67006 66782 67058 66834
rect 67342 66782 67394 66834
rect 67902 66782 67954 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 63422 66446 63474 66498
rect 68350 66446 68402 66498
rect 66110 66334 66162 66386
rect 67006 66334 67058 66386
rect 68126 66334 68178 66386
rect 63310 66222 63362 66274
rect 63870 66222 63922 66274
rect 64878 66222 64930 66274
rect 66334 66222 66386 66274
rect 66894 66222 66946 66274
rect 67902 66222 67954 66274
rect 1822 66110 1874 66162
rect 62414 66110 62466 66162
rect 62526 66110 62578 66162
rect 65886 66110 65938 66162
rect 78094 66110 78146 66162
rect 2158 65998 2210 66050
rect 2606 65998 2658 66050
rect 61966 65998 62018 66050
rect 65662 65998 65714 66050
rect 65774 65998 65826 66050
rect 67678 65998 67730 66050
rect 67790 65998 67842 66050
rect 77310 65998 77362 66050
rect 77758 65998 77810 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 66110 65662 66162 65714
rect 2158 65550 2210 65602
rect 64542 65550 64594 65602
rect 65886 65550 65938 65602
rect 77758 65550 77810 65602
rect 1934 65438 1986 65490
rect 61854 65438 61906 65490
rect 65662 65438 65714 65490
rect 65998 65438 66050 65490
rect 68014 65438 68066 65490
rect 68238 65438 68290 65490
rect 68686 65438 68738 65490
rect 77982 65438 78034 65490
rect 2606 65326 2658 65378
rect 61742 65326 61794 65378
rect 62302 65326 62354 65378
rect 67230 65326 67282 65378
rect 68126 65326 68178 65378
rect 68462 65326 68514 65378
rect 77310 65326 77362 65378
rect 64654 65214 64706 65266
rect 65438 65214 65490 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 65550 64766 65602 64818
rect 66446 64766 66498 64818
rect 67006 64766 67058 64818
rect 60734 64654 60786 64706
rect 61406 64654 61458 64706
rect 63534 64654 63586 64706
rect 64206 64654 64258 64706
rect 65774 64654 65826 64706
rect 67454 64654 67506 64706
rect 1822 64542 1874 64594
rect 66334 64542 66386 64594
rect 69358 64542 69410 64594
rect 76638 64542 76690 64594
rect 78094 64542 78146 64594
rect 2158 64430 2210 64482
rect 2606 64430 2658 64482
rect 61518 64430 61570 64482
rect 62078 64430 62130 64482
rect 63646 64430 63698 64482
rect 65102 64430 65154 64482
rect 65214 64430 65266 64482
rect 65326 64430 65378 64482
rect 67790 64430 67842 64482
rect 69694 64430 69746 64482
rect 77310 64430 77362 64482
rect 77758 64430 77810 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 65886 64094 65938 64146
rect 66446 64094 66498 64146
rect 67678 64094 67730 64146
rect 76862 64094 76914 64146
rect 2158 63982 2210 64034
rect 3054 63982 3106 64034
rect 3502 63982 3554 64034
rect 61182 63982 61234 64034
rect 62190 63982 62242 64034
rect 62526 63982 62578 64034
rect 63422 63982 63474 64034
rect 64542 63982 64594 64034
rect 68686 63982 68738 64034
rect 69022 63982 69074 64034
rect 77758 63982 77810 64034
rect 1934 63870 1986 63922
rect 2718 63870 2770 63922
rect 61070 63870 61122 63922
rect 61630 63870 61682 63922
rect 63198 63870 63250 63922
rect 64430 63870 64482 63922
rect 65550 63870 65602 63922
rect 66670 63870 66722 63922
rect 67342 63870 67394 63922
rect 76414 63870 76466 63922
rect 77198 63870 77250 63922
rect 77982 63870 78034 63922
rect 63310 63758 63362 63810
rect 63646 63758 63698 63810
rect 63870 63758 63922 63810
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 63758 63310 63810 63362
rect 2718 63198 2770 63250
rect 63534 63198 63586 63250
rect 64878 63198 64930 63250
rect 67006 63198 67058 63250
rect 61406 63086 61458 63138
rect 61966 63086 62018 63138
rect 63086 63086 63138 63138
rect 1822 62974 1874 63026
rect 59278 62974 59330 63026
rect 77310 62974 77362 63026
rect 78094 62974 78146 63026
rect 2158 62862 2210 62914
rect 3054 62862 3106 62914
rect 59390 62862 59442 62914
rect 59838 62862 59890 62914
rect 61518 62862 61570 62914
rect 63198 62862 63250 62914
rect 63310 62862 63362 62914
rect 65214 62862 65266 62914
rect 66110 62862 66162 62914
rect 77758 62862 77810 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 62638 62526 62690 62578
rect 62862 62526 62914 62578
rect 63646 62526 63698 62578
rect 68798 62526 68850 62578
rect 2158 62414 2210 62466
rect 77758 62414 77810 62466
rect 1934 62302 1986 62354
rect 59838 62302 59890 62354
rect 62526 62302 62578 62354
rect 63870 62302 63922 62354
rect 63982 62302 64034 62354
rect 77982 62302 78034 62354
rect 2606 62190 2658 62242
rect 59726 62190 59778 62242
rect 60286 62190 60338 62242
rect 62750 62190 62802 62242
rect 63758 62190 63810 62242
rect 64318 62190 64370 62242
rect 68238 62190 68290 62242
rect 68350 62190 68402 62242
rect 77310 62190 77362 62242
rect 62190 62078 62242 62130
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 62638 61742 62690 61794
rect 62750 61518 62802 61570
rect 64206 61518 64258 61570
rect 1822 61406 1874 61458
rect 2606 61406 2658 61458
rect 59726 61406 59778 61458
rect 60174 61406 60226 61458
rect 61406 61406 61458 61458
rect 62078 61406 62130 61458
rect 63310 61406 63362 61458
rect 63646 61406 63698 61458
rect 77310 61406 77362 61458
rect 78094 61406 78146 61458
rect 2158 61294 2210 61346
rect 60286 61294 60338 61346
rect 61518 61294 61570 61346
rect 77758 61294 77810 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 62302 60958 62354 61010
rect 65326 60958 65378 61010
rect 2158 60846 2210 60898
rect 59726 60846 59778 60898
rect 60622 60846 60674 60898
rect 62526 60846 62578 60898
rect 64654 60846 64706 60898
rect 77758 60846 77810 60898
rect 1934 60734 1986 60786
rect 57598 60734 57650 60786
rect 59390 60734 59442 60786
rect 60846 60734 60898 60786
rect 61854 60734 61906 60786
rect 63086 60734 63138 60786
rect 78094 60734 78146 60786
rect 2606 60622 2658 60674
rect 57486 60622 57538 60674
rect 58046 60622 58098 60674
rect 58830 60622 58882 60674
rect 60734 60622 60786 60674
rect 61070 60622 61122 60674
rect 62078 60622 62130 60674
rect 62414 60622 62466 60674
rect 77310 60622 77362 60674
rect 61294 60510 61346 60562
rect 64542 60510 64594 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 60398 60062 60450 60114
rect 61518 60062 61570 60114
rect 62078 60062 62130 60114
rect 66670 60062 66722 60114
rect 67230 60062 67282 60114
rect 57374 59950 57426 60002
rect 57934 59950 57986 60002
rect 59950 59950 60002 60002
rect 60622 59950 60674 60002
rect 66558 59950 66610 60002
rect 77982 59950 78034 60002
rect 1822 59838 1874 59890
rect 57486 59838 57538 59890
rect 58718 59838 58770 59890
rect 60174 59838 60226 59890
rect 2158 59726 2210 59778
rect 2606 59726 2658 59778
rect 58830 59726 58882 59778
rect 59278 59726 59330 59778
rect 60062 59726 60114 59778
rect 61406 59726 61458 59778
rect 76638 59726 76690 59778
rect 77310 59726 77362 59778
rect 77758 59726 77810 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 59838 59390 59890 59442
rect 61070 59390 61122 59442
rect 2158 59278 2210 59330
rect 3054 59278 3106 59330
rect 59614 59278 59666 59330
rect 76862 59278 76914 59330
rect 77758 59278 77810 59330
rect 1934 59166 1986 59218
rect 2718 59166 2770 59218
rect 3502 59166 3554 59218
rect 60286 59166 60338 59218
rect 61294 59166 61346 59218
rect 77198 59166 77250 59218
rect 78094 59166 78146 59218
rect 59726 59054 59778 59106
rect 60062 59054 60114 59106
rect 61854 59054 61906 59106
rect 76414 59054 76466 59106
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 2718 58494 2770 58546
rect 59390 58494 59442 58546
rect 60398 58494 60450 58546
rect 56142 58382 56194 58434
rect 56702 58382 56754 58434
rect 58494 58382 58546 58434
rect 59950 58382 60002 58434
rect 77982 58382 78034 58434
rect 1822 58270 1874 58322
rect 57262 58270 57314 58322
rect 57822 58270 57874 58322
rect 77310 58270 77362 58322
rect 2158 58158 2210 58210
rect 3054 58158 3106 58210
rect 56254 58158 56306 58210
rect 57374 58158 57426 58210
rect 58606 58158 58658 58210
rect 59278 58158 59330 58210
rect 77758 58158 77810 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 57598 57822 57650 57874
rect 59502 57822 59554 57874
rect 2158 57710 2210 57762
rect 77758 57710 77810 57762
rect 1934 57598 1986 57650
rect 55134 57598 55186 57650
rect 57822 57598 57874 57650
rect 58830 57598 58882 57650
rect 59278 57598 59330 57650
rect 62750 57598 62802 57650
rect 63198 57598 63250 57650
rect 78094 57598 78146 57650
rect 2606 57486 2658 57538
rect 55022 57486 55074 57538
rect 55582 57486 55634 57538
rect 57710 57486 57762 57538
rect 58046 57486 58098 57538
rect 59054 57486 59106 57538
rect 59390 57486 59442 57538
rect 77310 57486 77362 57538
rect 58270 57374 58322 57426
rect 62638 57374 62690 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 58494 57038 58546 57090
rect 59166 56926 59218 56978
rect 57822 56814 57874 56866
rect 58046 56814 58098 56866
rect 58158 56814 58210 56866
rect 77982 56814 78034 56866
rect 1822 56702 1874 56754
rect 56254 56702 56306 56754
rect 56702 56702 56754 56754
rect 2158 56590 2210 56642
rect 2606 56590 2658 56642
rect 56814 56590 56866 56642
rect 57934 56590 57986 56642
rect 59054 56590 59106 56642
rect 59726 56590 59778 56642
rect 77310 56590 77362 56642
rect 77758 56590 77810 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 56590 56254 56642 56306
rect 57822 56254 57874 56306
rect 2158 56142 2210 56194
rect 57598 56142 57650 56194
rect 77758 56142 77810 56194
rect 1934 56030 1986 56082
rect 52222 56030 52274 56082
rect 55358 56030 55410 56082
rect 55582 56030 55634 56082
rect 55694 56030 55746 56082
rect 56030 56030 56082 56082
rect 58270 56030 58322 56082
rect 78094 56030 78146 56082
rect 2606 55918 2658 55970
rect 52110 55918 52162 55970
rect 52670 55918 52722 55970
rect 54686 55918 54738 55970
rect 55470 55918 55522 55970
rect 56702 55918 56754 55970
rect 57710 55918 57762 55970
rect 58046 55918 58098 55970
rect 58718 55918 58770 55970
rect 77310 55918 77362 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 57598 55470 57650 55522
rect 57822 55470 57874 55522
rect 50318 55358 50370 55410
rect 50878 55358 50930 55410
rect 55582 55358 55634 55410
rect 54126 55246 54178 55298
rect 55134 55246 55186 55298
rect 55806 55246 55858 55298
rect 77982 55246 78034 55298
rect 1822 55134 1874 55186
rect 54350 55134 54402 55186
rect 56926 55134 56978 55186
rect 57262 55134 57314 55186
rect 2158 55022 2210 55074
rect 2606 55022 2658 55074
rect 50430 55022 50482 55074
rect 52446 55022 52498 55074
rect 53566 55022 53618 55074
rect 55246 55022 55298 55074
rect 55358 55022 55410 55074
rect 56254 55022 56306 55074
rect 57710 55022 57762 55074
rect 76638 55022 76690 55074
rect 77310 55022 77362 55074
rect 77758 55022 77810 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 56478 54686 56530 54738
rect 57822 54686 57874 54738
rect 76862 54686 76914 54738
rect 2158 54574 2210 54626
rect 3054 54574 3106 54626
rect 51662 54574 51714 54626
rect 52110 54574 52162 54626
rect 52782 54574 52834 54626
rect 53790 54574 53842 54626
rect 55918 54574 55970 54626
rect 56590 54574 56642 54626
rect 77758 54574 77810 54626
rect 1934 54462 1986 54514
rect 2718 54462 2770 54514
rect 3502 54462 3554 54514
rect 52894 54462 52946 54514
rect 54574 54462 54626 54514
rect 54798 54462 54850 54514
rect 55022 54462 55074 54514
rect 57486 54462 57538 54514
rect 77198 54462 77250 54514
rect 78094 54462 78146 54514
rect 54686 54350 54738 54402
rect 76414 54350 76466 54402
rect 52222 54238 52274 54290
rect 53902 54238 53954 54290
rect 55246 54238 55298 54290
rect 55806 54238 55858 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 54238 53902 54290 53954
rect 57150 53902 57202 53954
rect 57486 53902 57538 53954
rect 2718 53790 2770 53842
rect 54462 53678 54514 53730
rect 54686 53678 54738 53730
rect 54910 53678 54962 53730
rect 55918 53678 55970 53730
rect 56926 53678 56978 53730
rect 57486 53678 57538 53730
rect 1822 53566 1874 53618
rect 2158 53566 2210 53618
rect 52782 53566 52834 53618
rect 53454 53566 53506 53618
rect 55582 53566 55634 53618
rect 78094 53566 78146 53618
rect 3054 53454 3106 53506
rect 52110 53454 52162 53506
rect 53566 53454 53618 53506
rect 54798 53454 54850 53506
rect 77310 53454 77362 53506
rect 77758 53454 77810 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 47742 53118 47794 53170
rect 52670 53118 52722 53170
rect 57822 53118 57874 53170
rect 2158 53006 2210 53058
rect 48302 53006 48354 53058
rect 50318 53006 50370 53058
rect 51886 53006 51938 53058
rect 54350 53006 54402 53058
rect 56702 53006 56754 53058
rect 77758 53006 77810 53058
rect 1934 52894 1986 52946
rect 48414 52894 48466 52946
rect 51662 52894 51714 52946
rect 52894 52894 52946 52946
rect 53902 52894 53954 52946
rect 54574 52894 54626 52946
rect 57486 52894 57538 52946
rect 77982 52894 78034 52946
rect 2606 52782 2658 52834
rect 50206 52782 50258 52834
rect 50766 52782 50818 52834
rect 52782 52782 52834 52834
rect 53118 52782 53170 52834
rect 54126 52782 54178 52834
rect 54462 52782 54514 52834
rect 77310 52782 77362 52834
rect 53342 52670 53394 52722
rect 56590 52670 56642 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 52670 52334 52722 52386
rect 60286 52334 60338 52386
rect 46958 52222 47010 52274
rect 47518 52222 47570 52274
rect 48750 52222 48802 52274
rect 49310 52222 49362 52274
rect 51326 52222 51378 52274
rect 52446 52222 52498 52274
rect 59166 52222 59218 52274
rect 60398 52222 60450 52274
rect 61406 52222 61458 52274
rect 50878 52110 50930 52162
rect 56254 52110 56306 52162
rect 56814 52110 56866 52162
rect 57262 52110 57314 52162
rect 59278 52110 59330 52162
rect 59838 52110 59890 52162
rect 1822 51998 1874 52050
rect 2606 51998 2658 52050
rect 47070 51998 47122 52050
rect 52222 51998 52274 52050
rect 56030 51998 56082 52050
rect 78094 51998 78146 52050
rect 2158 51886 2210 51938
rect 48862 51886 48914 51938
rect 50542 51886 50594 51938
rect 51998 51886 52050 51938
rect 52110 51886 52162 51938
rect 77310 51886 77362 51938
rect 77758 51886 77810 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 51886 51550 51938 51602
rect 53342 51550 53394 51602
rect 56142 51550 56194 51602
rect 57822 51550 57874 51602
rect 2158 51438 2210 51490
rect 52110 51438 52162 51490
rect 53678 51438 53730 51490
rect 77758 51438 77810 51490
rect 1934 51326 1986 51378
rect 52334 51326 52386 51378
rect 52558 51326 52610 51378
rect 56366 51326 56418 51378
rect 57486 51326 57538 51378
rect 77982 51326 78034 51378
rect 2606 51214 2658 51266
rect 51998 51214 52050 51266
rect 55582 51214 55634 51266
rect 77310 51214 77362 51266
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 49198 50654 49250 50706
rect 49646 50654 49698 50706
rect 57150 50654 57202 50706
rect 68686 50654 68738 50706
rect 69358 50654 69410 50706
rect 70030 50654 70082 50706
rect 70702 50654 70754 50706
rect 77310 50654 77362 50706
rect 50766 50542 50818 50594
rect 51102 50542 51154 50594
rect 51662 50542 51714 50594
rect 51774 50542 51826 50594
rect 52334 50542 52386 50594
rect 53678 50542 53730 50594
rect 1822 50430 1874 50482
rect 3054 50430 3106 50482
rect 49758 50430 49810 50482
rect 50654 50430 50706 50482
rect 78094 50430 78146 50482
rect 2158 50318 2210 50370
rect 2718 50318 2770 50370
rect 50430 50318 50482 50370
rect 50542 50318 50594 50370
rect 53454 50318 53506 50370
rect 69470 50318 69522 50370
rect 70142 50318 70194 50370
rect 77758 50318 77810 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 46622 49982 46674 50034
rect 50206 49982 50258 50034
rect 50990 49982 51042 50034
rect 51214 49982 51266 50034
rect 69806 49982 69858 50034
rect 2158 49870 2210 49922
rect 3054 49870 3106 49922
rect 52334 49870 52386 49922
rect 77758 49870 77810 49922
rect 1822 49758 1874 49810
rect 2718 49758 2770 49810
rect 49982 49758 50034 49810
rect 68910 49758 68962 49810
rect 69582 49758 69634 49810
rect 70254 49758 70306 49810
rect 77982 49758 78034 49810
rect 3502 49646 3554 49698
rect 46510 49646 46562 49698
rect 47070 49646 47122 49698
rect 49758 49646 49810 49698
rect 50094 49646 50146 49698
rect 51102 49646 51154 49698
rect 51438 49646 51490 49698
rect 52782 49646 52834 49698
rect 69694 49646 69746 49698
rect 70030 49646 70082 49698
rect 70702 49646 70754 49698
rect 77310 49646 77362 49698
rect 49534 49534 49586 49586
rect 51662 49534 51714 49586
rect 52222 49534 52274 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 48078 49198 48130 49250
rect 47966 49086 48018 49138
rect 48526 49086 48578 49138
rect 49646 49086 49698 49138
rect 68014 49086 68066 49138
rect 68574 49086 68626 49138
rect 69582 49086 69634 49138
rect 70702 49086 70754 49138
rect 3054 48974 3106 49026
rect 49198 48974 49250 49026
rect 49870 48974 49922 49026
rect 50430 48974 50482 49026
rect 69358 48974 69410 49026
rect 2158 48862 2210 48914
rect 50542 48862 50594 48914
rect 78094 48862 78146 48914
rect 3502 48750 3554 48802
rect 49310 48750 49362 48802
rect 49422 48750 49474 48802
rect 51102 48750 51154 48802
rect 68126 48750 68178 48802
rect 69806 48750 69858 48802
rect 69918 48750 69970 48802
rect 70030 48750 70082 48802
rect 76638 48750 76690 48802
rect 77310 48750 77362 48802
rect 77758 48750 77810 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 48526 48414 48578 48466
rect 49758 48414 49810 48466
rect 50318 48414 50370 48466
rect 68910 48414 68962 48466
rect 69358 48414 69410 48466
rect 49870 48302 49922 48354
rect 68798 48302 68850 48354
rect 3054 48190 3106 48242
rect 75070 48190 75122 48242
rect 76974 48190 77026 48242
rect 2046 48078 2098 48130
rect 3614 48078 3666 48130
rect 47294 48078 47346 48130
rect 47854 48078 47906 48130
rect 48414 48078 48466 48130
rect 69918 48078 69970 48130
rect 74622 48078 74674 48130
rect 76078 48078 76130 48130
rect 77870 48078 77922 48130
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 3054 47406 3106 47458
rect 2158 47294 2210 47346
rect 47518 47294 47570 47346
rect 48190 47294 48242 47346
rect 48974 47294 49026 47346
rect 3502 47182 3554 47234
rect 47182 47182 47234 47234
rect 48526 47182 48578 47234
rect 76638 47182 76690 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 46510 46734 46562 46786
rect 47854 46734 47906 46786
rect 3054 46622 3106 46674
rect 46846 46622 46898 46674
rect 47630 46622 47682 46674
rect 75070 46622 75122 46674
rect 77086 46622 77138 46674
rect 2046 46510 2098 46562
rect 3614 46510 3666 46562
rect 46062 46510 46114 46562
rect 48302 46510 48354 46562
rect 74622 46510 74674 46562
rect 76078 46510 76130 46562
rect 77758 46510 77810 46562
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 3054 45838 3106 45890
rect 47742 45838 47794 45890
rect 48078 45838 48130 45890
rect 75294 45838 75346 45890
rect 2158 45726 2210 45778
rect 46174 45726 46226 45778
rect 46846 45726 46898 45778
rect 47182 45726 47234 45778
rect 76190 45726 76242 45778
rect 3502 45614 3554 45666
rect 45838 45614 45890 45666
rect 74734 45614 74786 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 44382 45278 44434 45330
rect 46510 45278 46562 45330
rect 45278 45166 45330 45218
rect 3054 45054 3106 45106
rect 43934 45054 43986 45106
rect 44606 45054 44658 45106
rect 45614 45054 45666 45106
rect 46286 45054 46338 45106
rect 75070 45054 75122 45106
rect 76862 45054 76914 45106
rect 2046 44942 2098 44994
rect 3614 44942 3666 44994
rect 46958 44942 47010 44994
rect 47406 44942 47458 44994
rect 74622 44942 74674 44994
rect 76078 44942 76130 44994
rect 77870 44942 77922 44994
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 3054 44270 3106 44322
rect 46398 44270 46450 44322
rect 2158 44158 2210 44210
rect 43710 44158 43762 44210
rect 44046 44158 44098 44210
rect 44606 44158 44658 44210
rect 45502 44158 45554 44210
rect 45838 44158 45890 44210
rect 3502 44046 3554 44098
rect 46734 44046 46786 44098
rect 76526 44046 76578 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 42926 43710 42978 43762
rect 44382 43710 44434 43762
rect 3054 43486 3106 43538
rect 43262 43486 43314 43538
rect 44158 43486 44210 43538
rect 76862 43486 76914 43538
rect 2046 43374 2098 43426
rect 3614 43374 3666 43426
rect 42478 43374 42530 43426
rect 44830 43374 44882 43426
rect 45278 43374 45330 43426
rect 46062 43374 46114 43426
rect 76414 43374 76466 43426
rect 77870 43374 77922 43426
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 3054 42702 3106 42754
rect 41918 42702 41970 42754
rect 42590 42702 42642 42754
rect 43374 42702 43426 42754
rect 2158 42590 2210 42642
rect 42366 42590 42418 42642
rect 3502 42478 3554 42530
rect 43710 42478 43762 42530
rect 44158 42478 44210 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 41694 42142 41746 42194
rect 43038 42030 43090 42082
rect 3054 41918 3106 41970
rect 42030 41918 42082 41970
rect 42814 41918 42866 41970
rect 75070 41918 75122 41970
rect 76862 41918 76914 41970
rect 77758 41918 77810 41970
rect 2046 41806 2098 41858
rect 3614 41806 3666 41858
rect 43486 41806 43538 41858
rect 43934 41806 43986 41858
rect 74622 41806 74674 41858
rect 76078 41806 76130 41858
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 3054 41134 3106 41186
rect 42142 41134 42194 41186
rect 2158 41022 2210 41074
rect 41022 41022 41074 41074
rect 41358 41022 41410 41074
rect 42366 41022 42418 41074
rect 3502 40910 3554 40962
rect 40014 40910 40066 40962
rect 40574 40910 40626 40962
rect 42814 40910 42866 40962
rect 76638 40910 76690 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 40238 40574 40290 40626
rect 39342 40462 39394 40514
rect 41918 40462 41970 40514
rect 77758 40462 77810 40514
rect 3054 40350 3106 40402
rect 3614 40350 3666 40402
rect 39678 40350 39730 40402
rect 40574 40350 40626 40402
rect 41582 40350 41634 40402
rect 42366 40350 42418 40402
rect 74622 40350 74674 40402
rect 75070 40350 75122 40402
rect 75966 40350 76018 40402
rect 76862 40350 76914 40402
rect 2046 40238 2098 40290
rect 38894 40238 38946 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 77198 39678 77250 39730
rect 2158 39566 2210 39618
rect 3054 39566 3106 39618
rect 75294 39566 75346 39618
rect 3614 39454 3666 39506
rect 38782 39454 38834 39506
rect 39118 39454 39170 39506
rect 39678 39454 39730 39506
rect 40574 39454 40626 39506
rect 40910 39454 40962 39506
rect 76190 39454 76242 39506
rect 38334 39342 38386 39394
rect 40014 39342 40066 39394
rect 41358 39342 41410 39394
rect 74734 39342 74786 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 2158 38894 2210 38946
rect 38334 38894 38386 38946
rect 39790 38894 39842 38946
rect 77758 38894 77810 38946
rect 3054 38782 3106 38834
rect 3614 38782 3666 38834
rect 38670 38782 38722 38834
rect 39566 38782 39618 38834
rect 40686 38782 40738 38834
rect 75070 38782 75122 38834
rect 76862 38782 76914 38834
rect 37886 38670 37938 38722
rect 40238 38670 40290 38722
rect 74622 38670 74674 38722
rect 76078 38670 76130 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 2046 38110 2098 38162
rect 76638 38110 76690 38162
rect 3054 37998 3106 38050
rect 37998 37886 38050 37938
rect 38670 37886 38722 37938
rect 39454 37886 39506 37938
rect 3614 37774 3666 37826
rect 37662 37774 37714 37826
rect 39006 37774 39058 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 2158 37326 2210 37378
rect 36990 37326 37042 37378
rect 38334 37326 38386 37378
rect 77758 37326 77810 37378
rect 3054 37214 3106 37266
rect 37214 37214 37266 37266
rect 37998 37214 38050 37266
rect 75070 37214 75122 37266
rect 76862 37214 76914 37266
rect 3614 37102 3666 37154
rect 36542 37102 36594 37154
rect 38782 37102 38834 37154
rect 74622 37102 74674 37154
rect 76078 37102 76130 37154
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 2046 36542 2098 36594
rect 38334 36542 38386 36594
rect 76638 36542 76690 36594
rect 3054 36430 3106 36482
rect 35870 36318 35922 36370
rect 36654 36318 36706 36370
rect 37550 36318 37602 36370
rect 38782 36318 38834 36370
rect 3614 36206 3666 36258
rect 35310 36206 35362 36258
rect 36318 36206 36370 36258
rect 37886 36206 37938 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 2158 35758 2210 35810
rect 34638 35758 34690 35810
rect 35534 35758 35586 35810
rect 35870 35758 35922 35810
rect 36990 35758 37042 35810
rect 77758 35758 77810 35810
rect 3054 35646 3106 35698
rect 4846 35646 4898 35698
rect 34974 35646 35026 35698
rect 36766 35646 36818 35698
rect 37438 35646 37490 35698
rect 75070 35646 75122 35698
rect 76862 35646 76914 35698
rect 3838 35534 3890 35586
rect 5406 35534 5458 35586
rect 74622 35534 74674 35586
rect 76078 35534 76130 35586
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 2046 34974 2098 35026
rect 3614 34974 3666 35026
rect 77198 34974 77250 35026
rect 3054 34862 3106 34914
rect 33742 34862 33794 34914
rect 34526 34862 34578 34914
rect 35198 34862 35250 34914
rect 36094 34862 36146 34914
rect 75294 34862 75346 34914
rect 34190 34750 34242 34802
rect 36318 34750 36370 34802
rect 76190 34750 76242 34802
rect 4062 34638 4114 34690
rect 35422 34638 35474 34690
rect 36766 34638 36818 34690
rect 74734 34638 74786 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 2158 34190 2210 34242
rect 33630 34190 33682 34242
rect 35086 34190 35138 34242
rect 77758 34190 77810 34242
rect 3054 34078 3106 34130
rect 32958 34078 33010 34130
rect 33966 34078 34018 34130
rect 34862 34078 34914 34130
rect 75070 34078 75122 34130
rect 76862 34078 76914 34130
rect 3614 33966 3666 34018
rect 35646 33966 35698 34018
rect 36094 33966 36146 34018
rect 74622 33966 74674 34018
rect 76078 33966 76130 34018
rect 35982 33854 36034 33906
rect 36206 33854 36258 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 2046 33406 2098 33458
rect 76638 33406 76690 33458
rect 3054 33294 3106 33346
rect 32510 33294 32562 33346
rect 33182 33294 33234 33346
rect 34078 33294 34130 33346
rect 3614 33070 3666 33122
rect 32958 33070 33010 33122
rect 34414 33070 34466 33122
rect 34862 33070 34914 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 34414 32734 34466 32786
rect 2158 32622 2210 32674
rect 32174 32622 32226 32674
rect 33966 32622 34018 32674
rect 77758 32622 77810 32674
rect 3054 32510 3106 32562
rect 32510 32510 32562 32562
rect 33630 32510 33682 32562
rect 74622 32510 74674 32562
rect 75070 32510 75122 32562
rect 76862 32510 76914 32562
rect 3614 32398 3666 32450
rect 31726 32398 31778 32450
rect 76078 32398 76130 32450
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 2046 31838 2098 31890
rect 33406 31838 33458 31890
rect 76638 31838 76690 31890
rect 3054 31726 3106 31778
rect 31166 31614 31218 31666
rect 31950 31614 32002 31666
rect 32622 31614 32674 31666
rect 33854 31614 33906 31666
rect 3614 31502 3666 31554
rect 30718 31502 30770 31554
rect 31614 31502 31666 31554
rect 32958 31502 33010 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 2158 31054 2210 31106
rect 30046 31054 30098 31106
rect 30942 31054 30994 31106
rect 32286 31054 32338 31106
rect 77758 31054 77810 31106
rect 3054 30942 3106 30994
rect 4846 30942 4898 30994
rect 30270 30942 30322 30994
rect 31278 30942 31330 30994
rect 32062 30942 32114 30994
rect 32734 30942 32786 30994
rect 75070 30942 75122 30994
rect 76862 30942 76914 30994
rect 3838 30830 3890 30882
rect 5406 30830 5458 30882
rect 74622 30830 74674 30882
rect 76078 30830 76130 30882
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 32062 30270 32114 30322
rect 77198 30270 77250 30322
rect 2158 30158 2210 30210
rect 3054 30158 3106 30210
rect 3614 30158 3666 30210
rect 75294 30158 75346 30210
rect 30382 30046 30434 30098
rect 31278 30046 31330 30098
rect 31614 30046 31666 30098
rect 76190 30046 76242 30098
rect 4062 29934 4114 29986
rect 29934 29934 29986 29986
rect 30718 29934 30770 29986
rect 74734 29934 74786 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 29598 29598 29650 29650
rect 2158 29486 2210 29538
rect 28702 29486 28754 29538
rect 30830 29486 30882 29538
rect 77758 29486 77810 29538
rect 3054 29374 3106 29426
rect 29038 29374 29090 29426
rect 29934 29374 29986 29426
rect 30494 29374 30546 29426
rect 75070 29374 75122 29426
rect 76862 29374 76914 29426
rect 3614 29262 3666 29314
rect 28254 29262 28306 29314
rect 31278 29262 31330 29314
rect 74622 29262 74674 29314
rect 76078 29262 76130 29314
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 30270 28814 30322 28866
rect 30942 28814 30994 28866
rect 2046 28702 2098 28754
rect 76638 28702 76690 28754
rect 3054 28590 3106 28642
rect 3614 28590 3666 28642
rect 27806 28590 27858 28642
rect 30382 28590 30434 28642
rect 30830 28590 30882 28642
rect 28254 28478 28306 28530
rect 28590 28478 28642 28530
rect 29598 28478 29650 28530
rect 29934 28366 29986 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 2158 27918 2210 27970
rect 27582 27918 27634 27970
rect 28926 27918 28978 27970
rect 77758 27918 77810 27970
rect 3054 27806 3106 27858
rect 27134 27806 27186 27858
rect 27918 27806 27970 27858
rect 28590 27806 28642 27858
rect 29822 27806 29874 27858
rect 75070 27806 75122 27858
rect 76862 27806 76914 27858
rect 3614 27694 3666 27746
rect 29374 27694 29426 27746
rect 74622 27694 74674 27746
rect 76078 27694 76130 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 2046 27134 2098 27186
rect 76638 27134 76690 27186
rect 3054 27022 3106 27074
rect 3614 27022 3666 27074
rect 26462 26910 26514 26962
rect 27246 26910 27298 26962
rect 28030 26910 28082 26962
rect 28814 26910 28866 26962
rect 26910 26798 26962 26850
rect 28366 26798 28418 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 2158 26350 2210 26402
rect 26238 26350 26290 26402
rect 27694 26350 27746 26402
rect 77758 26350 77810 26402
rect 2942 26238 2994 26290
rect 4846 26238 4898 26290
rect 26462 26238 26514 26290
rect 27358 26238 27410 26290
rect 75070 26238 75122 26290
rect 76862 26238 76914 26290
rect 3838 26126 3890 26178
rect 5406 26126 5458 26178
rect 25790 26126 25842 26178
rect 74622 26126 74674 26178
rect 76078 26126 76130 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 2046 25566 2098 25618
rect 77198 25566 77250 25618
rect 3054 25454 3106 25506
rect 25566 25454 25618 25506
rect 27582 25454 27634 25506
rect 75294 25454 75346 25506
rect 4062 25342 4114 25394
rect 24334 25342 24386 25394
rect 24670 25342 24722 25394
rect 25230 25342 25282 25394
rect 26350 25342 26402 25394
rect 27134 25342 27186 25394
rect 76190 25342 76242 25394
rect 3614 25230 3666 25282
rect 26686 25230 26738 25282
rect 74734 25230 74786 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 2158 24782 2210 24834
rect 24110 24782 24162 24834
rect 26126 24782 26178 24834
rect 77758 24782 77810 24834
rect 3054 24670 3106 24722
rect 24446 24670 24498 24722
rect 25902 24670 25954 24722
rect 75070 24670 75122 24722
rect 76862 24670 76914 24722
rect 3614 24558 3666 24610
rect 24894 24558 24946 24610
rect 26574 24558 26626 24610
rect 27022 24558 27074 24610
rect 74622 24558 74674 24610
rect 76078 24558 76130 24610
rect 26350 24446 26402 24498
rect 26574 24446 26626 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 2046 23998 2098 24050
rect 76638 23998 76690 24050
rect 3054 23886 3106 23938
rect 25566 23886 25618 23938
rect 23998 23774 24050 23826
rect 26350 23774 26402 23826
rect 26686 23774 26738 23826
rect 3614 23662 3666 23714
rect 23102 23662 23154 23714
rect 23662 23662 23714 23714
rect 24670 23662 24722 23714
rect 25790 23662 25842 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 26014 23326 26066 23378
rect 2158 23214 2210 23266
rect 22430 23214 22482 23266
rect 23886 23214 23938 23266
rect 77758 23214 77810 23266
rect 3054 23102 3106 23154
rect 22766 23102 22818 23154
rect 23662 23102 23714 23154
rect 24782 23102 24834 23154
rect 75070 23102 75122 23154
rect 76862 23102 76914 23154
rect 3614 22990 3666 23042
rect 24334 22990 24386 23042
rect 25566 22990 25618 23042
rect 74622 22990 74674 23042
rect 76078 22990 76130 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 2046 22430 2098 22482
rect 76638 22430 76690 22482
rect 3054 22318 3106 22370
rect 3614 22206 3666 22258
rect 22094 22206 22146 22258
rect 22430 22206 22482 22258
rect 22990 22206 23042 22258
rect 21646 22094 21698 22146
rect 23326 22094 23378 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 2158 21646 2210 21698
rect 21646 21646 21698 21698
rect 23998 21646 24050 21698
rect 77758 21646 77810 21698
rect 2942 21534 2994 21586
rect 4846 21534 4898 21586
rect 21870 21534 21922 21586
rect 23662 21534 23714 21586
rect 75070 21534 75122 21586
rect 76862 21534 76914 21586
rect 3838 21422 3890 21474
rect 5406 21422 5458 21474
rect 22654 21422 22706 21474
rect 23102 21422 23154 21474
rect 74622 21422 74674 21474
rect 76078 21422 76130 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 2046 20862 2098 20914
rect 77198 20862 77250 20914
rect 3054 20750 3106 20802
rect 75294 20750 75346 20802
rect 4062 20638 4114 20690
rect 21646 20638 21698 20690
rect 21982 20638 22034 20690
rect 23214 20638 23266 20690
rect 76190 20638 76242 20690
rect 3614 20526 3666 20578
rect 20638 20526 20690 20578
rect 22430 20526 22482 20578
rect 23550 20526 23602 20578
rect 74734 20526 74786 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 19966 20190 20018 20242
rect 2158 20078 2210 20130
rect 21198 20078 21250 20130
rect 77758 20078 77810 20130
rect 3054 19966 3106 20018
rect 19518 19966 19570 20018
rect 20302 19966 20354 20018
rect 20862 19966 20914 20018
rect 75070 19966 75122 20018
rect 76862 19966 76914 20018
rect 3614 19854 3666 19906
rect 21758 19854 21810 19906
rect 22206 19854 22258 19906
rect 22878 19854 22930 19906
rect 74622 19854 74674 19906
rect 76078 19854 76130 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 2046 19294 2098 19346
rect 76638 19294 76690 19346
rect 3054 19182 3106 19234
rect 20526 19182 20578 19234
rect 18958 19070 19010 19122
rect 19518 19070 19570 19122
rect 19854 19070 19906 19122
rect 21646 19070 21698 19122
rect 21982 19070 22034 19122
rect 3614 18958 3666 19010
rect 18174 18958 18226 19010
rect 18622 18958 18674 19010
rect 20750 18958 20802 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 21534 18622 21586 18674
rect 56254 18622 56306 18674
rect 2158 18510 2210 18562
rect 18622 18510 18674 18562
rect 21086 18510 21138 18562
rect 55582 18510 55634 18562
rect 3054 18398 3106 18450
rect 18958 18398 19010 18450
rect 20750 18398 20802 18450
rect 55806 18398 55858 18450
rect 56030 18398 56082 18450
rect 56254 18398 56306 18450
rect 75070 18398 75122 18450
rect 76862 18398 76914 18450
rect 77758 18398 77810 18450
rect 3614 18286 3666 18338
rect 18174 18286 18226 18338
rect 19630 18286 19682 18338
rect 20078 18286 20130 18338
rect 54574 18286 54626 18338
rect 55022 18286 55074 18338
rect 74622 18286 74674 18338
rect 76078 18286 76130 18338
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 20526 17838 20578 17890
rect 20750 17838 20802 17890
rect 56142 17838 56194 17890
rect 2046 17726 2098 17778
rect 21982 17726 22034 17778
rect 26126 17726 26178 17778
rect 55582 17726 55634 17778
rect 3054 17614 3106 17666
rect 20078 17614 20130 17666
rect 20302 17614 20354 17666
rect 76638 17614 76690 17666
rect 18062 17502 18114 17554
rect 18622 17502 18674 17554
rect 18958 17502 19010 17554
rect 20862 17502 20914 17554
rect 21534 17502 21586 17554
rect 25790 17502 25842 17554
rect 27022 17502 27074 17554
rect 54798 17502 54850 17554
rect 55470 17502 55522 17554
rect 56030 17502 56082 17554
rect 3614 17390 3666 17442
rect 16382 17390 16434 17442
rect 17166 17390 17218 17442
rect 17726 17390 17778 17442
rect 19406 17390 19458 17442
rect 26014 17390 26066 17442
rect 26574 17390 26626 17442
rect 53566 17390 53618 17442
rect 54014 17390 54066 17442
rect 55022 17390 55074 17442
rect 55246 17390 55298 17442
rect 56590 17390 56642 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 19854 17054 19906 17106
rect 20302 17054 20354 17106
rect 20750 17054 20802 17106
rect 22990 17054 23042 17106
rect 74622 17054 74674 17106
rect 2158 16942 2210 16994
rect 15710 16942 15762 16994
rect 16606 16942 16658 16994
rect 18622 16942 18674 16994
rect 25790 16942 25842 16994
rect 26014 16942 26066 16994
rect 77758 16942 77810 16994
rect 3054 16830 3106 16882
rect 4846 16830 4898 16882
rect 5406 16830 5458 16882
rect 15934 16830 15986 16882
rect 16942 16830 16994 16882
rect 18286 16830 18338 16882
rect 19518 16830 19570 16882
rect 21534 16830 21586 16882
rect 21870 16830 21922 16882
rect 22990 16830 23042 16882
rect 24446 16830 24498 16882
rect 24894 16830 24946 16882
rect 25678 16830 25730 16882
rect 26238 16830 26290 16882
rect 26686 16830 26738 16882
rect 54462 16830 54514 16882
rect 75070 16830 75122 16882
rect 75966 16830 76018 16882
rect 76862 16830 76914 16882
rect 3838 16718 3890 16770
rect 17726 16718 17778 16770
rect 22318 16718 22370 16770
rect 23326 16718 23378 16770
rect 23550 16718 23602 16770
rect 23102 16606 23154 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 16942 16270 16994 16322
rect 17726 16270 17778 16322
rect 18510 16270 18562 16322
rect 22878 16270 22930 16322
rect 23214 16270 23266 16322
rect 2046 16158 2098 16210
rect 3614 16158 3666 16210
rect 16830 16158 16882 16210
rect 18958 16158 19010 16210
rect 77198 16158 77250 16210
rect 3054 16046 3106 16098
rect 18286 16046 18338 16098
rect 18734 16046 18786 16098
rect 19070 16046 19122 16098
rect 22654 16046 22706 16098
rect 75294 16046 75346 16098
rect 15710 15934 15762 15986
rect 16046 15934 16098 15986
rect 19630 15934 19682 15986
rect 76190 15934 76242 15986
rect 4062 15822 4114 15874
rect 17278 15822 17330 15874
rect 17726 15822 17778 15874
rect 19966 15822 20018 15874
rect 23886 15822 23938 15874
rect 74734 15822 74786 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 19294 15486 19346 15538
rect 2158 15374 2210 15426
rect 14702 15374 14754 15426
rect 55918 15374 55970 15426
rect 77758 15374 77810 15426
rect 3054 15262 3106 15314
rect 15038 15262 15090 15314
rect 55022 15262 55074 15314
rect 55582 15262 55634 15314
rect 75070 15262 75122 15314
rect 76862 15262 76914 15314
rect 3614 15150 3666 15202
rect 15486 15150 15538 15202
rect 16270 15150 16322 15202
rect 17054 15150 17106 15202
rect 17726 15150 17778 15202
rect 18174 15150 18226 15202
rect 74622 15150 74674 15202
rect 76078 15150 76130 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 54798 14702 54850 14754
rect 2046 14590 2098 14642
rect 53902 14590 53954 14642
rect 76638 14590 76690 14642
rect 3054 14478 3106 14530
rect 55022 14478 55074 14530
rect 55246 14478 55298 14530
rect 55918 14478 55970 14530
rect 56590 14478 56642 14530
rect 14366 14366 14418 14418
rect 14814 14366 14866 14418
rect 53454 14366 53506 14418
rect 56142 14366 56194 14418
rect 3614 14254 3666 14306
rect 14030 14254 14082 14306
rect 55134 14254 55186 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 2158 13806 2210 13858
rect 12462 13806 12514 13858
rect 13358 13806 13410 13858
rect 55582 13806 55634 13858
rect 57822 13806 57874 13858
rect 77758 13806 77810 13858
rect 3054 13694 3106 13746
rect 12014 13694 12066 13746
rect 12798 13694 12850 13746
rect 13694 13694 13746 13746
rect 55246 13694 55298 13746
rect 56702 13694 56754 13746
rect 57486 13694 57538 13746
rect 74622 13694 74674 13746
rect 75070 13694 75122 13746
rect 76862 13694 76914 13746
rect 3614 13582 3666 13634
rect 14142 13582 14194 13634
rect 54350 13582 54402 13634
rect 76078 13582 76130 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 2046 13022 2098 13074
rect 54910 13022 54962 13074
rect 76638 13022 76690 13074
rect 3054 12910 3106 12962
rect 3614 12686 3666 12738
rect 12014 12686 12066 12738
rect 13022 12686 13074 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 2158 12238 2210 12290
rect 11342 12238 11394 12290
rect 12238 12238 12290 12290
rect 13582 12238 13634 12290
rect 77758 12238 77810 12290
rect 3054 12126 3106 12178
rect 4846 12126 4898 12178
rect 11678 12126 11730 12178
rect 12574 12126 12626 12178
rect 13246 12126 13298 12178
rect 14030 12126 14082 12178
rect 75070 12126 75122 12178
rect 76862 12126 76914 12178
rect 3838 12014 3890 12066
rect 74622 12014 74674 12066
rect 76078 12014 76130 12066
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 2046 11454 2098 11506
rect 3614 11454 3666 11506
rect 4062 11454 4114 11506
rect 77198 11454 77250 11506
rect 3054 11342 3106 11394
rect 75294 11342 75346 11394
rect 10782 11230 10834 11282
rect 11118 11230 11170 11282
rect 11678 11230 11730 11282
rect 12574 11230 12626 11282
rect 12910 11230 12962 11282
rect 76190 11230 76242 11282
rect 12014 11118 12066 11170
rect 74734 11118 74786 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 2158 10670 2210 10722
rect 10110 10670 10162 10722
rect 11454 10670 11506 10722
rect 77758 10670 77810 10722
rect 3054 10558 3106 10610
rect 10446 10558 10498 10610
rect 11118 10558 11170 10610
rect 75070 10558 75122 10610
rect 76862 10558 76914 10610
rect 12238 10446 12290 10498
rect 74622 10446 74674 10498
rect 76078 10446 76130 10498
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 2046 9886 2098 9938
rect 76638 9886 76690 9938
rect 3054 9774 3106 9826
rect 9662 9774 9714 9826
rect 9438 9662 9490 9714
rect 10558 9662 10610 9714
rect 10894 9550 10946 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 2158 9102 2210 9154
rect 8654 9102 8706 9154
rect 10222 9102 10274 9154
rect 77758 9102 77810 9154
rect 3054 8990 3106 9042
rect 8990 8990 9042 9042
rect 9886 8990 9938 9042
rect 74622 8990 74674 9042
rect 75070 8990 75122 9042
rect 76862 8990 76914 9042
rect 76078 8878 76130 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 2046 8318 2098 8370
rect 76638 8318 76690 8370
rect 3054 8206 3106 8258
rect 7982 8094 8034 8146
rect 8318 8094 8370 8146
rect 9102 8094 9154 8146
rect 9438 7982 9490 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 2158 7534 2210 7586
rect 6526 7534 6578 7586
rect 7422 7534 7474 7586
rect 8766 7534 8818 7586
rect 77758 7534 77810 7586
rect 3054 7422 3106 7474
rect 4846 7422 4898 7474
rect 6862 7422 6914 7474
rect 7646 7422 7698 7474
rect 8430 7422 8482 7474
rect 75070 7422 75122 7474
rect 76862 7422 76914 7474
rect 3838 7310 3890 7362
rect 74622 7310 74674 7362
rect 76078 7310 76130 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 77198 6750 77250 6802
rect 2158 6638 2210 6690
rect 3054 6638 3106 6690
rect 7758 6638 7810 6690
rect 75294 6638 75346 6690
rect 5966 6526 6018 6578
rect 6302 6526 6354 6578
rect 6862 6526 6914 6578
rect 8094 6526 8146 6578
rect 76190 6526 76242 6578
rect 7198 6414 7250 6466
rect 74734 6414 74786 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 54238 6078 54290 6130
rect 55022 6078 55074 6130
rect 57374 6078 57426 6130
rect 58158 6078 58210 6130
rect 58718 6078 58770 6130
rect 59166 6078 59218 6130
rect 60286 6078 60338 6130
rect 60734 6078 60786 6130
rect 61182 6078 61234 6130
rect 61630 6078 61682 6130
rect 62078 6078 62130 6130
rect 64206 6078 64258 6130
rect 65326 6078 65378 6130
rect 65774 6078 65826 6130
rect 66222 6078 66274 6130
rect 66782 6078 66834 6130
rect 67678 6078 67730 6130
rect 69022 6078 69074 6130
rect 69470 6078 69522 6130
rect 2158 5966 2210 6018
rect 5294 5966 5346 6018
rect 6750 5966 6802 6018
rect 77758 5966 77810 6018
rect 3054 5854 3106 5906
rect 5630 5854 5682 5906
rect 6414 5854 6466 5906
rect 75070 5854 75122 5906
rect 76862 5854 76914 5906
rect 56366 5742 56418 5794
rect 67230 5742 67282 5794
rect 68126 5742 68178 5794
rect 74622 5742 74674 5794
rect 76078 5742 76130 5794
rect 66222 5630 66274 5682
rect 66558 5630 66610 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 2046 5182 2098 5234
rect 49310 5182 49362 5234
rect 49982 5182 50034 5234
rect 50318 5182 50370 5234
rect 51102 5182 51154 5234
rect 51774 5182 51826 5234
rect 52334 5182 52386 5234
rect 52782 5182 52834 5234
rect 54126 5182 54178 5234
rect 55918 5182 55970 5234
rect 57486 5182 57538 5234
rect 59502 5182 59554 5234
rect 62078 5182 62130 5234
rect 63534 5182 63586 5234
rect 65550 5182 65602 5234
rect 68014 5182 68066 5234
rect 70030 5182 70082 5234
rect 74398 5182 74450 5234
rect 76638 5182 76690 5234
rect 3054 5070 3106 5122
rect 53454 5070 53506 5122
rect 55246 5070 55298 5122
rect 58494 5070 58546 5122
rect 60286 5070 60338 5122
rect 61406 5070 61458 5122
rect 64318 5070 64370 5122
rect 66334 5070 66386 5122
rect 67342 5070 67394 5122
rect 69358 5070 69410 5122
rect 4622 4958 4674 5010
rect 4958 4958 5010 5010
rect 5742 4958 5794 5010
rect 72046 4958 72098 5010
rect 72382 4958 72434 5010
rect 6078 4846 6130 4898
rect 10334 4846 10386 4898
rect 12126 4846 12178 4898
rect 14254 4846 14306 4898
rect 16046 4846 16098 4898
rect 18174 4846 18226 4898
rect 20862 4846 20914 4898
rect 24782 4846 24834 4898
rect 26014 4846 26066 4898
rect 29934 4846 29986 4898
rect 30830 4846 30882 4898
rect 32734 4846 32786 4898
rect 35646 4846 35698 4898
rect 37774 4846 37826 4898
rect 47630 4846 47682 4898
rect 71038 4846 71090 4898
rect 71598 4846 71650 4898
rect 72830 4846 72882 4898
rect 73390 4846 73442 4898
rect 74062 4846 74114 4898
rect 74958 4846 75010 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 5854 4510 5906 4562
rect 6862 4510 6914 4562
rect 9774 4510 9826 4562
rect 11902 4510 11954 4562
rect 13918 4510 13970 4562
rect 15934 4510 15986 4562
rect 18062 4510 18114 4562
rect 20638 4510 20690 4562
rect 21982 4510 22034 4562
rect 24670 4510 24722 4562
rect 26686 4510 26738 4562
rect 29374 4510 29426 4562
rect 30718 4510 30770 4562
rect 32734 4510 32786 4562
rect 35422 4510 35474 4562
rect 37438 4510 37490 4562
rect 39454 4510 39506 4562
rect 41918 4510 41970 4562
rect 44158 4510 44210 4562
rect 46846 4510 46898 4562
rect 48190 4510 48242 4562
rect 71150 4510 71202 4562
rect 71710 4510 71762 4562
rect 73726 4510 73778 4562
rect 74286 4510 74338 4562
rect 75182 4510 75234 4562
rect 47854 4398 47906 4450
rect 5518 4286 5570 4338
rect 7086 4286 7138 4338
rect 9998 4286 10050 4338
rect 11566 4286 11618 4338
rect 13582 4286 13634 4338
rect 15150 4286 15202 4338
rect 15598 4286 15650 4338
rect 17054 4286 17106 4338
rect 17726 4286 17778 4338
rect 19854 4286 19906 4338
rect 20302 4286 20354 4338
rect 21198 4286 21250 4338
rect 21646 4286 21698 4338
rect 23886 4286 23938 4338
rect 24334 4286 24386 4338
rect 25902 4286 25954 4338
rect 26350 4286 26402 4338
rect 29038 4286 29090 4338
rect 30382 4286 30434 4338
rect 32398 4286 32450 4338
rect 35086 4286 35138 4338
rect 37102 4286 37154 4338
rect 38670 4286 38722 4338
rect 39118 4286 39170 4338
rect 41582 4286 41634 4338
rect 43822 4286 43874 4338
rect 46510 4286 46562 4338
rect 49534 4286 49586 4338
rect 51326 4286 51378 4338
rect 53118 4286 53170 4338
rect 55918 4286 55970 4338
rect 56590 4286 56642 4338
rect 57598 4286 57650 4338
rect 59278 4286 59330 4338
rect 61070 4286 61122 4338
rect 63870 4286 63922 4338
rect 64542 4286 64594 4338
rect 65662 4286 65714 4338
rect 67454 4286 67506 4338
rect 69134 4286 69186 4338
rect 70814 4286 70866 4338
rect 72046 4286 72098 4338
rect 72494 4286 72546 4338
rect 73390 4286 73442 4338
rect 74510 4286 74562 4338
rect 75406 4286 75458 4338
rect 5070 4174 5122 4226
rect 6414 4174 6466 4226
rect 7646 4174 7698 4226
rect 8094 4174 8146 4226
rect 8654 4174 8706 4226
rect 8990 4174 9042 4226
rect 10670 4174 10722 4226
rect 11118 4174 11170 4226
rect 12686 4174 12738 4226
rect 13134 4174 13186 4226
rect 14702 4174 14754 4226
rect 16606 4174 16658 4226
rect 18846 4174 18898 4226
rect 19406 4174 19458 4226
rect 22430 4174 22482 4226
rect 22878 4174 22930 4226
rect 23438 4174 23490 4226
rect 27134 4174 27186 4226
rect 27582 4174 27634 4226
rect 28142 4174 28194 4226
rect 28590 4174 28642 4226
rect 29934 4174 29986 4226
rect 31502 4174 31554 4226
rect 31950 4174 32002 4226
rect 33630 4174 33682 4226
rect 34190 4174 34242 4226
rect 34638 4174 34690 4226
rect 36206 4174 36258 4226
rect 36654 4174 36706 4226
rect 38222 4174 38274 4226
rect 39902 4174 39954 4226
rect 40350 4174 40402 4226
rect 40910 4174 40962 4226
rect 42478 4174 42530 4226
rect 42926 4174 42978 4226
rect 43374 4174 43426 4226
rect 44718 4174 44770 4226
rect 45614 4174 45666 4226
rect 46062 4174 46114 4226
rect 47294 4174 47346 4226
rect 48638 4174 48690 4226
rect 50206 4174 50258 4226
rect 52110 4174 52162 4226
rect 53790 4174 53842 4226
rect 55134 4174 55186 4226
rect 58158 4174 58210 4226
rect 59950 4174 60002 4226
rect 61854 4174 61906 4226
rect 63086 4174 63138 4226
rect 66110 4174 66162 4226
rect 67902 4174 67954 4226
rect 69694 4174 69746 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 53454 3614 53506 3666
rect 55246 3614 55298 3666
rect 57374 3614 57426 3666
rect 61294 3614 61346 3666
rect 65214 3614 65266 3666
rect 67006 3614 67058 3666
rect 73166 3614 73218 3666
rect 5966 3502 6018 3554
rect 12574 3502 12626 3554
rect 14702 3502 14754 3554
rect 15598 3502 15650 3554
rect 16606 3502 16658 3554
rect 17950 3502 18002 3554
rect 18622 3502 18674 3554
rect 19406 3502 19458 3554
rect 20638 3502 20690 3554
rect 21646 3502 21698 3554
rect 22766 3502 22818 3554
rect 23438 3502 23490 3554
rect 24558 3502 24610 3554
rect 25790 3502 25842 3554
rect 26686 3502 26738 3554
rect 27470 3502 27522 3554
rect 29598 3502 29650 3554
rect 36206 3502 36258 3554
rect 38222 3502 38274 3554
rect 39342 3502 39394 3554
rect 40238 3502 40290 3554
rect 42702 3502 42754 3554
rect 43598 3502 43650 3554
rect 44942 3502 44994 3554
rect 45838 3502 45890 3554
rect 47070 3502 47122 3554
rect 47966 3502 48018 3554
rect 50094 3502 50146 3554
rect 50878 3502 50930 3554
rect 52782 3502 52834 3554
rect 54686 3502 54738 3554
rect 56702 3502 56754 3554
rect 58494 3502 58546 3554
rect 60622 3502 60674 3554
rect 62414 3502 62466 3554
rect 64542 3502 64594 3554
rect 66558 3502 66610 3554
rect 68462 3502 68514 3554
rect 70590 3502 70642 3554
rect 71262 3502 71314 3554
rect 74286 3502 74338 3554
rect 5070 3390 5122 3442
rect 6190 3390 6242 3442
rect 6750 3390 6802 3442
rect 7086 3390 7138 3442
rect 7646 3390 7698 3442
rect 7982 3390 8034 3442
rect 8542 3390 8594 3442
rect 10110 3390 10162 3442
rect 10670 3390 10722 3442
rect 11902 3390 11954 3442
rect 14030 3390 14082 3442
rect 28142 3390 28194 3442
rect 30606 3390 30658 3442
rect 31502 3390 31554 3442
rect 32398 3390 32450 3442
rect 33630 3390 33682 3442
rect 34190 3390 34242 3442
rect 35422 3390 35474 3442
rect 37550 3390 37602 3442
rect 41358 3390 41410 3442
rect 41806 3390 41858 3442
rect 49198 3390 49250 3442
rect 51550 3390 51602 3442
rect 59390 3390 59442 3442
rect 63310 3390 63362 3442
rect 69358 3390 69410 3442
rect 72718 3390 72770 3442
rect 74958 3390 75010 3442
rect 8878 3278 8930 3330
rect 9774 3278 9826 3330
rect 11006 3278 11058 3330
rect 11566 3278 11618 3330
rect 12798 3278 12850 3330
rect 13694 3278 13746 3330
rect 14926 3278 14978 3330
rect 15822 3278 15874 3330
rect 16382 3278 16434 3330
rect 17614 3278 17666 3330
rect 18846 3278 18898 3330
rect 19742 3278 19794 3330
rect 20302 3278 20354 3330
rect 21870 3278 21922 3330
rect 22430 3278 22482 3330
rect 23662 3278 23714 3330
rect 24222 3278 24274 3330
rect 25454 3278 25506 3330
rect 26350 3278 26402 3330
rect 27246 3278 27298 3330
rect 28478 3278 28530 3330
rect 29374 3278 29426 3330
rect 30270 3278 30322 3330
rect 31166 3278 31218 3330
rect 32062 3278 32114 3330
rect 33294 3278 33346 3330
rect 34526 3278 34578 3330
rect 35086 3278 35138 3330
rect 35982 3278 36034 3330
rect 37214 3278 37266 3330
rect 38446 3278 38498 3330
rect 39006 3278 39058 3330
rect 39902 3278 39954 3330
rect 42142 3278 42194 3330
rect 43038 3278 43090 3330
rect 43934 3278 43986 3330
rect 45278 3278 45330 3330
rect 46174 3278 46226 3330
rect 46734 3278 46786 3330
rect 47630 3278 47682 3330
rect 72382 3278 72434 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 3052 74898 3108 74910
rect 3052 74846 3054 74898
rect 3106 74846 3108 74898
rect 2044 74786 2100 74798
rect 2044 74734 2046 74786
rect 2098 74734 2100 74786
rect 2044 74564 2100 74734
rect 3052 74788 3108 74846
rect 73724 74900 73780 74910
rect 3052 74722 3108 74732
rect 3612 74786 3668 74798
rect 3612 74734 3614 74786
rect 3666 74734 3668 74786
rect 2044 74498 2100 74508
rect 3052 74116 3108 74126
rect 3052 74022 3108 74060
rect 2156 74002 2212 74014
rect 2156 73950 2158 74002
rect 2210 73950 2212 74002
rect 2044 73218 2100 73230
rect 2044 73166 2046 73218
rect 2098 73166 2100 73218
rect 2044 72548 2100 73166
rect 2156 73220 2212 73950
rect 3612 74002 3668 74734
rect 4060 74788 4116 74798
rect 4060 74694 4116 74732
rect 4844 74788 4900 74798
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 3612 73950 3614 74002
rect 3666 73950 3668 74002
rect 3612 73892 3668 73950
rect 4284 74116 4340 74126
rect 4284 74004 4340 74060
rect 4396 74004 4452 74014
rect 4284 74002 4452 74004
rect 4284 73950 4398 74002
rect 4450 73950 4452 74002
rect 4284 73948 4452 73950
rect 3612 73826 3668 73836
rect 3948 73892 4004 73902
rect 3948 73890 4228 73892
rect 3948 73838 3950 73890
rect 4002 73838 4228 73890
rect 3948 73836 4228 73838
rect 3948 73826 4004 73836
rect 2156 73154 2212 73164
rect 3052 73330 3108 73342
rect 3052 73278 3054 73330
rect 3106 73278 3108 73330
rect 3052 73220 3108 73278
rect 3052 73154 3108 73164
rect 3612 73220 3668 73230
rect 3612 73126 3668 73164
rect 2044 72482 2100 72492
rect 3052 72546 3108 72558
rect 3052 72494 3054 72546
rect 3106 72494 3108 72546
rect 2156 72434 2212 72446
rect 2156 72382 2158 72434
rect 2210 72382 2212 72434
rect 2156 71876 2212 72382
rect 3052 72324 3108 72494
rect 3500 72324 3556 72334
rect 3052 72322 3556 72324
rect 3052 72270 3502 72322
rect 3554 72270 3556 72322
rect 3052 72268 3556 72270
rect 2156 71810 2212 71820
rect 3500 71876 3556 72268
rect 3500 71810 3556 71820
rect 3052 71762 3108 71774
rect 3052 71710 3054 71762
rect 3106 71710 3108 71762
rect 2044 71650 2100 71662
rect 2044 71598 2046 71650
rect 2098 71598 2100 71650
rect 2044 71204 2100 71598
rect 3052 71652 3108 71710
rect 3052 71586 3108 71596
rect 3612 71652 3668 71662
rect 3612 71558 3668 71596
rect 2044 71138 2100 71148
rect 3052 70978 3108 70990
rect 3052 70926 3054 70978
rect 3106 70926 3108 70978
rect 2156 70866 2212 70878
rect 2156 70814 2158 70866
rect 2210 70814 2212 70866
rect 2156 70532 2212 70814
rect 3052 70756 3108 70926
rect 3500 70756 3556 70766
rect 3052 70754 3556 70756
rect 3052 70702 3502 70754
rect 3554 70702 3556 70754
rect 3052 70700 3556 70702
rect 2156 70466 2212 70476
rect 3500 70308 3556 70700
rect 3500 70242 3556 70252
rect 3052 70194 3108 70206
rect 3052 70142 3054 70194
rect 3106 70142 3108 70194
rect 2044 70082 2100 70094
rect 2044 70030 2046 70082
rect 2098 70030 2100 70082
rect 2044 69860 2100 70030
rect 3052 70084 3108 70142
rect 3052 70018 3108 70028
rect 3612 70084 3668 70094
rect 3612 69990 3668 70028
rect 2044 69794 2100 69804
rect 1820 69300 1876 69310
rect 1820 67956 1876 69244
rect 2716 69298 2772 69310
rect 2716 69246 2718 69298
rect 2770 69246 2772 69298
rect 2156 69188 2212 69198
rect 2716 69188 2772 69246
rect 3948 69300 4004 69310
rect 3948 69206 4004 69244
rect 2156 69186 2324 69188
rect 2156 69134 2158 69186
rect 2210 69134 2324 69186
rect 2156 69132 2324 69134
rect 2156 69122 2212 69132
rect 2156 68740 2212 68750
rect 2044 68738 2212 68740
rect 2044 68686 2158 68738
rect 2210 68686 2212 68738
rect 2044 68684 2212 68686
rect 1820 67890 1876 67900
rect 1932 68628 1988 68638
rect 1820 67730 1876 67742
rect 1820 67678 1822 67730
rect 1874 67678 1876 67730
rect 1820 67172 1876 67678
rect 1932 67284 1988 68572
rect 2044 67396 2100 68684
rect 2156 68674 2212 68684
rect 2268 67844 2324 69132
rect 2716 69122 2772 69132
rect 3052 69188 3108 69198
rect 3500 69188 3556 69198
rect 3052 69186 3220 69188
rect 3052 69134 3054 69186
rect 3106 69134 3220 69186
rect 3052 69132 3220 69134
rect 3052 69122 3108 69132
rect 3052 68740 3108 68750
rect 3052 68646 3108 68684
rect 2716 68626 2772 68638
rect 2716 68574 2718 68626
rect 2770 68574 2772 68626
rect 2716 68516 2772 68574
rect 2716 67954 2772 68460
rect 3164 68516 3220 69132
rect 3500 69094 3556 69132
rect 3500 68628 3556 68638
rect 3500 68534 3556 68572
rect 3164 68450 3220 68460
rect 2716 67902 2718 67954
rect 2770 67902 2772 67954
rect 2716 67890 2772 67902
rect 2268 67778 2324 67788
rect 2156 67620 2212 67630
rect 2156 67618 2436 67620
rect 2156 67566 2158 67618
rect 2210 67566 2436 67618
rect 2156 67564 2436 67566
rect 2156 67554 2212 67564
rect 2044 67340 2324 67396
rect 1932 67218 1988 67228
rect 2156 67172 2212 67182
rect 1820 66500 1876 67116
rect 2044 67170 2212 67172
rect 2044 67118 2158 67170
rect 2210 67118 2212 67170
rect 2044 67116 2212 67118
rect 1820 66434 1876 66444
rect 1932 67058 1988 67070
rect 1932 67006 1934 67058
rect 1986 67006 1988 67058
rect 1932 66948 1988 67006
rect 1820 66162 1876 66174
rect 1820 66110 1822 66162
rect 1874 66110 1876 66162
rect 1820 65156 1876 66110
rect 1932 65828 1988 66892
rect 1932 65762 1988 65772
rect 1820 65090 1876 65100
rect 1932 65490 1988 65502
rect 1932 65438 1934 65490
rect 1986 65438 1988 65490
rect 1932 65380 1988 65438
rect 2044 65492 2100 67116
rect 2156 67106 2212 67116
rect 2268 66276 2324 67340
rect 2268 66210 2324 66220
rect 2156 66052 2212 66062
rect 2380 66052 2436 67564
rect 3052 67618 3108 67630
rect 3052 67566 3054 67618
rect 3106 67566 3108 67618
rect 3052 67172 3108 67566
rect 3052 67106 3108 67116
rect 2604 66948 2660 66958
rect 2604 66854 2660 66892
rect 2604 66052 2660 66062
rect 2156 66050 2324 66052
rect 2156 65998 2158 66050
rect 2210 65998 2324 66050
rect 2156 65996 2324 65998
rect 2156 65986 2212 65996
rect 2044 65426 2100 65436
rect 2156 65602 2212 65614
rect 2156 65550 2158 65602
rect 2210 65550 2212 65602
rect 1820 64596 1876 64606
rect 1708 64594 1876 64596
rect 1708 64542 1822 64594
rect 1874 64542 1876 64594
rect 1708 64540 1876 64542
rect 1708 63700 1764 64540
rect 1820 64530 1876 64540
rect 1932 64484 1988 65324
rect 2156 64708 2212 65550
rect 1932 64418 1988 64428
rect 2044 64652 2212 64708
rect 2268 64708 2324 65996
rect 2380 65986 2436 65996
rect 2492 66050 2660 66052
rect 2492 65998 2606 66050
rect 2658 65998 2660 66050
rect 2492 65996 2660 65998
rect 2492 65156 2548 65996
rect 2604 65986 2660 65996
rect 2604 65380 2660 65390
rect 2604 65286 2660 65324
rect 2492 65090 2548 65100
rect 1708 63140 1764 63644
rect 1708 63074 1764 63084
rect 1932 64036 1988 64046
rect 1932 63922 1988 63980
rect 1932 63870 1934 63922
rect 1986 63870 1988 63922
rect 1820 63026 1876 63038
rect 1820 62974 1822 63026
rect 1874 62974 1876 63026
rect 1820 61796 1876 62974
rect 1932 62580 1988 63870
rect 2044 63924 2100 64652
rect 2268 64642 2324 64652
rect 2156 64484 2212 64494
rect 2156 64482 2436 64484
rect 2156 64430 2158 64482
rect 2210 64430 2436 64482
rect 2156 64428 2436 64430
rect 2156 64418 2212 64428
rect 2044 63858 2100 63868
rect 2156 64034 2212 64046
rect 2156 63982 2158 64034
rect 2210 63982 2212 64034
rect 2156 63140 2212 63982
rect 2156 63074 2212 63084
rect 2156 62916 2212 62926
rect 2156 62914 2324 62916
rect 2156 62862 2158 62914
rect 2210 62862 2324 62914
rect 2156 62860 2324 62862
rect 2156 62850 2212 62860
rect 1932 62514 1988 62524
rect 2156 62468 2212 62478
rect 2044 62466 2212 62468
rect 2044 62414 2158 62466
rect 2210 62414 2212 62466
rect 2044 62412 2212 62414
rect 1820 61730 1876 61740
rect 1932 62354 1988 62366
rect 1932 62302 1934 62354
rect 1986 62302 1988 62354
rect 1932 62132 1988 62302
rect 1820 61460 1876 61470
rect 1708 61404 1820 61460
rect 1708 60452 1764 61404
rect 1820 61328 1876 61404
rect 1932 61124 1988 62076
rect 1932 61058 1988 61068
rect 1708 60386 1764 60396
rect 1932 60786 1988 60798
rect 1932 60734 1934 60786
rect 1986 60734 1988 60786
rect 1932 60452 1988 60734
rect 2044 60676 2100 62412
rect 2156 62402 2212 62412
rect 2268 61572 2324 62860
rect 2380 62244 2436 64428
rect 2604 64482 2660 64494
rect 2604 64430 2606 64482
rect 2658 64430 2660 64482
rect 2604 63700 2660 64430
rect 3052 64036 3108 64046
rect 3500 64036 3556 64046
rect 3052 64034 3220 64036
rect 3052 63982 3054 64034
rect 3106 63982 3220 64034
rect 3052 63980 3220 63982
rect 3052 63970 3108 63980
rect 2604 63634 2660 63644
rect 2716 63922 2772 63934
rect 2716 63870 2718 63922
rect 2770 63870 2772 63922
rect 2716 63812 2772 63870
rect 2716 63250 2772 63756
rect 2716 63198 2718 63250
rect 2770 63198 2772 63250
rect 2716 63186 2772 63198
rect 3052 62914 3108 62926
rect 3052 62862 3054 62914
rect 3106 62862 3108 62914
rect 2380 62178 2436 62188
rect 2604 62242 2660 62254
rect 2604 62190 2606 62242
rect 2658 62190 2660 62242
rect 2604 62132 2660 62190
rect 2604 62066 2660 62076
rect 3052 61796 3108 62862
rect 3164 62916 3220 63980
rect 3500 63942 3556 63980
rect 3164 62850 3220 62860
rect 3052 61730 3108 61740
rect 2268 61506 2324 61516
rect 2604 61460 2660 61470
rect 2604 61366 2660 61404
rect 2156 61348 2212 61358
rect 2156 61346 2324 61348
rect 2156 61294 2158 61346
rect 2210 61294 2324 61346
rect 2156 61292 2324 61294
rect 2156 61282 2212 61292
rect 2044 60610 2100 60620
rect 2156 60898 2212 60910
rect 2156 60846 2158 60898
rect 2210 60846 2212 60898
rect 1820 59892 1876 59902
rect 1708 59890 1876 59892
rect 1708 59838 1822 59890
rect 1874 59838 1876 59890
rect 1708 59836 1876 59838
rect 1708 58436 1764 59836
rect 1820 59826 1876 59836
rect 1932 59780 1988 60396
rect 2156 60004 2212 60846
rect 2268 60116 2324 61292
rect 2604 60674 2660 60686
rect 2604 60622 2606 60674
rect 2658 60622 2660 60674
rect 2604 60452 2660 60622
rect 2604 60386 2660 60396
rect 2268 60050 2324 60060
rect 2156 59938 2212 59948
rect 1932 59714 1988 59724
rect 2156 59780 2212 59790
rect 2156 59778 2324 59780
rect 2156 59726 2158 59778
rect 2210 59726 2324 59778
rect 2156 59724 2324 59726
rect 2156 59714 2212 59724
rect 2156 59330 2212 59342
rect 2156 59278 2158 59330
rect 2210 59278 2212 59330
rect 1708 58370 1764 58380
rect 1932 59220 1988 59230
rect 1820 58322 1876 58334
rect 1820 58270 1822 58322
rect 1874 58270 1876 58322
rect 1820 57092 1876 58270
rect 1932 57876 1988 59164
rect 2156 58660 2212 59278
rect 2156 58594 2212 58604
rect 2268 58548 2324 59724
rect 2268 58482 2324 58492
rect 2604 59778 2660 59790
rect 2604 59726 2606 59778
rect 2658 59726 2660 59778
rect 2604 58436 2660 59726
rect 3052 59330 3108 59342
rect 3052 59278 3054 59330
rect 3106 59278 3108 59330
rect 2716 59218 2772 59230
rect 2716 59166 2718 59218
rect 2770 59166 2772 59218
rect 2716 59108 2772 59166
rect 2716 58546 2772 59052
rect 2716 58494 2718 58546
rect 2770 58494 2772 58546
rect 2716 58482 2772 58494
rect 2604 58370 2660 58380
rect 3052 58436 3108 59278
rect 3500 59220 3556 59230
rect 3500 59126 3556 59164
rect 3052 58370 3108 58380
rect 3276 58660 3332 58670
rect 2156 58212 2212 58222
rect 2156 58210 2772 58212
rect 2156 58158 2158 58210
rect 2210 58158 2772 58210
rect 2156 58156 2772 58158
rect 2156 58146 2212 58156
rect 1932 57810 1988 57820
rect 2156 57764 2212 57774
rect 2044 57762 2212 57764
rect 2044 57710 2158 57762
rect 2210 57710 2212 57762
rect 2044 57708 2212 57710
rect 1820 57026 1876 57036
rect 1932 57650 1988 57662
rect 1932 57598 1934 57650
rect 1986 57598 1988 57650
rect 1932 56980 1988 57598
rect 1820 56754 1876 56766
rect 1820 56702 1822 56754
rect 1874 56702 1876 56754
rect 1820 56644 1876 56702
rect 1820 55748 1876 56588
rect 1932 56420 1988 56924
rect 1932 56354 1988 56364
rect 1820 55682 1876 55692
rect 1932 56082 1988 56094
rect 1932 56030 1934 56082
rect 1986 56030 1988 56082
rect 1820 55188 1876 55198
rect 1708 55186 1876 55188
rect 1708 55134 1822 55186
rect 1874 55134 1876 55186
rect 1708 55132 1876 55134
rect 1708 53732 1764 55132
rect 1820 55122 1876 55132
rect 1932 55076 1988 56030
rect 2044 55972 2100 57708
rect 2156 57698 2212 57708
rect 2604 57538 2660 57550
rect 2604 57486 2606 57538
rect 2658 57486 2660 57538
rect 2604 56980 2660 57486
rect 2604 56914 2660 56924
rect 2716 56756 2772 58156
rect 3052 58210 3108 58222
rect 3052 58158 3054 58210
rect 3106 58158 3108 58210
rect 3052 57092 3108 58158
rect 3276 57540 3332 58604
rect 3276 57474 3332 57484
rect 3052 57026 3108 57036
rect 2716 56690 2772 56700
rect 2156 56644 2212 56654
rect 2604 56644 2660 56654
rect 2156 56642 2324 56644
rect 2156 56590 2158 56642
rect 2210 56590 2324 56642
rect 2156 56588 2324 56590
rect 2156 56578 2212 56588
rect 2044 55906 2100 55916
rect 2156 56194 2212 56206
rect 2156 56142 2158 56194
rect 2210 56142 2212 56194
rect 2156 55468 2212 56142
rect 1932 55010 1988 55020
rect 2044 55412 2212 55468
rect 2268 55412 2324 56588
rect 2604 56550 2660 56588
rect 2604 55970 2660 55982
rect 2604 55918 2606 55970
rect 2658 55918 2660 55970
rect 2604 55468 2660 55918
rect 2044 54740 2100 55412
rect 2268 55346 2324 55356
rect 2492 55412 2660 55468
rect 2156 55076 2212 55086
rect 2492 55076 2548 55412
rect 2156 55074 2436 55076
rect 2156 55022 2158 55074
rect 2210 55022 2436 55074
rect 2156 55020 2436 55022
rect 2156 55010 2212 55020
rect 2044 54674 2100 54684
rect 2156 54628 2212 54638
rect 2156 54626 2324 54628
rect 2156 54574 2158 54626
rect 2210 54574 2324 54626
rect 2156 54572 2324 54574
rect 2156 54562 2212 54572
rect 1708 53666 1764 53676
rect 1932 54516 1988 54526
rect 1820 53618 1876 53630
rect 1820 53566 1822 53618
rect 1874 53566 1876 53618
rect 1820 53508 1876 53566
rect 1820 52388 1876 53452
rect 1932 53172 1988 54460
rect 2156 53620 2212 53630
rect 2156 53526 2212 53564
rect 2268 53396 2324 54572
rect 2268 53330 2324 53340
rect 1932 53106 1988 53116
rect 2156 53060 2212 53070
rect 2380 53060 2436 55020
rect 2492 55010 2548 55020
rect 2604 55074 2660 55086
rect 2604 55022 2606 55074
rect 2658 55022 2660 55074
rect 2604 53732 2660 55022
rect 3052 54628 3108 54638
rect 3052 54534 3108 54572
rect 2716 54514 2772 54526
rect 2716 54462 2718 54514
rect 2770 54462 2772 54514
rect 2716 54404 2772 54462
rect 3500 54516 3556 54526
rect 3500 54422 3556 54460
rect 2716 53842 2772 54348
rect 2716 53790 2718 53842
rect 2770 53790 2772 53842
rect 2716 53778 2772 53790
rect 2604 53666 2660 53676
rect 3052 53508 3108 53518
rect 3052 53414 3108 53452
rect 2380 53004 2772 53060
rect 2156 52966 2212 53004
rect 1820 52322 1876 52332
rect 1932 52946 1988 52958
rect 1932 52894 1934 52946
rect 1986 52894 1988 52946
rect 1932 52836 1988 52894
rect 2604 52836 2660 52846
rect 1932 52834 2660 52836
rect 1932 52782 2606 52834
rect 2658 52782 2660 52834
rect 1932 52780 2660 52782
rect 1820 52052 1876 52062
rect 1820 51044 1876 51996
rect 1932 51716 1988 52780
rect 2604 52770 2660 52780
rect 2716 52836 2772 53004
rect 2716 52770 2772 52780
rect 2604 52052 2660 52062
rect 2604 51958 2660 51996
rect 2156 51940 2212 51950
rect 2156 51846 2212 51884
rect 1932 51650 1988 51660
rect 2156 51492 2212 51502
rect 2156 51490 2996 51492
rect 2156 51438 2158 51490
rect 2210 51438 2996 51490
rect 2156 51436 2996 51438
rect 2156 51426 2212 51436
rect 1820 50978 1876 50988
rect 1932 51378 1988 51390
rect 1932 51326 1934 51378
rect 1986 51326 1988 51378
rect 1932 51268 1988 51326
rect 2604 51268 2660 51278
rect 1932 51266 2660 51268
rect 1932 51214 2606 51266
rect 2658 51214 2660 51266
rect 1932 51212 2660 51214
rect 1820 50484 1876 50494
rect 1708 50482 1876 50484
rect 1708 50430 1822 50482
rect 1874 50430 1876 50482
rect 1708 50428 1876 50430
rect 1708 50260 1764 50428
rect 1820 50418 1876 50428
rect 1932 50372 1988 51212
rect 2604 51202 2660 51212
rect 1932 50306 1988 50316
rect 2156 50372 2212 50382
rect 2156 50370 2324 50372
rect 2156 50318 2158 50370
rect 2210 50318 2324 50370
rect 2156 50316 2324 50318
rect 2156 50306 2212 50316
rect 1708 49028 1764 50204
rect 2156 49924 2212 49934
rect 2156 49830 2212 49868
rect 1708 48962 1764 48972
rect 1820 49810 1876 49822
rect 1820 49758 1822 49810
rect 1874 49758 1876 49810
rect 1820 49588 1876 49758
rect 1820 48356 1876 49532
rect 1820 48290 1876 48300
rect 2156 48914 2212 48926
rect 2156 48862 2158 48914
rect 2210 48862 2212 48914
rect 2044 48130 2100 48142
rect 2044 48078 2046 48130
rect 2098 48078 2100 48130
rect 2044 47012 2100 48078
rect 2156 47684 2212 48862
rect 2268 48132 2324 50316
rect 2716 50370 2772 50382
rect 2716 50318 2718 50370
rect 2770 50318 2772 50370
rect 2716 49810 2772 50318
rect 2716 49758 2718 49810
rect 2770 49758 2772 49810
rect 2716 49700 2772 49758
rect 2716 49634 2772 49644
rect 2940 49700 2996 51436
rect 4172 50708 4228 73836
rect 4284 72436 4340 73948
rect 4396 73938 4452 73948
rect 4844 73108 4900 74732
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 73388 73890 73444 73902
rect 73388 73838 73390 73890
rect 73442 73838 73444 73890
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 69356 73444 69412 73454
rect 69356 73350 69412 73388
rect 4844 73042 4900 73052
rect 69132 73332 69188 73342
rect 69132 73106 69188 73276
rect 70028 73332 70084 73342
rect 70028 73238 70084 73276
rect 73276 73332 73332 73342
rect 69132 73054 69134 73106
rect 69186 73054 69188 73106
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 4284 72370 4340 72380
rect 69132 72436 69188 73054
rect 69244 73218 69300 73230
rect 69244 73166 69246 73218
rect 69298 73166 69300 73218
rect 69244 73108 69300 73166
rect 69244 73042 69300 73052
rect 71820 73220 71876 73230
rect 69804 72660 69860 72670
rect 69356 72436 69412 72446
rect 69132 72434 69412 72436
rect 69132 72382 69358 72434
rect 69410 72382 69412 72434
rect 69132 72380 69412 72382
rect 68684 72324 68740 72334
rect 69132 72324 69188 72380
rect 69356 72370 69412 72380
rect 69468 72436 69524 72446
rect 69468 72342 69524 72380
rect 68684 72322 69188 72324
rect 68684 72270 68686 72322
rect 68738 72270 69188 72322
rect 68684 72268 69188 72270
rect 68684 72258 68740 72268
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 67340 68740 67396 68750
rect 67340 68646 67396 68684
rect 67676 68740 67732 68750
rect 66780 68516 66836 68526
rect 66780 68422 66836 68460
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 67676 67956 67732 68684
rect 68684 68740 68740 68750
rect 68684 68646 68740 68684
rect 67788 68516 67844 68526
rect 67788 68422 67844 68460
rect 67900 68404 67956 68414
rect 67900 68402 68404 68404
rect 67900 68350 67902 68402
rect 67954 68350 68404 68402
rect 67900 68348 68404 68350
rect 67900 68338 67956 68348
rect 67788 67956 67844 67966
rect 67676 67954 67844 67956
rect 67676 67902 67790 67954
rect 67842 67902 67844 67954
rect 67676 67900 67844 67902
rect 67788 67890 67844 67900
rect 66668 67844 66724 67854
rect 66668 67750 66724 67788
rect 67116 67844 67172 67854
rect 67116 67750 67172 67788
rect 67228 67618 67284 67630
rect 67228 67566 67230 67618
rect 67282 67566 67284 67618
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 67228 67228 67284 67566
rect 67900 67618 67956 67630
rect 67900 67566 67902 67618
rect 67954 67566 67956 67618
rect 67900 67228 67956 67566
rect 67228 67172 67396 67228
rect 63420 67060 63476 67070
rect 65772 67060 65828 67070
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 63420 66498 63476 67004
rect 63420 66446 63422 66498
rect 63474 66446 63476 66498
rect 63420 66434 63476 66446
rect 65660 67058 65828 67060
rect 65660 67006 65774 67058
rect 65826 67006 65828 67058
rect 65660 67004 65828 67006
rect 63308 66276 63364 66286
rect 63308 66182 63364 66220
rect 63868 66276 63924 66286
rect 63868 66182 63924 66220
rect 64540 66276 64596 66286
rect 62412 66162 62468 66174
rect 62412 66110 62414 66162
rect 62466 66110 62468 66162
rect 61964 66052 62020 66062
rect 61964 65958 62020 65996
rect 62412 66052 62468 66110
rect 62524 66164 62580 66174
rect 62524 66070 62580 66108
rect 62412 65986 62468 65996
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 61852 65604 61908 65614
rect 61852 65490 61908 65548
rect 64540 65602 64596 66220
rect 64876 66276 64932 66286
rect 64876 66182 64932 66220
rect 65660 66052 65716 67004
rect 65772 66994 65828 67004
rect 65996 67060 66052 67070
rect 65996 66966 66052 67004
rect 65884 66946 65940 66958
rect 65884 66894 65886 66946
rect 65938 66894 65940 66946
rect 65884 66836 65940 66894
rect 66220 66948 66276 66958
rect 67116 66948 67172 66958
rect 66220 66946 66388 66948
rect 66220 66894 66222 66946
rect 66274 66894 66388 66946
rect 66220 66892 66388 66894
rect 66220 66882 66276 66892
rect 65772 66780 65940 66836
rect 65772 66388 65828 66780
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 66332 66500 66388 66892
rect 67116 66854 67172 66892
rect 66444 66836 66500 66846
rect 67004 66836 67060 66846
rect 66444 66834 67060 66836
rect 66444 66782 66446 66834
rect 66498 66782 67006 66834
rect 67058 66782 67060 66834
rect 66444 66780 67060 66782
rect 66444 66770 66500 66780
rect 67004 66770 67060 66780
rect 67340 66834 67396 67172
rect 67340 66782 67342 66834
rect 67394 66782 67396 66834
rect 67340 66770 67396 66782
rect 67564 67172 67620 67182
rect 67900 67172 68068 67228
rect 66108 66444 66388 66500
rect 65772 66332 66052 66388
rect 65884 66164 65940 66174
rect 65884 66070 65940 66108
rect 65660 65986 65716 65996
rect 65772 66050 65828 66062
rect 65772 65998 65774 66050
rect 65826 65998 65828 66050
rect 64540 65550 64542 65602
rect 64594 65550 64596 65602
rect 64540 65538 64596 65550
rect 65660 65828 65716 65838
rect 65660 65492 65716 65772
rect 61852 65438 61854 65490
rect 61906 65438 61908 65490
rect 61852 65426 61908 65438
rect 65548 65490 65716 65492
rect 65548 65438 65662 65490
rect 65714 65438 65716 65490
rect 65548 65436 65716 65438
rect 61740 65380 61796 65390
rect 61740 65286 61796 65324
rect 62300 65380 62356 65390
rect 62300 65286 62356 65324
rect 64652 65268 64708 65278
rect 65436 65268 65492 65278
rect 64652 65266 65492 65268
rect 64652 65214 64654 65266
rect 64706 65214 65438 65266
rect 65490 65214 65492 65266
rect 64652 65212 65492 65214
rect 64652 65202 64708 65212
rect 65436 65202 65492 65212
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 65548 64818 65604 65436
rect 65660 65426 65716 65436
rect 65772 64932 65828 65998
rect 65996 65716 66052 66332
rect 66108 66386 66164 66444
rect 66108 66334 66110 66386
rect 66162 66334 66164 66386
rect 66108 66322 66164 66334
rect 65996 65650 66052 65660
rect 66108 65940 66164 65950
rect 66108 65714 66164 65884
rect 66220 65828 66276 66444
rect 67004 66388 67060 66398
rect 67004 66294 67060 66332
rect 67564 66388 67620 67116
rect 67564 66322 67620 66332
rect 67676 67060 67732 67070
rect 66332 66276 66388 66286
rect 66892 66276 66948 66286
rect 66332 66274 66948 66276
rect 66332 66222 66334 66274
rect 66386 66222 66894 66274
rect 66946 66222 66948 66274
rect 66332 66220 66948 66222
rect 66332 66210 66388 66220
rect 66892 66210 66948 66220
rect 67676 66050 67732 67004
rect 67900 66834 67956 66846
rect 67900 66782 67902 66834
rect 67954 66782 67956 66834
rect 67900 66274 67956 66782
rect 67900 66222 67902 66274
rect 67954 66222 67956 66274
rect 67900 66210 67956 66222
rect 67676 65998 67678 66050
rect 67730 65998 67732 66050
rect 66668 65940 66724 65950
rect 66220 65762 66276 65772
rect 66444 65828 66500 65838
rect 66108 65662 66110 65714
rect 66162 65662 66164 65714
rect 66108 65650 66164 65662
rect 65884 65604 65940 65614
rect 65884 65510 65940 65548
rect 65996 65492 66052 65502
rect 65996 65490 66388 65492
rect 65996 65438 65998 65490
rect 66050 65438 66388 65490
rect 65996 65436 66388 65438
rect 65996 65426 66052 65436
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 66332 64932 66388 65436
rect 65548 64766 65550 64818
rect 65602 64766 65604 64818
rect 60732 64708 60788 64718
rect 60732 64614 60788 64652
rect 61404 64708 61460 64718
rect 61404 64614 61460 64652
rect 63532 64708 63588 64718
rect 63532 64614 63588 64652
rect 64204 64708 64260 64718
rect 64204 64614 64260 64652
rect 61516 64484 61572 64494
rect 61516 64390 61572 64428
rect 62076 64484 62132 64494
rect 63644 64484 63700 64494
rect 62076 64482 62244 64484
rect 62076 64430 62078 64482
rect 62130 64430 62244 64482
rect 62076 64428 62244 64430
rect 62076 64418 62132 64428
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 59500 64148 59556 64158
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 59276 63026 59332 63038
rect 59276 62974 59278 63026
rect 59330 62974 59332 63026
rect 59276 62916 59332 62974
rect 59276 62850 59332 62860
rect 59388 62914 59444 62926
rect 59388 62862 59390 62914
rect 59442 62862 59444 62914
rect 59388 62804 59444 62862
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 59388 62738 59444 62748
rect 50556 62682 50820 62692
rect 59500 62188 59556 64092
rect 62188 64148 62244 64428
rect 63644 64482 63812 64484
rect 63644 64430 63646 64482
rect 63698 64430 63812 64482
rect 63644 64428 63812 64430
rect 63644 64418 63700 64428
rect 61180 64036 61236 64046
rect 61180 63942 61236 63980
rect 62188 64034 62244 64092
rect 62188 63982 62190 64034
rect 62242 63982 62244 64034
rect 62188 63970 62244 63982
rect 62524 64034 62580 64046
rect 62524 63982 62526 64034
rect 62578 63982 62580 64034
rect 61068 63924 61124 63934
rect 61068 63830 61124 63868
rect 61628 63924 61684 63934
rect 61628 63830 61684 63868
rect 62524 63812 62580 63982
rect 63420 64036 63476 64046
rect 63420 63942 63476 63980
rect 61404 63140 61460 63150
rect 61404 63046 61460 63084
rect 61964 63140 62020 63150
rect 61964 63046 62020 63084
rect 59836 62916 59892 62926
rect 59836 62822 59892 62860
rect 61516 62914 61572 62926
rect 61516 62862 61518 62914
rect 61570 62862 61572 62914
rect 61516 62580 61572 62862
rect 61516 62514 61572 62524
rect 59836 62356 59892 62366
rect 59836 62262 59892 62300
rect 62524 62354 62580 63756
rect 63196 63922 63252 63934
rect 63196 63870 63198 63922
rect 63250 63870 63252 63922
rect 63084 63140 63140 63150
rect 63196 63140 63252 63870
rect 63532 63924 63588 63934
rect 63308 63810 63364 63822
rect 63308 63758 63310 63810
rect 63362 63758 63364 63810
rect 63308 63252 63364 63758
rect 63420 63812 63476 63822
rect 63420 63252 63476 63756
rect 63532 63476 63588 63868
rect 63644 63812 63700 63822
rect 63756 63812 63812 64428
rect 65100 64482 65156 64494
rect 65100 64430 65102 64482
rect 65154 64430 65156 64482
rect 65100 64372 65156 64430
rect 65100 64306 65156 64316
rect 65212 64482 65268 64494
rect 65212 64430 65214 64482
rect 65266 64430 65268 64482
rect 64540 64260 64596 64270
rect 64540 64034 64596 64204
rect 64540 63982 64542 64034
rect 64594 63982 64596 64034
rect 64540 63970 64596 63982
rect 64876 64260 64932 64270
rect 64428 63924 64484 63934
rect 64428 63830 64484 63868
rect 63868 63812 63924 63822
rect 63756 63810 63924 63812
rect 63756 63758 63870 63810
rect 63922 63758 63924 63810
rect 63756 63756 63924 63758
rect 63644 63718 63700 63756
rect 63868 63746 63924 63756
rect 63980 63812 64036 63822
rect 63532 63420 63812 63476
rect 63756 63362 63812 63420
rect 63756 63310 63758 63362
rect 63810 63310 63812 63362
rect 63756 63298 63812 63310
rect 63532 63252 63588 63262
rect 63420 63250 63588 63252
rect 63420 63198 63534 63250
rect 63586 63198 63588 63250
rect 63420 63196 63588 63198
rect 63308 63186 63364 63196
rect 63532 63186 63588 63196
rect 62860 63138 63196 63140
rect 62860 63086 63086 63138
rect 63138 63086 63196 63138
rect 62860 63084 63196 63086
rect 62636 62580 62692 62590
rect 62636 62486 62692 62524
rect 62860 62578 62916 63084
rect 62860 62526 62862 62578
rect 62914 62526 62916 62578
rect 62860 62514 62916 62526
rect 62524 62302 62526 62354
rect 62578 62302 62580 62354
rect 62524 62290 62580 62302
rect 59388 62132 59556 62188
rect 59724 62244 59780 62254
rect 59724 62150 59780 62188
rect 60284 62244 60340 62254
rect 60284 62150 60340 62188
rect 62748 62242 62804 62254
rect 62748 62190 62750 62242
rect 62802 62190 62804 62242
rect 62748 62188 62804 62190
rect 63084 62188 63140 63084
rect 63196 63074 63252 63084
rect 63644 63140 63700 63150
rect 62188 62132 62244 62142
rect 62748 62132 62916 62188
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 57596 60788 57652 60798
rect 57596 60694 57652 60732
rect 59388 60786 59444 62132
rect 62188 62130 62692 62132
rect 62188 62078 62190 62130
rect 62242 62078 62692 62130
rect 62188 62076 62692 62078
rect 62188 62066 62244 62076
rect 62636 61794 62692 62076
rect 62636 61742 62638 61794
rect 62690 61742 62692 61794
rect 62636 61730 62692 61742
rect 62748 61572 62804 61582
rect 62748 61478 62804 61516
rect 59724 61460 59780 61470
rect 59724 61366 59780 61404
rect 60172 61460 60228 61470
rect 60172 61366 60228 61404
rect 61404 61460 61460 61470
rect 61404 61366 61460 61404
rect 62076 61460 62132 61470
rect 62076 61366 62132 61404
rect 60284 61346 60340 61358
rect 60284 61294 60286 61346
rect 60338 61294 60340 61346
rect 60284 61012 60340 61294
rect 61516 61348 61572 61358
rect 61516 61346 61908 61348
rect 61516 61294 61518 61346
rect 61570 61294 61908 61346
rect 61516 61292 61908 61294
rect 61516 61282 61572 61292
rect 60284 60946 60340 60956
rect 59388 60734 59390 60786
rect 59442 60734 59444 60786
rect 57484 60676 57540 60686
rect 57484 60582 57540 60620
rect 58044 60676 58100 60686
rect 58044 60582 58100 60620
rect 58380 60676 58436 60686
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 57372 60004 57428 60014
rect 57372 59910 57428 59948
rect 57932 60004 57988 60014
rect 57932 59910 57988 59948
rect 57484 59892 57540 59902
rect 57484 59798 57540 59836
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 56140 58436 56196 58446
rect 56140 58342 56196 58380
rect 56700 58436 56756 58446
rect 56700 58342 56756 58380
rect 57260 58324 57316 58334
rect 57260 58230 57316 58268
rect 57820 58324 57876 58334
rect 57820 58230 57876 58268
rect 56252 58210 56308 58222
rect 56252 58158 56254 58210
rect 56306 58158 56308 58210
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 55132 57652 55188 57662
rect 55132 57558 55188 57596
rect 55020 57540 55076 57550
rect 55020 57446 55076 57484
rect 55580 57540 55636 57550
rect 55580 57446 55636 57484
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 56252 56980 56308 58158
rect 57372 58210 57428 58222
rect 57372 58158 57374 58210
rect 57426 58158 57428 58210
rect 57372 57764 57428 58158
rect 57596 57988 57652 57998
rect 57596 57874 57652 57932
rect 57596 57822 57598 57874
rect 57650 57822 57652 57874
rect 57596 57810 57652 57822
rect 57932 57988 57988 57998
rect 57372 57698 57428 57708
rect 57820 57652 57876 57662
rect 57820 57558 57876 57596
rect 57708 57538 57764 57550
rect 57708 57486 57710 57538
rect 57762 57486 57764 57538
rect 57708 56980 57764 57486
rect 56252 56914 56308 56924
rect 57372 56924 57764 56980
rect 56252 56756 56308 56766
rect 56252 56662 56308 56700
rect 56700 56756 56756 56766
rect 56700 56662 56756 56700
rect 56812 56642 56868 56654
rect 56812 56590 56814 56642
rect 56866 56590 56868 56642
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 56028 56364 56644 56420
rect 52220 56084 52276 56094
rect 52220 55990 52276 56028
rect 55356 56082 55412 56094
rect 55356 56030 55358 56082
rect 55410 56030 55412 56082
rect 52108 55972 52164 55982
rect 52108 55878 52164 55916
rect 52668 55972 52724 55982
rect 52668 55878 52724 55916
rect 54684 55970 54740 55982
rect 54684 55918 54686 55970
rect 54738 55918 54740 55970
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 50316 55412 50372 55422
rect 50316 55318 50372 55356
rect 50876 55412 50932 55422
rect 50876 55318 50932 55356
rect 52332 55300 52388 55310
rect 50428 55076 50484 55086
rect 50428 54982 50484 55020
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 51660 54628 51716 54638
rect 51660 54534 51716 54572
rect 52108 54628 52164 54638
rect 52108 54534 52164 54572
rect 52220 54290 52276 54302
rect 52220 54238 52222 54290
rect 52274 54238 52276 54290
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 52220 53732 52276 54238
rect 52220 53666 52276 53676
rect 46956 53620 47012 53630
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 46956 52276 47012 53564
rect 47740 53508 47796 53518
rect 47740 53170 47796 53452
rect 47740 53118 47742 53170
rect 47794 53118 47796 53170
rect 47740 53106 47796 53118
rect 48300 53508 48356 53518
rect 52108 53508 52164 53518
rect 52332 53508 52388 55244
rect 54124 55300 54180 55310
rect 54124 55206 54180 55244
rect 54684 55300 54740 55918
rect 54684 55234 54740 55244
rect 55132 55300 55188 55310
rect 55356 55300 55412 56030
rect 55580 56084 55636 56094
rect 55580 55990 55636 56028
rect 55692 56082 55748 56094
rect 55692 56030 55694 56082
rect 55746 56030 55748 56082
rect 55132 55298 55412 55300
rect 55132 55246 55134 55298
rect 55186 55246 55412 55298
rect 55132 55244 55412 55246
rect 55468 55970 55524 55982
rect 55468 55918 55470 55970
rect 55522 55918 55524 55970
rect 54348 55188 54404 55198
rect 52444 55074 52500 55086
rect 52444 55022 52446 55074
rect 52498 55022 52500 55074
rect 52444 54740 52500 55022
rect 53564 55074 53620 55086
rect 53564 55022 53566 55074
rect 53618 55022 53620 55074
rect 52444 54674 52500 54684
rect 52780 54740 52836 54750
rect 52780 54626 52836 54684
rect 53564 54740 53620 55022
rect 53564 54674 53620 54684
rect 53788 54740 53844 54750
rect 52780 54574 52782 54626
rect 52834 54574 52836 54626
rect 52780 54562 52836 54574
rect 53788 54626 53844 54684
rect 53788 54574 53790 54626
rect 53842 54574 53844 54626
rect 53788 54562 53844 54574
rect 52892 54516 52948 54526
rect 52892 54422 52948 54460
rect 53900 54292 53956 54302
rect 53900 54290 54292 54292
rect 53900 54238 53902 54290
rect 53954 54238 54292 54290
rect 53900 54236 54292 54238
rect 53900 54226 53956 54236
rect 54236 53954 54292 54236
rect 54236 53902 54238 53954
rect 54290 53902 54292 53954
rect 54236 53890 54292 53902
rect 54348 53732 54404 55132
rect 55132 54852 55188 55244
rect 54572 54796 55188 54852
rect 55244 55074 55300 55086
rect 55244 55022 55246 55074
rect 55298 55022 55300 55074
rect 54572 54514 54628 54796
rect 54572 54462 54574 54514
rect 54626 54462 54628 54514
rect 54572 54450 54628 54462
rect 54796 54516 54852 54526
rect 54796 54422 54852 54460
rect 54684 54404 54740 54414
rect 54684 54310 54740 54348
rect 54572 54180 54628 54190
rect 54460 53732 54516 53742
rect 54348 53730 54516 53732
rect 54348 53678 54462 53730
rect 54514 53678 54516 53730
rect 54348 53676 54516 53678
rect 54460 53666 54516 53676
rect 52780 53620 52836 53630
rect 52780 53526 52836 53564
rect 53452 53620 53508 53630
rect 53452 53526 53508 53564
rect 48300 53058 48356 53452
rect 51660 53506 52388 53508
rect 51660 53454 52110 53506
rect 52162 53454 52388 53506
rect 51660 53452 52388 53454
rect 53564 53508 53620 53518
rect 53564 53506 53956 53508
rect 53564 53454 53566 53506
rect 53618 53454 53956 53506
rect 53564 53452 53956 53454
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 48300 53006 48302 53058
rect 48354 53006 48356 53058
rect 48300 52994 48356 53006
rect 48748 53060 48804 53070
rect 48412 52948 48468 52958
rect 48412 52854 48468 52892
rect 46956 52144 47012 52220
rect 47516 52276 47572 52286
rect 47516 52182 47572 52220
rect 48748 52276 48804 53004
rect 50316 53060 50372 53070
rect 50316 52966 50372 53004
rect 51660 52948 51716 53452
rect 52108 53442 52164 53452
rect 53564 53442 53620 53452
rect 52668 53172 52724 53182
rect 52668 53078 52724 53116
rect 53228 53172 53284 53182
rect 51324 52946 51716 52948
rect 51324 52894 51662 52946
rect 51714 52894 51716 52946
rect 51324 52892 51716 52894
rect 50204 52836 50260 52846
rect 50204 52742 50260 52780
rect 50764 52836 50820 52846
rect 50764 52742 50820 52780
rect 48748 52144 48804 52220
rect 49308 52276 49364 52286
rect 51324 52276 51380 52892
rect 51660 52882 51716 52892
rect 51884 53058 51940 53070
rect 51884 53006 51886 53058
rect 51938 53006 51940 53058
rect 51884 52836 51940 53006
rect 52892 52948 52948 52958
rect 52892 52854 52948 52892
rect 51884 52770 51940 52780
rect 52444 52836 52500 52846
rect 52444 52276 52500 52780
rect 52780 52834 52836 52846
rect 52780 52782 52782 52834
rect 52834 52782 52836 52834
rect 52668 52388 52724 52398
rect 52668 52294 52724 52332
rect 49308 52182 49364 52220
rect 50876 52274 51380 52276
rect 50876 52222 51326 52274
rect 51378 52222 51380 52274
rect 50876 52220 51380 52222
rect 50876 52162 50932 52220
rect 51324 52210 51380 52220
rect 52332 52274 52500 52276
rect 52332 52222 52446 52274
rect 52498 52222 52500 52274
rect 52332 52220 52500 52222
rect 50876 52110 50878 52162
rect 50930 52110 50932 52162
rect 50876 52098 50932 52110
rect 47068 52052 47124 52062
rect 47068 51958 47124 51996
rect 52220 52052 52276 52062
rect 52220 51958 52276 51996
rect 48860 51938 48916 51950
rect 48860 51886 48862 51938
rect 48914 51886 48916 51938
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 48860 51604 48916 51886
rect 48860 51538 48916 51548
rect 49196 51940 49252 51950
rect 50540 51940 50596 51950
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 4172 50642 4228 50652
rect 49196 50708 49252 51884
rect 50428 51938 50596 51940
rect 50428 51886 50542 51938
rect 50594 51886 50596 51938
rect 50428 51884 50596 51886
rect 49644 50708 49700 50718
rect 49196 50706 49700 50708
rect 49196 50654 49198 50706
rect 49250 50654 49646 50706
rect 49698 50654 49700 50706
rect 49196 50652 49700 50654
rect 50428 50708 50484 51884
rect 50540 51874 50596 51884
rect 51996 51940 52052 51950
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 51884 51604 51940 51614
rect 51996 51604 52052 51884
rect 52108 51938 52164 51950
rect 52108 51886 52110 51938
rect 52162 51886 52164 51938
rect 52108 51716 52164 51886
rect 52108 51660 52276 51716
rect 51884 51602 52052 51604
rect 51884 51550 51886 51602
rect 51938 51550 52052 51602
rect 51884 51548 52052 51550
rect 51884 51538 51940 51548
rect 52108 51492 52164 51502
rect 52108 51398 52164 51436
rect 51996 51266 52052 51278
rect 51996 51214 51998 51266
rect 52050 51214 52052 51266
rect 50428 50652 50820 50708
rect 49196 50642 49252 50652
rect 49644 50642 49700 50652
rect 50764 50594 50820 50652
rect 50764 50542 50766 50594
rect 50818 50542 50820 50594
rect 3052 50482 3108 50494
rect 3052 50430 3054 50482
rect 3106 50430 3108 50482
rect 3052 50260 3108 50430
rect 49756 50484 49812 50494
rect 49756 50390 49812 50428
rect 50652 50484 50708 50522
rect 50652 50418 50708 50428
rect 50764 50428 50820 50542
rect 51100 50596 51156 50606
rect 51660 50596 51716 50606
rect 51100 50594 51716 50596
rect 51100 50542 51102 50594
rect 51154 50542 51662 50594
rect 51714 50542 51716 50594
rect 51100 50540 51716 50542
rect 51100 50530 51156 50540
rect 51660 50530 51716 50540
rect 51772 50596 51828 50634
rect 51772 50530 51828 50540
rect 50428 50370 50484 50382
rect 50428 50318 50430 50370
rect 50482 50318 50484 50370
rect 3052 50194 3108 50204
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 46620 50036 46676 50046
rect 46620 49942 46676 49980
rect 50204 50036 50260 50046
rect 50428 50036 50484 50318
rect 50540 50372 50596 50410
rect 50764 50372 50932 50428
rect 50540 50306 50596 50316
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50204 50034 50484 50036
rect 50204 49982 50206 50034
rect 50258 49982 50484 50034
rect 50204 49980 50484 49982
rect 50204 49970 50260 49980
rect 3052 49922 3108 49934
rect 3052 49870 3054 49922
rect 3106 49870 3108 49922
rect 3052 49812 3108 49870
rect 3052 49746 3108 49756
rect 47964 49812 48020 49822
rect 2940 49634 2996 49644
rect 3500 49698 3556 49710
rect 3500 49646 3502 49698
rect 3554 49646 3556 49698
rect 3500 49588 3556 49646
rect 46508 49700 46564 49710
rect 46508 49606 46564 49644
rect 47068 49700 47124 49710
rect 47068 49606 47124 49644
rect 3500 49522 3556 49532
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 47964 49140 48020 49756
rect 49980 49810 50036 49822
rect 49980 49758 49982 49810
rect 50034 49758 50036 49810
rect 49756 49700 49812 49710
rect 49644 49644 49756 49700
rect 49196 49588 49252 49598
rect 48076 49252 48132 49262
rect 48076 49158 48132 49196
rect 3052 49028 3108 49038
rect 3052 49026 3556 49028
rect 3052 48974 3054 49026
rect 3106 48974 3556 49026
rect 47964 49008 48020 49084
rect 48524 49140 48580 49150
rect 48524 49046 48580 49084
rect 49196 49026 49252 49532
rect 3052 48972 3556 48974
rect 3052 48962 3108 48972
rect 3500 48802 3556 48972
rect 49196 48974 49198 49026
rect 49250 48974 49252 49026
rect 49196 48962 49252 48974
rect 49532 49586 49588 49598
rect 49532 49534 49534 49586
rect 49586 49534 49588 49586
rect 3500 48750 3502 48802
rect 3554 48750 3556 48802
rect 3052 48244 3108 48254
rect 3052 48150 3108 48188
rect 2268 48066 2324 48076
rect 3500 47908 3556 48750
rect 48636 48804 48692 48814
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 48524 48468 48580 48478
rect 48636 48468 48692 48748
rect 48524 48466 48692 48468
rect 48524 48414 48526 48466
rect 48578 48414 48692 48466
rect 48524 48412 48692 48414
rect 49308 48802 49364 48814
rect 49308 48750 49310 48802
rect 49362 48750 49364 48802
rect 48524 48402 48580 48412
rect 3612 48244 3668 48254
rect 3612 48132 3668 48188
rect 47292 48132 47348 48142
rect 3612 48130 3780 48132
rect 3612 48078 3614 48130
rect 3666 48078 3780 48130
rect 3612 48076 3780 48078
rect 3612 48066 3668 48076
rect 3500 47852 3668 47908
rect 2156 47618 2212 47628
rect 3052 47460 3108 47470
rect 3052 47458 3556 47460
rect 3052 47406 3054 47458
rect 3106 47406 3556 47458
rect 3052 47404 3556 47406
rect 3052 47394 3108 47404
rect 2044 46946 2100 46956
rect 2156 47346 2212 47358
rect 2156 47294 2158 47346
rect 2210 47294 2212 47346
rect 2044 46562 2100 46574
rect 2044 46510 2046 46562
rect 2098 46510 2100 46562
rect 2044 45668 2100 46510
rect 2156 46340 2212 47294
rect 3500 47234 3556 47404
rect 3500 47182 3502 47234
rect 3554 47182 3556 47234
rect 3052 46676 3108 46686
rect 3052 46582 3108 46620
rect 2156 46274 2212 46284
rect 3052 45890 3108 45902
rect 3052 45838 3054 45890
rect 3106 45838 3108 45890
rect 2044 45602 2100 45612
rect 2156 45778 2212 45790
rect 2156 45726 2158 45778
rect 2210 45726 2212 45778
rect 2044 44994 2100 45006
rect 2044 44942 2046 44994
rect 2098 44942 2100 44994
rect 2044 44324 2100 44942
rect 2156 44996 2212 45726
rect 3052 45668 3108 45838
rect 3500 45892 3556 47182
rect 3612 47236 3668 47852
rect 3612 47170 3668 47180
rect 3724 46788 3780 48076
rect 47292 48038 47348 48076
rect 47852 48130 47908 48142
rect 47852 48078 47854 48130
rect 47906 48078 47908 48130
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 47516 47348 47572 47358
rect 47516 47254 47572 47292
rect 47852 47348 47908 48078
rect 48412 48132 48468 48142
rect 48412 48038 48468 48076
rect 47852 47282 47908 47292
rect 48188 47348 48244 47358
rect 47180 47236 47236 47246
rect 47180 47142 47236 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 3724 46722 3780 46732
rect 46508 46788 46564 46798
rect 46508 46694 46564 46732
rect 47852 46788 47908 46798
rect 47852 46694 47908 46732
rect 3500 45826 3556 45836
rect 3612 46676 3668 46686
rect 3612 46562 3668 46620
rect 46844 46674 46900 46686
rect 46844 46622 46846 46674
rect 46898 46622 46900 46674
rect 3612 46510 3614 46562
rect 3666 46510 3668 46562
rect 3500 45668 3556 45678
rect 3052 45666 3556 45668
rect 3052 45614 3502 45666
rect 3554 45614 3556 45666
rect 3052 45612 3556 45614
rect 3500 45332 3556 45612
rect 3500 45266 3556 45276
rect 3612 45220 3668 46510
rect 46060 46564 46116 46574
rect 46060 46470 46116 46508
rect 46844 46564 46900 46622
rect 46844 46498 46900 46508
rect 47628 46674 47684 46686
rect 47628 46622 47630 46674
rect 47682 46622 47684 46674
rect 47628 46564 47684 46622
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 46172 45780 46228 45790
rect 46172 45686 46228 45724
rect 46844 45780 46900 45790
rect 45836 45668 45892 45678
rect 45836 45574 45892 45612
rect 46508 45668 46564 45678
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 44380 45332 44436 45342
rect 44380 45238 44436 45276
rect 46508 45330 46564 45612
rect 46508 45278 46510 45330
rect 46562 45278 46564 45330
rect 46508 45266 46564 45278
rect 3612 45154 3668 45164
rect 45276 45220 45332 45230
rect 45276 45126 45332 45164
rect 2156 44930 2212 44940
rect 3052 45106 3108 45118
rect 3052 45054 3054 45106
rect 3106 45054 3108 45106
rect 3052 44996 3108 45054
rect 43932 45108 43988 45118
rect 43932 45014 43988 45052
rect 44604 45108 44660 45118
rect 44604 45014 44660 45052
rect 45612 45108 45668 45118
rect 45612 45014 45668 45052
rect 46284 45108 46340 45118
rect 46284 45014 46340 45052
rect 3052 44930 3108 44940
rect 3612 44996 3668 45006
rect 3612 44902 3668 44940
rect 43708 44996 43764 45006
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 2044 44258 2100 44268
rect 3052 44322 3108 44334
rect 3052 44270 3054 44322
rect 3106 44270 3108 44322
rect 2156 44210 2212 44222
rect 2156 44158 2158 44210
rect 2210 44158 2212 44210
rect 2156 43652 2212 44158
rect 3052 44100 3108 44270
rect 43708 44210 43764 44940
rect 46396 44996 46452 45006
rect 46396 44322 46452 44940
rect 46396 44270 46398 44322
rect 46450 44270 46452 44322
rect 43708 44158 43710 44210
rect 43762 44158 43764 44210
rect 43708 44146 43764 44158
rect 44044 44212 44100 44222
rect 44044 44118 44100 44156
rect 44604 44212 44660 44222
rect 44604 44118 44660 44156
rect 45276 44212 45332 44222
rect 3052 44034 3108 44044
rect 3500 44100 3556 44110
rect 3500 44006 3556 44044
rect 42924 44100 42980 44110
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 42924 43762 42980 44044
rect 42924 43710 42926 43762
rect 42978 43710 42980 43762
rect 42924 43698 42980 43710
rect 44380 43764 44436 43802
rect 44380 43698 44436 43708
rect 2156 43586 2212 43596
rect 3052 43538 3108 43550
rect 3052 43486 3054 43538
rect 3106 43486 3108 43538
rect 2044 43426 2100 43438
rect 2044 43374 2046 43426
rect 2098 43374 2100 43426
rect 2044 42980 2100 43374
rect 3052 43428 3108 43486
rect 43260 43538 43316 43550
rect 43260 43486 43262 43538
rect 43314 43486 43316 43538
rect 3052 43362 3108 43372
rect 3612 43428 3668 43438
rect 3612 43334 3668 43372
rect 42252 43428 42308 43438
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 2044 42914 2100 42924
rect 3052 42754 3108 42766
rect 3052 42702 3054 42754
rect 3106 42702 3108 42754
rect 2156 42642 2212 42654
rect 2156 42590 2158 42642
rect 2210 42590 2212 42642
rect 2156 42308 2212 42590
rect 3052 42532 3108 42702
rect 41916 42756 41972 42766
rect 41916 42662 41972 42700
rect 42252 42644 42308 43372
rect 42476 43428 42532 43438
rect 42476 43334 42532 43372
rect 43260 43428 43316 43486
rect 44156 43540 44212 43550
rect 44156 43538 44324 43540
rect 44156 43486 44158 43538
rect 44210 43486 44324 43538
rect 44156 43484 44324 43486
rect 44156 43474 44212 43484
rect 43260 43362 43316 43372
rect 44268 43428 44324 43484
rect 42588 42756 42644 42766
rect 42588 42662 42644 42700
rect 43372 42756 43428 42766
rect 43372 42662 43428 42700
rect 42364 42644 42420 42654
rect 42252 42642 42420 42644
rect 42252 42590 42366 42642
rect 42418 42590 42420 42642
rect 42252 42588 42420 42590
rect 42364 42578 42420 42588
rect 44044 42644 44100 42654
rect 3052 42466 3108 42476
rect 3500 42532 3556 42542
rect 3500 42438 3556 42476
rect 41692 42532 41748 42542
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 2156 42242 2212 42252
rect 41692 42194 41748 42476
rect 43708 42532 43764 42542
rect 43708 42438 43764 42476
rect 44044 42532 44100 42588
rect 44156 42532 44212 42542
rect 44044 42530 44212 42532
rect 44044 42478 44158 42530
rect 44210 42478 44212 42530
rect 44044 42476 44212 42478
rect 41692 42142 41694 42194
rect 41746 42142 41748 42194
rect 41692 42130 41748 42142
rect 43036 42082 43092 42094
rect 43036 42030 43038 42082
rect 43090 42030 43092 42082
rect 3052 41970 3108 41982
rect 3052 41918 3054 41970
rect 3106 41918 3108 41970
rect 2044 41858 2100 41870
rect 2044 41806 2046 41858
rect 2098 41806 2100 41858
rect 2044 41636 2100 41806
rect 3052 41860 3108 41918
rect 42028 41970 42084 41982
rect 42028 41918 42030 41970
rect 42082 41918 42084 41970
rect 3052 41794 3108 41804
rect 3612 41860 3668 41870
rect 3612 41766 3668 41804
rect 41020 41860 41076 41870
rect 2044 41570 2100 41580
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 3052 41186 3108 41198
rect 3052 41134 3054 41186
rect 3106 41134 3108 41186
rect 2156 41074 2212 41086
rect 2156 41022 2158 41074
rect 2210 41022 2212 41074
rect 2156 40964 2212 41022
rect 2156 40898 2212 40908
rect 3052 40964 3108 41134
rect 41020 41074 41076 41804
rect 42028 41860 42084 41918
rect 42812 41972 42868 41982
rect 42812 41970 42980 41972
rect 42812 41918 42814 41970
rect 42866 41918 42980 41970
rect 42812 41916 42980 41918
rect 42812 41906 42868 41916
rect 42028 41794 42084 41804
rect 42924 41860 42980 41916
rect 42140 41186 42196 41198
rect 42140 41134 42142 41186
rect 42194 41134 42196 41186
rect 41020 41022 41022 41074
rect 41074 41022 41076 41074
rect 41020 41010 41076 41022
rect 41356 41074 41412 41086
rect 41356 41022 41358 41074
rect 41410 41022 41412 41074
rect 3052 40898 3108 40908
rect 3500 40964 3556 40974
rect 40012 40964 40068 40974
rect 3500 40870 3556 40908
rect 39900 40962 40068 40964
rect 39900 40910 40014 40962
rect 40066 40910 40068 40962
rect 39900 40908 40068 40910
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 39340 40514 39396 40526
rect 39340 40462 39342 40514
rect 39394 40462 39396 40514
rect 3052 40404 3108 40414
rect 3052 40310 3108 40348
rect 3612 40404 3668 40414
rect 3612 40310 3668 40348
rect 39340 40404 39396 40462
rect 39340 40338 39396 40348
rect 39676 40404 39732 40414
rect 39900 40404 39956 40908
rect 40012 40898 40068 40908
rect 40236 40964 40292 40974
rect 40236 40626 40292 40908
rect 40572 40964 40628 40974
rect 40572 40870 40628 40908
rect 41356 40964 41412 41022
rect 41356 40898 41412 40908
rect 42140 40964 42196 41134
rect 42364 41076 42420 41086
rect 42364 40982 42420 41020
rect 40236 40574 40238 40626
rect 40290 40574 40292 40626
rect 40236 40562 40292 40574
rect 41916 40516 41972 40526
rect 41916 40422 41972 40460
rect 39676 40402 39956 40404
rect 39676 40350 39678 40402
rect 39730 40350 39956 40402
rect 39676 40348 39956 40350
rect 39676 40338 39732 40348
rect 2044 40292 2100 40302
rect 2044 40198 2100 40236
rect 38892 40290 38948 40302
rect 38892 40238 38894 40290
rect 38946 40238 38948 40290
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 2156 39620 2212 39630
rect 2156 39526 2212 39564
rect 3052 39618 3108 39630
rect 3052 39566 3054 39618
rect 3106 39566 3108 39618
rect 3052 39508 3108 39566
rect 3052 39442 3108 39452
rect 3612 39508 3668 39518
rect 3612 39414 3668 39452
rect 38780 39508 38836 39518
rect 38780 39414 38836 39452
rect 38332 39396 38388 39406
rect 38332 39302 38388 39340
rect 38892 39396 38948 40238
rect 38892 39330 38948 39340
rect 39116 39508 39172 39518
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 2156 38948 2212 38958
rect 2156 38854 2212 38892
rect 38332 38946 38388 38958
rect 38332 38894 38334 38946
rect 38386 38894 38388 38946
rect 3052 38836 3108 38846
rect 3052 38742 3108 38780
rect 3612 38836 3668 38846
rect 3612 38742 3668 38780
rect 38332 38836 38388 38894
rect 38332 38770 38388 38780
rect 38668 38836 38724 38846
rect 38668 38742 38724 38780
rect 37884 38724 37940 38734
rect 37884 38630 37940 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 2044 38276 2100 38286
rect 2044 38162 2100 38220
rect 2044 38110 2046 38162
rect 2098 38110 2100 38162
rect 2044 38098 2100 38110
rect 3052 38050 3108 38062
rect 3052 37998 3054 38050
rect 3106 37998 3108 38050
rect 3052 37828 3108 37998
rect 37996 37940 38052 37950
rect 37996 37846 38052 37884
rect 38668 37940 38724 37950
rect 3052 37762 3108 37772
rect 3612 37828 3668 37838
rect 3612 37734 3668 37772
rect 37660 37828 37716 37838
rect 37660 37734 37716 37772
rect 19836 37660 20100 37670
rect 2156 37604 2212 37614
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 2156 37378 2212 37548
rect 2156 37326 2158 37378
rect 2210 37326 2212 37378
rect 2156 37314 2212 37326
rect 36988 37378 37044 37390
rect 36988 37326 36990 37378
rect 37042 37326 37044 37378
rect 3052 37266 3108 37278
rect 3052 37214 3054 37266
rect 3106 37214 3108 37266
rect 3052 37044 3108 37214
rect 3052 36978 3108 36988
rect 3612 37154 3668 37166
rect 3612 37102 3614 37154
rect 3666 37102 3668 37154
rect 3612 37044 3668 37102
rect 36540 37156 36596 37166
rect 36540 37062 36596 37100
rect 3612 36978 3668 36988
rect 36988 37044 37044 37326
rect 38332 37380 38388 37390
rect 38332 37286 38388 37324
rect 36988 36978 37044 36988
rect 37212 37266 37268 37278
rect 37212 37214 37214 37266
rect 37266 37214 37268 37266
rect 37212 37156 37268 37214
rect 2044 36932 2100 36942
rect 2044 36594 2100 36876
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 2044 36542 2046 36594
rect 2098 36542 2100 36594
rect 2044 36530 2100 36542
rect 3052 36482 3108 36494
rect 3052 36430 3054 36482
rect 3106 36430 3108 36482
rect 2156 36260 2212 36270
rect 2156 35810 2212 36204
rect 3052 36260 3108 36430
rect 35868 36372 35924 36382
rect 35868 36278 35924 36316
rect 36652 36372 36708 36382
rect 36652 36278 36708 36316
rect 3052 36194 3108 36204
rect 3612 36260 3668 36270
rect 3612 36166 3668 36204
rect 35308 36258 35364 36270
rect 35308 36206 35310 36258
rect 35362 36206 35364 36258
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 2156 35758 2158 35810
rect 2210 35758 2212 35810
rect 2156 35746 2212 35758
rect 3052 35812 3108 35822
rect 3052 35698 3108 35756
rect 3052 35646 3054 35698
rect 3106 35646 3108 35698
rect 3052 35634 3108 35646
rect 3612 35812 3668 35822
rect 2044 35588 2100 35598
rect 2044 35026 2100 35532
rect 2044 34974 2046 35026
rect 2098 34974 2100 35026
rect 2044 34962 2100 34974
rect 3612 35026 3668 35756
rect 34636 35810 34692 35822
rect 34636 35758 34638 35810
rect 34690 35758 34692 35810
rect 4844 35698 4900 35710
rect 4844 35646 4846 35698
rect 4898 35646 4900 35698
rect 3612 34974 3614 35026
rect 3666 34974 3668 35026
rect 3612 34962 3668 34974
rect 3836 35586 3892 35598
rect 3836 35534 3838 35586
rect 3890 35534 3892 35586
rect 3052 34914 3108 34926
rect 3052 34862 3054 34914
rect 3106 34862 3108 34914
rect 3052 34692 3108 34862
rect 3836 34916 3892 35534
rect 4844 35588 4900 35646
rect 4844 35522 4900 35532
rect 5404 35588 5460 35598
rect 5404 35494 5460 35532
rect 34188 35588 34244 35598
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 3836 34850 3892 34860
rect 33740 34916 33796 34926
rect 33740 34822 33796 34860
rect 34188 34802 34244 35532
rect 34524 34916 34580 34926
rect 34524 34822 34580 34860
rect 34188 34750 34190 34802
rect 34242 34750 34244 34802
rect 34188 34738 34244 34750
rect 3052 34626 3108 34636
rect 4060 34692 4116 34702
rect 4060 34598 4116 34636
rect 34636 34692 34692 35758
rect 34972 35700 35028 35710
rect 34972 35606 35028 35644
rect 35308 35700 35364 36206
rect 36316 36260 36372 36270
rect 36316 36166 36372 36204
rect 35532 35812 35588 35822
rect 35532 35718 35588 35756
rect 35868 35812 35924 35822
rect 35868 35718 35924 35756
rect 36764 35812 36820 35822
rect 35308 35634 35364 35644
rect 36092 35700 36148 35710
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 34916 35252 34926
rect 35252 34860 35588 34916
rect 35196 34784 35252 34860
rect 34636 34626 34692 34636
rect 35420 34692 35476 34702
rect 35420 34598 35476 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 2156 34244 2212 34254
rect 2156 34150 2212 34188
rect 33628 34242 33684 34254
rect 33628 34190 33630 34242
rect 33682 34190 33684 34242
rect 3052 34130 3108 34142
rect 3052 34078 3054 34130
rect 3106 34078 3108 34130
rect 3052 33908 3108 34078
rect 32956 34132 33012 34142
rect 32956 34038 33012 34076
rect 3052 33842 3108 33852
rect 3612 34018 3668 34030
rect 3612 33966 3614 34018
rect 3666 33966 3668 34018
rect 3612 33908 3668 33966
rect 3612 33842 3668 33852
rect 33628 33908 33684 34190
rect 35084 34244 35140 34254
rect 35084 34150 35140 34188
rect 33964 34132 34020 34142
rect 33964 34038 34020 34076
rect 34860 34132 34916 34142
rect 33628 33842 33684 33852
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 2044 33572 2100 33582
rect 2044 33458 2100 33516
rect 2044 33406 2046 33458
rect 2098 33406 2100 33458
rect 2044 33394 2100 33406
rect 3052 33346 3108 33358
rect 3052 33294 3054 33346
rect 3106 33294 3108 33346
rect 3052 33124 3108 33294
rect 32508 33348 32564 33358
rect 32508 33254 32564 33292
rect 33180 33348 33236 33358
rect 3052 33058 3108 33068
rect 3612 33124 3668 33134
rect 3612 33030 3668 33068
rect 32956 33124 33012 33134
rect 32956 33030 33012 33068
rect 19836 32956 20100 32966
rect 2156 32900 2212 32910
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 2156 32674 2212 32844
rect 2156 32622 2158 32674
rect 2210 32622 2212 32674
rect 2156 32610 2212 32622
rect 32172 32674 32228 32686
rect 32172 32622 32174 32674
rect 32226 32622 32228 32674
rect 3052 32562 3108 32574
rect 3052 32510 3054 32562
rect 3106 32510 3108 32562
rect 3052 32340 3108 32510
rect 3052 32274 3108 32284
rect 3612 32450 3668 32462
rect 3612 32398 3614 32450
rect 3666 32398 3668 32450
rect 3612 32340 3668 32398
rect 31724 32452 31780 32462
rect 31724 32358 31780 32396
rect 3612 32274 3668 32284
rect 32172 32340 32228 32622
rect 32172 32274 32228 32284
rect 32508 32564 32564 32574
rect 2044 32228 2100 32238
rect 2044 31890 2100 32172
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 32508 31948 32564 32508
rect 2044 31838 2046 31890
rect 2098 31838 2100 31890
rect 2044 31826 2100 31838
rect 32172 31892 32564 31948
rect 33180 31948 33236 33292
rect 34076 33348 34132 33358
rect 34132 33292 34356 33348
rect 34076 33254 34132 33292
rect 34300 32788 34356 33292
rect 34412 33124 34468 33134
rect 34412 33030 34468 33068
rect 34860 33122 34916 34076
rect 35532 34020 35588 34860
rect 36092 34914 36148 35644
rect 36092 34862 36094 34914
rect 36146 34862 36148 34914
rect 35644 34020 35700 34030
rect 35532 34018 35700 34020
rect 35532 33966 35646 34018
rect 35698 33966 35700 34018
rect 35532 33964 35700 33966
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34860 33070 34862 33122
rect 34914 33070 34916 33122
rect 34412 32788 34468 32798
rect 34300 32786 34468 32788
rect 34300 32734 34414 32786
rect 34466 32734 34468 32786
rect 34300 32732 34468 32734
rect 34412 32722 34468 32732
rect 33964 32676 34020 32686
rect 33964 32582 34020 32620
rect 33404 32564 33460 32574
rect 33180 31892 33348 31948
rect 3052 31778 3108 31790
rect 3052 31726 3054 31778
rect 3106 31726 3108 31778
rect 2156 31556 2212 31566
rect 2156 31106 2212 31500
rect 3052 31556 3108 31726
rect 31164 31668 31220 31678
rect 31164 31574 31220 31612
rect 31948 31668 32004 31678
rect 31948 31574 32004 31612
rect 3052 31490 3108 31500
rect 3612 31556 3668 31566
rect 3612 31462 3668 31500
rect 30716 31554 30772 31566
rect 30716 31502 30718 31554
rect 30770 31502 30772 31554
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 2156 31054 2158 31106
rect 2210 31054 2212 31106
rect 2156 31042 2212 31054
rect 3052 31108 3108 31118
rect 3052 30994 3108 31052
rect 3052 30942 3054 30994
rect 3106 30942 3108 30994
rect 3052 30930 3108 30942
rect 3612 31108 3668 31118
rect 2156 30884 2212 30894
rect 2156 30210 2212 30828
rect 2156 30158 2158 30210
rect 2210 30158 2212 30210
rect 2156 30146 2212 30158
rect 3052 30210 3108 30222
rect 3052 30158 3054 30210
rect 3106 30158 3108 30210
rect 3052 29988 3108 30158
rect 3612 30210 3668 31052
rect 30044 31106 30100 31118
rect 30044 31054 30046 31106
rect 30098 31054 30100 31106
rect 4844 30994 4900 31006
rect 4844 30942 4846 30994
rect 4898 30942 4900 30994
rect 3612 30158 3614 30210
rect 3666 30158 3668 30210
rect 3612 30146 3668 30158
rect 3836 30882 3892 30894
rect 3836 30830 3838 30882
rect 3890 30830 3892 30882
rect 3836 30212 3892 30830
rect 4844 30884 4900 30942
rect 4844 30818 4900 30828
rect 5404 30884 5460 30894
rect 5404 30790 5460 30828
rect 29596 30884 29652 30894
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 3836 30146 3892 30156
rect 3052 29922 3108 29932
rect 4060 29988 4116 29998
rect 4060 29894 4116 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 29596 29650 29652 30828
rect 29596 29598 29598 29650
rect 29650 29598 29652 29650
rect 29596 29586 29652 29598
rect 29932 29986 29988 29998
rect 29932 29934 29934 29986
rect 29986 29934 29988 29986
rect 2156 29540 2212 29550
rect 2156 29446 2212 29484
rect 28700 29538 28756 29550
rect 28700 29486 28702 29538
rect 28754 29486 28756 29538
rect 3052 29426 3108 29438
rect 3052 29374 3054 29426
rect 3106 29374 3108 29426
rect 3052 29204 3108 29374
rect 3052 29138 3108 29148
rect 3612 29314 3668 29326
rect 3612 29262 3614 29314
rect 3666 29262 3668 29314
rect 3612 29204 3668 29262
rect 28252 29316 28308 29326
rect 28252 29222 28308 29260
rect 3612 29138 3668 29148
rect 28700 29204 28756 29486
rect 28700 29138 28756 29148
rect 29036 29426 29092 29438
rect 29036 29374 29038 29426
rect 29090 29374 29092 29426
rect 29036 29316 29092 29374
rect 29932 29428 29988 29934
rect 30044 29988 30100 31054
rect 30044 29922 30100 29932
rect 30268 30996 30324 31006
rect 30716 30996 30772 31502
rect 31612 31556 31668 31566
rect 31612 31462 31668 31500
rect 30940 31108 30996 31118
rect 30940 31014 30996 31052
rect 30268 30994 30772 30996
rect 30268 30942 30270 30994
rect 30322 30942 30772 30994
rect 30268 30940 30772 30942
rect 31276 30996 31332 31006
rect 29932 29334 29988 29372
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 2044 28868 2100 28878
rect 2044 28754 2100 28812
rect 2044 28702 2046 28754
rect 2098 28702 2100 28754
rect 2044 28690 2100 28702
rect 3052 28644 3108 28654
rect 3052 28550 3108 28588
rect 3612 28644 3668 28654
rect 3612 28550 3668 28588
rect 27804 28642 27860 28654
rect 27804 28590 27806 28642
rect 27858 28590 27860 28642
rect 27804 28532 27860 28590
rect 27804 28466 27860 28476
rect 28252 28644 28308 28654
rect 28252 28530 28308 28588
rect 29036 28644 29092 29260
rect 30268 28866 30324 30940
rect 31276 30902 31332 30940
rect 32060 30996 32116 31006
rect 32060 30322 32116 30940
rect 32060 30270 32062 30322
rect 32114 30270 32116 30322
rect 30380 30098 30436 30110
rect 30380 30046 30382 30098
rect 30434 30046 30436 30098
rect 30380 29428 30436 30046
rect 31276 30098 31332 30110
rect 31276 30046 31278 30098
rect 31330 30046 31332 30098
rect 30716 29988 30772 29998
rect 30716 29894 30772 29932
rect 30828 29540 30884 29550
rect 30828 29446 30884 29484
rect 30380 29362 30436 29372
rect 30492 29426 30548 29438
rect 30492 29374 30494 29426
rect 30546 29374 30548 29426
rect 30268 28814 30270 28866
rect 30322 28814 30324 28866
rect 29036 28578 29092 28588
rect 29708 28644 29764 28654
rect 28252 28478 28254 28530
rect 28306 28478 28308 28530
rect 28252 28466 28308 28478
rect 28588 28532 28644 28542
rect 28588 28438 28644 28476
rect 29372 28532 29428 28542
rect 29596 28532 29652 28542
rect 29428 28530 29652 28532
rect 29428 28478 29598 28530
rect 29650 28478 29652 28530
rect 29428 28476 29652 28478
rect 19836 28252 20100 28262
rect 2156 28196 2212 28206
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 2156 27970 2212 28140
rect 2156 27918 2158 27970
rect 2210 27918 2212 27970
rect 2156 27906 2212 27918
rect 27580 27970 27636 27982
rect 27580 27918 27582 27970
rect 27634 27918 27636 27970
rect 3052 27858 3108 27870
rect 3052 27806 3054 27858
rect 3106 27806 3108 27858
rect 3052 27748 3108 27806
rect 27132 27860 27188 27870
rect 27132 27766 27188 27804
rect 3052 27682 3108 27692
rect 3612 27748 3668 27758
rect 3612 27654 3668 27692
rect 27580 27748 27636 27918
rect 28924 27972 28980 27982
rect 28924 27878 28980 27916
rect 27916 27860 27972 27870
rect 27916 27766 27972 27804
rect 28476 27860 28532 27870
rect 28588 27860 28644 27870
rect 28532 27858 28644 27860
rect 28532 27806 28590 27858
rect 28642 27806 28644 27858
rect 28532 27804 28644 27806
rect 27580 27682 27636 27692
rect 2044 27524 2100 27534
rect 2044 27186 2100 27468
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 2044 27134 2046 27186
rect 2098 27134 2100 27186
rect 2044 27122 2100 27134
rect 3052 27076 3108 27086
rect 3052 26982 3108 27020
rect 3612 27076 3668 27086
rect 3612 26982 3668 27020
rect 26908 27076 26964 27086
rect 26460 26964 26516 26974
rect 26460 26870 26516 26908
rect 2156 26852 2212 26862
rect 2156 26402 2212 26796
rect 26908 26850 26964 27020
rect 26908 26798 26910 26850
rect 26962 26798 26964 26850
rect 26908 26786 26964 26798
rect 27244 26964 27300 26974
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 2156 26350 2158 26402
rect 2210 26350 2212 26402
rect 2156 26338 2212 26350
rect 26236 26402 26292 26414
rect 26236 26350 26238 26402
rect 26290 26350 26292 26402
rect 2940 26290 2996 26302
rect 2940 26238 2942 26290
rect 2994 26238 2996 26290
rect 2044 26180 2100 26190
rect 2044 25618 2100 26124
rect 2044 25566 2046 25618
rect 2098 25566 2100 25618
rect 2044 25554 2100 25566
rect 2940 25284 2996 26238
rect 4844 26290 4900 26302
rect 4844 26238 4846 26290
rect 4898 26238 4900 26290
rect 3836 26178 3892 26190
rect 3836 26126 3838 26178
rect 3890 26126 3892 26178
rect 3052 25506 3108 25518
rect 3052 25454 3054 25506
rect 3106 25454 3108 25506
rect 3052 25396 3108 25454
rect 3836 25508 3892 26126
rect 4844 26180 4900 26238
rect 4844 26114 4900 26124
rect 5404 26180 5460 26190
rect 5404 26086 5460 26124
rect 24332 26180 24388 26190
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 3836 25442 3892 25452
rect 3052 25330 3108 25340
rect 4060 25396 4116 25406
rect 4060 25302 4116 25340
rect 24332 25394 24388 26124
rect 25788 26180 25844 26190
rect 25788 26086 25844 26124
rect 25564 25508 25620 25518
rect 25564 25414 25620 25452
rect 24332 25342 24334 25394
rect 24386 25342 24388 25394
rect 24332 25330 24388 25342
rect 24668 25396 24724 25406
rect 25228 25396 25284 25406
rect 24668 25394 24836 25396
rect 24668 25342 24670 25394
rect 24722 25342 24836 25394
rect 24668 25340 24836 25342
rect 24668 25330 24724 25340
rect 2940 25218 2996 25228
rect 3612 25284 3668 25294
rect 3612 25190 3668 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 2156 24836 2212 24846
rect 2156 24742 2212 24780
rect 24108 24834 24164 24846
rect 24108 24782 24110 24834
rect 24162 24782 24164 24834
rect 3052 24722 3108 24734
rect 3052 24670 3054 24722
rect 3106 24670 3108 24722
rect 3052 24612 3108 24670
rect 3052 24546 3108 24556
rect 3612 24612 3668 24622
rect 3612 24518 3668 24556
rect 24108 24612 24164 24782
rect 24108 24546 24164 24556
rect 24444 24722 24500 24734
rect 24444 24670 24446 24722
rect 24498 24670 24500 24722
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 2044 24164 2100 24174
rect 2044 24050 2100 24108
rect 2044 23998 2046 24050
rect 2098 23998 2100 24050
rect 2044 23986 2100 23998
rect 3052 23938 3108 23950
rect 3052 23886 3054 23938
rect 3106 23886 3108 23938
rect 3052 23716 3108 23886
rect 23996 23826 24052 23838
rect 23996 23774 23998 23826
rect 24050 23774 24052 23826
rect 3052 23650 3108 23660
rect 3612 23716 3668 23726
rect 3612 23622 3668 23660
rect 23100 23714 23156 23726
rect 23100 23662 23102 23714
rect 23154 23662 23156 23714
rect 19836 23548 20100 23558
rect 2156 23492 2212 23502
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 2156 23266 2212 23436
rect 2156 23214 2158 23266
rect 2210 23214 2212 23266
rect 2156 23202 2212 23214
rect 22428 23266 22484 23278
rect 22428 23214 22430 23266
rect 22482 23214 22484 23266
rect 3052 23154 3108 23166
rect 3052 23102 3054 23154
rect 3106 23102 3108 23154
rect 3052 23044 3108 23102
rect 3052 22978 3108 22988
rect 3612 23044 3668 23054
rect 3612 22950 3668 22988
rect 22428 23044 22484 23214
rect 22764 23156 22820 23166
rect 22764 23062 22820 23100
rect 23100 23156 23156 23662
rect 23660 23716 23716 23726
rect 23660 23622 23716 23660
rect 23996 23604 24052 23774
rect 24444 23716 24500 24670
rect 24780 24612 24836 25340
rect 25228 25302 25284 25340
rect 26236 25284 26292 26350
rect 26460 26290 26516 26302
rect 26460 26238 26462 26290
rect 26514 26238 26516 26290
rect 26460 26180 26516 26238
rect 26236 25218 26292 25228
rect 26348 25508 26404 25518
rect 26348 25394 26404 25452
rect 26348 25342 26350 25394
rect 26402 25342 26404 25394
rect 26124 24836 26180 24846
rect 26124 24742 26180 24780
rect 25900 24722 25956 24734
rect 25900 24670 25902 24722
rect 25954 24670 25956 24722
rect 24892 24612 24948 24622
rect 24780 24556 24892 24612
rect 24892 24518 24948 24556
rect 25900 24612 25956 24670
rect 25564 23938 25620 23950
rect 25564 23886 25566 23938
rect 25618 23886 25620 23938
rect 24668 23716 24724 23726
rect 24444 23660 24668 23716
rect 24668 23622 24724 23660
rect 25564 23716 25620 23886
rect 23884 23268 23940 23278
rect 23884 23174 23940 23212
rect 23100 23090 23156 23100
rect 23660 23156 23716 23166
rect 23716 23100 23828 23156
rect 23660 23024 23716 23100
rect 22428 22978 22484 22988
rect 2044 22820 2100 22830
rect 2044 22482 2100 22764
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 2044 22430 2046 22482
rect 2098 22430 2100 22482
rect 2044 22418 2100 22430
rect 3052 22370 3108 22382
rect 3052 22318 3054 22370
rect 3106 22318 3108 22370
rect 3052 22260 3108 22318
rect 3052 22194 3108 22204
rect 3612 22260 3668 22270
rect 3612 22166 3668 22204
rect 22092 22260 22148 22270
rect 22092 22166 22148 22204
rect 22428 22260 22484 22270
rect 2156 22148 2212 22158
rect 2156 21698 2212 22092
rect 21644 22148 21700 22158
rect 21644 22054 21700 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 21644 21700 21700 21710
rect 2156 21646 2158 21698
rect 2210 21646 2212 21698
rect 2156 21634 2212 21646
rect 21532 21698 21700 21700
rect 21532 21646 21646 21698
rect 21698 21646 21700 21698
rect 21532 21644 21700 21646
rect 2940 21586 2996 21598
rect 2940 21534 2942 21586
rect 2994 21534 2996 21586
rect 2044 21476 2100 21486
rect 2044 20914 2100 21420
rect 2044 20862 2046 20914
rect 2098 20862 2100 20914
rect 2044 20850 2100 20862
rect 2940 20580 2996 21534
rect 4844 21586 4900 21598
rect 4844 21534 4846 21586
rect 4898 21534 4900 21586
rect 3836 21474 3892 21486
rect 3836 21422 3838 21474
rect 3890 21422 3892 21474
rect 3052 20802 3108 20814
rect 3052 20750 3054 20802
rect 3106 20750 3108 20802
rect 3052 20692 3108 20750
rect 3836 20804 3892 21422
rect 4844 21476 4900 21534
rect 4844 21410 4900 21420
rect 5404 21476 5460 21486
rect 5404 21382 5460 21420
rect 19628 21476 19684 21486
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 3836 20738 3892 20748
rect 3052 20626 3108 20636
rect 4060 20692 4116 20702
rect 4060 20598 4116 20636
rect 2940 20514 2996 20524
rect 3612 20580 3668 20590
rect 3612 20486 3668 20524
rect 19628 20244 19684 21420
rect 20636 20578 20692 20590
rect 20636 20526 20638 20578
rect 20690 20526 20692 20578
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19964 20244 20020 20254
rect 19628 20242 20020 20244
rect 19628 20190 19966 20242
rect 20018 20190 20020 20242
rect 19628 20188 20020 20190
rect 19964 20178 20020 20188
rect 2156 20132 2212 20142
rect 2156 20038 2212 20076
rect 3052 20018 3108 20030
rect 3052 19966 3054 20018
rect 3106 19966 3108 20018
rect 3052 19908 3108 19966
rect 19516 20020 19572 20030
rect 19516 19926 19572 19964
rect 20300 20020 20356 20030
rect 3052 19842 3108 19852
rect 3612 19908 3668 19918
rect 3612 19814 3668 19852
rect 19404 19908 19460 19918
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 2044 19460 2100 19470
rect 2044 19346 2100 19404
rect 2044 19294 2046 19346
rect 2098 19294 2100 19346
rect 2044 19282 2100 19294
rect 3052 19234 3108 19246
rect 3052 19182 3054 19234
rect 3106 19182 3108 19234
rect 3052 18900 3108 19182
rect 18956 19122 19012 19134
rect 18956 19070 18958 19122
rect 19010 19070 19012 19122
rect 3052 18834 3108 18844
rect 3612 19010 3668 19022
rect 3612 18958 3614 19010
rect 3666 18958 3668 19010
rect 3612 18900 3668 18958
rect 3612 18834 3668 18844
rect 18172 19010 18228 19022
rect 18172 18958 18174 19010
rect 18226 18958 18228 19010
rect 2156 18788 2212 18798
rect 2156 18562 2212 18732
rect 18172 18676 18228 18958
rect 18620 19010 18676 19022
rect 18620 18958 18622 19010
rect 18674 18958 18676 19010
rect 18620 18900 18676 18958
rect 18620 18834 18676 18844
rect 18172 18610 18228 18620
rect 18956 18676 19012 19070
rect 19404 19124 19460 19852
rect 19516 19124 19572 19134
rect 19404 19122 19572 19124
rect 19404 19070 19518 19122
rect 19570 19070 19572 19122
rect 19404 19068 19572 19070
rect 19516 19058 19572 19068
rect 19852 19124 19908 19134
rect 19852 19030 19908 19068
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 18956 18610 19012 18620
rect 2156 18510 2158 18562
rect 2210 18510 2212 18562
rect 2156 18498 2212 18510
rect 18620 18562 18676 18574
rect 18620 18510 18622 18562
rect 18674 18510 18676 18562
rect 3052 18450 3108 18462
rect 3052 18398 3054 18450
rect 3106 18398 3108 18450
rect 3052 18340 3108 18398
rect 3052 18274 3108 18284
rect 3612 18340 3668 18350
rect 3612 18246 3668 18284
rect 18172 18338 18228 18350
rect 18172 18286 18174 18338
rect 18226 18286 18228 18338
rect 2044 18116 2100 18126
rect 2044 17778 2100 18060
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 2044 17726 2046 17778
rect 2098 17726 2100 17778
rect 2044 17714 2100 17726
rect 3052 17666 3108 17678
rect 3052 17614 3054 17666
rect 3106 17614 3108 17666
rect 2156 17444 2212 17454
rect 2156 16994 2212 17388
rect 3052 17444 3108 17614
rect 18060 17556 18116 17566
rect 18172 17556 18228 18286
rect 18620 18340 18676 18510
rect 20076 18564 20132 18574
rect 18956 18452 19012 18462
rect 18956 18450 19124 18452
rect 18956 18398 18958 18450
rect 19010 18398 19124 18450
rect 18956 18396 19124 18398
rect 18956 18386 19012 18396
rect 18620 18274 18676 18284
rect 18956 17892 19012 17902
rect 18620 17556 18676 17566
rect 18060 17554 18228 17556
rect 18060 17502 18062 17554
rect 18114 17502 18228 17554
rect 18060 17500 18228 17502
rect 18508 17554 18676 17556
rect 18508 17502 18622 17554
rect 18674 17502 18676 17554
rect 18508 17500 18676 17502
rect 3052 17378 3108 17388
rect 3612 17444 3668 17454
rect 3612 17350 3668 17388
rect 16380 17442 16436 17454
rect 17164 17444 17220 17454
rect 16380 17390 16382 17442
rect 16434 17390 16436 17442
rect 2156 16942 2158 16994
rect 2210 16942 2212 16994
rect 2156 16930 2212 16942
rect 3052 16996 3108 17006
rect 3052 16882 3108 16940
rect 3052 16830 3054 16882
rect 3106 16830 3108 16882
rect 3052 16818 3108 16830
rect 3612 16996 3668 17006
rect 2044 16772 2100 16782
rect 2044 16210 2100 16716
rect 2044 16158 2046 16210
rect 2098 16158 2100 16210
rect 2044 16146 2100 16158
rect 3612 16210 3668 16940
rect 15708 16996 15764 17006
rect 15708 16994 15876 16996
rect 15708 16942 15710 16994
rect 15762 16942 15876 16994
rect 15708 16940 15876 16942
rect 15708 16930 15764 16940
rect 4844 16884 4900 16894
rect 4844 16790 4900 16828
rect 5404 16884 5460 16894
rect 5404 16790 5460 16828
rect 15596 16884 15652 16894
rect 3612 16158 3614 16210
rect 3666 16158 3668 16210
rect 3612 16146 3668 16158
rect 3836 16770 3892 16782
rect 3836 16718 3838 16770
rect 3890 16718 3892 16770
rect 3052 16098 3108 16110
rect 3052 16046 3054 16098
rect 3106 16046 3108 16098
rect 3052 15876 3108 16046
rect 3836 16100 3892 16718
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 3836 16034 3892 16044
rect 15596 15988 15652 16828
rect 15708 15988 15764 15998
rect 15596 15986 15764 15988
rect 15596 15934 15710 15986
rect 15762 15934 15764 15986
rect 15596 15932 15764 15934
rect 15708 15922 15764 15932
rect 3052 15810 3108 15820
rect 4060 15876 4116 15886
rect 4060 15782 4116 15820
rect 15820 15876 15876 16940
rect 15820 15810 15876 15820
rect 15932 16884 15988 16894
rect 16380 16884 16436 17390
rect 17052 17442 17220 17444
rect 17052 17390 17166 17442
rect 17218 17390 17220 17442
rect 17052 17388 17220 17390
rect 16604 16996 16660 17006
rect 16604 16902 16660 16940
rect 15932 16882 16436 16884
rect 15932 16830 15934 16882
rect 15986 16830 16436 16882
rect 15932 16828 16436 16830
rect 16940 16882 16996 16894
rect 16940 16830 16942 16882
rect 16994 16830 16996 16882
rect 2156 15428 2212 15438
rect 2156 15334 2212 15372
rect 14700 15426 14756 15438
rect 14700 15374 14702 15426
rect 14754 15374 14756 15426
rect 3052 15314 3108 15326
rect 3052 15262 3054 15314
rect 3106 15262 3108 15314
rect 3052 15204 3108 15262
rect 3052 15138 3108 15148
rect 3612 15204 3668 15214
rect 3612 15110 3668 15148
rect 14700 15204 14756 15374
rect 15036 15314 15092 15326
rect 15036 15262 15038 15314
rect 15090 15262 15092 15314
rect 15036 15204 15092 15262
rect 15484 15316 15540 15326
rect 15484 15204 15540 15260
rect 15036 15202 15540 15204
rect 15036 15150 15486 15202
rect 15538 15150 15540 15202
rect 15036 15148 15540 15150
rect 15932 15204 15988 16828
rect 16940 16322 16996 16830
rect 16940 16270 16942 16322
rect 16994 16270 16996 16322
rect 16828 16212 16884 16222
rect 16940 16212 16996 16270
rect 16828 16210 16996 16212
rect 16828 16158 16830 16210
rect 16882 16158 16996 16210
rect 16828 16156 16996 16158
rect 17052 16884 17108 17388
rect 17164 17378 17220 17388
rect 17724 17444 17780 17454
rect 17724 17350 17780 17388
rect 16828 16146 16884 16156
rect 16044 15986 16100 15998
rect 16044 15934 16046 15986
rect 16098 15934 16100 15986
rect 16044 15876 16100 15934
rect 16044 15204 16100 15820
rect 16268 15204 16324 15214
rect 16044 15202 16324 15204
rect 16044 15150 16270 15202
rect 16322 15150 16324 15202
rect 16044 15148 16324 15150
rect 14700 15138 14756 15148
rect 15484 15092 15876 15148
rect 15932 15138 15988 15148
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 2044 14756 2100 14766
rect 2044 14642 2100 14700
rect 2044 14590 2046 14642
rect 2098 14590 2100 14642
rect 2044 14578 2100 14590
rect 3052 14530 3108 14542
rect 3052 14478 3054 14530
rect 3106 14478 3108 14530
rect 3052 14308 3108 14478
rect 14364 14420 14420 14430
rect 14364 14326 14420 14364
rect 14812 14420 14868 14430
rect 3052 14242 3108 14252
rect 3612 14308 3668 14318
rect 3612 14214 3668 14252
rect 14028 14308 14084 14318
rect 14028 14214 14084 14252
rect 2156 14084 2212 14094
rect 2156 13858 2212 14028
rect 2156 13806 2158 13858
rect 2210 13806 2212 13858
rect 2156 13794 2212 13806
rect 12460 13858 12516 13870
rect 12460 13806 12462 13858
rect 12514 13806 12516 13858
rect 3052 13746 3108 13758
rect 3052 13694 3054 13746
rect 3106 13694 3108 13746
rect 3052 13636 3108 13694
rect 12012 13748 12068 13758
rect 12012 13654 12068 13692
rect 3052 13570 3108 13580
rect 3612 13636 3668 13646
rect 3612 13542 3668 13580
rect 2044 13412 2100 13422
rect 2044 13074 2100 13356
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 2044 13022 2046 13074
rect 2098 13022 2100 13074
rect 2044 13010 2100 13022
rect 3052 12962 3108 12974
rect 3052 12910 3054 12962
rect 3106 12910 3108 12962
rect 2156 12740 2212 12750
rect 2156 12290 2212 12684
rect 3052 12740 3108 12910
rect 3052 12674 3108 12684
rect 3612 12740 3668 12750
rect 3612 12646 3668 12684
rect 12012 12738 12068 12750
rect 12012 12686 12014 12738
rect 12066 12686 12068 12738
rect 2156 12238 2158 12290
rect 2210 12238 2212 12290
rect 2156 12226 2212 12238
rect 3052 12292 3108 12302
rect 3052 12178 3108 12236
rect 3052 12126 3054 12178
rect 3106 12126 3108 12178
rect 3052 12114 3108 12126
rect 3612 12292 3668 12302
rect 2044 12068 2100 12078
rect 2044 11506 2100 12012
rect 2044 11454 2046 11506
rect 2098 11454 2100 11506
rect 2044 11442 2100 11454
rect 3052 11508 3108 11518
rect 3052 11394 3108 11452
rect 3612 11506 3668 12236
rect 11340 12290 11396 12302
rect 11340 12238 11342 12290
rect 11394 12238 11396 12290
rect 4844 12178 4900 12190
rect 4844 12126 4846 12178
rect 4898 12126 4900 12178
rect 3612 11454 3614 11506
rect 3666 11454 3668 11506
rect 3612 11442 3668 11454
rect 3836 12066 3892 12078
rect 3836 12014 3838 12066
rect 3890 12014 3892 12066
rect 3052 11342 3054 11394
rect 3106 11342 3108 11394
rect 3052 11330 3108 11342
rect 3836 11396 3892 12014
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4060 11508 4116 11518
rect 4060 11414 4116 11452
rect 3836 11330 3892 11340
rect 4844 11284 4900 12126
rect 11340 11508 11396 12238
rect 11676 12180 11732 12190
rect 12012 12180 12068 12686
rect 12460 12740 12516 13806
rect 13356 13858 13412 13870
rect 13356 13806 13358 13858
rect 13410 13806 13412 13858
rect 12796 13748 12852 13758
rect 12796 13654 12852 13692
rect 13356 13636 13412 13806
rect 13356 13570 13412 13580
rect 13692 13746 13748 13758
rect 13692 13694 13694 13746
rect 13746 13694 13748 13746
rect 13692 13524 13748 13694
rect 12460 12674 12516 12684
rect 13020 12738 13076 12750
rect 13020 12686 13022 12738
rect 13074 12686 13076 12738
rect 12236 12292 12292 12302
rect 12236 12198 12292 12236
rect 11676 12178 12068 12180
rect 11676 12126 11678 12178
rect 11730 12126 12068 12178
rect 11676 12124 12068 12126
rect 12572 12180 12628 12190
rect 12684 12180 12740 12190
rect 12572 12178 12684 12180
rect 12572 12126 12574 12178
rect 12626 12126 12684 12178
rect 12572 12124 12684 12126
rect 11676 12114 11732 12124
rect 11340 11442 11396 11452
rect 4844 11218 4900 11228
rect 10780 11284 10836 11294
rect 10780 11190 10836 11228
rect 11116 11284 11172 11294
rect 11676 11284 11732 11294
rect 11116 11282 11732 11284
rect 11116 11230 11118 11282
rect 11170 11230 11678 11282
rect 11730 11230 11732 11282
rect 11116 11228 11732 11230
rect 11116 11218 11172 11228
rect 2156 10724 2212 10734
rect 2156 10630 2212 10668
rect 3052 10724 3108 10734
rect 3052 10610 3108 10668
rect 10108 10724 10164 10734
rect 10108 10630 10164 10668
rect 11452 10724 11508 10734
rect 11452 10630 11508 10668
rect 3052 10558 3054 10610
rect 3106 10558 3108 10610
rect 3052 10546 3108 10558
rect 10444 10612 10500 10622
rect 11116 10612 11172 10622
rect 10444 10610 11172 10612
rect 10444 10558 10446 10610
rect 10498 10558 11118 10610
rect 11170 10558 11172 10610
rect 10444 10556 11172 10558
rect 10444 10546 10500 10556
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 2044 10052 2100 10062
rect 2044 9938 2100 9996
rect 2044 9886 2046 9938
rect 2098 9886 2100 9938
rect 2044 9874 2100 9886
rect 3052 9826 3108 9838
rect 3052 9774 3054 9826
rect 3106 9774 3108 9826
rect 3052 9716 3108 9774
rect 9660 9826 9716 9838
rect 9660 9774 9662 9826
rect 9714 9774 9716 9826
rect 3052 9650 3108 9660
rect 9436 9716 9492 9726
rect 9436 9622 9492 9660
rect 9660 9716 9716 9774
rect 2156 9380 2212 9390
rect 2156 9154 2212 9324
rect 2156 9102 2158 9154
rect 2210 9102 2212 9154
rect 2156 9090 2212 9102
rect 3052 9156 3108 9166
rect 3052 9042 3108 9100
rect 8652 9156 8708 9166
rect 8652 9062 8708 9100
rect 3052 8990 3054 9042
rect 3106 8990 3108 9042
rect 3052 8978 3108 8990
rect 8988 9044 9044 9054
rect 2044 8708 2100 8718
rect 2044 8370 2100 8652
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 8988 8428 9044 8988
rect 2044 8318 2046 8370
rect 2098 8318 2100 8370
rect 2044 8306 2100 8318
rect 8876 8372 9044 8428
rect 3052 8258 3108 8270
rect 3052 8206 3054 8258
rect 3106 8206 3108 8258
rect 3052 8148 3108 8206
rect 3052 8082 3108 8092
rect 7980 8148 8036 8158
rect 7980 8054 8036 8092
rect 8316 8148 8372 8158
rect 8316 8054 8372 8092
rect 2156 8036 2212 8046
rect 2156 7586 2212 7980
rect 2156 7534 2158 7586
rect 2210 7534 2212 7586
rect 2156 7522 2212 7534
rect 3052 7588 3108 7598
rect 3052 7474 3108 7532
rect 6524 7586 6580 7598
rect 6524 7534 6526 7586
rect 6578 7534 6580 7586
rect 3052 7422 3054 7474
rect 3106 7422 3108 7474
rect 3052 7410 3108 7422
rect 4844 7474 4900 7486
rect 4844 7422 4846 7474
rect 4898 7422 4900 7474
rect 2156 7364 2212 7374
rect 2156 6690 2212 7308
rect 3836 7362 3892 7374
rect 3836 7310 3838 7362
rect 3890 7310 3892 7362
rect 2156 6638 2158 6690
rect 2210 6638 2212 6690
rect 2156 6626 2212 6638
rect 3052 6804 3108 6814
rect 3052 6690 3108 6748
rect 3052 6638 3054 6690
rect 3106 6638 3108 6690
rect 3052 6626 3108 6638
rect 3836 6692 3892 7310
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 3836 6626 3892 6636
rect 4844 6580 4900 7422
rect 6524 6804 6580 7534
rect 7420 7588 7476 7598
rect 7420 7494 7476 7532
rect 8764 7588 8820 7598
rect 8764 7494 8820 7532
rect 6860 7476 6916 7486
rect 7644 7476 7700 7486
rect 6860 7474 7028 7476
rect 6860 7422 6862 7474
rect 6914 7422 7028 7474
rect 6860 7420 7028 7422
rect 6860 7410 6916 7420
rect 6524 6738 6580 6748
rect 6972 6692 7028 7420
rect 4844 6514 4900 6524
rect 5964 6580 6020 6590
rect 5964 6486 6020 6524
rect 6300 6580 6356 6590
rect 6300 6486 6356 6524
rect 6860 6580 6916 6590
rect 2156 6020 2212 6030
rect 2156 5926 2212 5964
rect 3052 6020 3108 6030
rect 3052 5906 3108 5964
rect 5292 6020 5348 6030
rect 5292 5926 5348 5964
rect 6748 6020 6804 6030
rect 6748 5926 6804 5964
rect 3052 5854 3054 5906
rect 3106 5854 3108 5906
rect 3052 5842 3108 5854
rect 5628 5908 5684 5918
rect 6412 5908 6468 5918
rect 5628 5906 6468 5908
rect 5628 5854 5630 5906
rect 5682 5854 6414 5906
rect 6466 5854 6468 5906
rect 5628 5852 6468 5854
rect 5628 5842 5684 5852
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 2044 5348 2100 5358
rect 2044 5234 2100 5292
rect 2044 5182 2046 5234
rect 2098 5182 2100 5234
rect 2044 5170 2100 5182
rect 3052 5122 3108 5134
rect 3052 5070 3054 5122
rect 3106 5070 3108 5122
rect 3052 5012 3108 5070
rect 3052 4946 3108 4956
rect 4620 5012 4676 5022
rect 4620 4918 4676 4956
rect 4956 5012 5012 5022
rect 4956 4918 5012 4956
rect 5740 5012 5796 5022
rect 5740 4564 5796 4956
rect 6076 4900 6132 4910
rect 6076 4806 6132 4844
rect 5852 4564 5908 4574
rect 5740 4562 5908 4564
rect 5740 4510 5854 4562
rect 5906 4510 5908 4562
rect 5740 4508 5908 4510
rect 5852 4498 5908 4508
rect 5516 4338 5572 4350
rect 5516 4286 5518 4338
rect 5570 4286 5572 4338
rect 5068 4228 5124 4238
rect 5516 4228 5572 4286
rect 5068 4226 5572 4228
rect 5068 4174 5070 4226
rect 5122 4174 5572 4226
rect 5068 4172 5572 4174
rect 5068 4162 5124 4172
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 5068 3444 5124 3454
rect 5068 3350 5124 3388
rect 5292 800 5348 4172
rect 5964 3554 6020 3566
rect 5964 3502 5966 3554
rect 6018 3502 6020 3554
rect 5964 3444 6020 3502
rect 5964 800 6020 3388
rect 6188 3444 6244 3454
rect 6300 3444 6356 5852
rect 6412 5842 6468 5852
rect 6860 4562 6916 6524
rect 6860 4510 6862 4562
rect 6914 4510 6916 4562
rect 6860 4498 6916 4510
rect 6412 4340 6468 4350
rect 6972 4340 7028 6636
rect 7196 6468 7252 6478
rect 7196 6374 7252 6412
rect 7644 6132 7700 7420
rect 8428 7476 8484 7486
rect 8428 7382 8484 7420
rect 7756 6692 7812 6702
rect 7756 6598 7812 6636
rect 8092 6580 8148 6590
rect 8092 6486 8148 6524
rect 7644 6076 7812 6132
rect 6412 4226 6468 4284
rect 6412 4174 6414 4226
rect 6466 4174 6468 4226
rect 6412 3780 6468 4174
rect 6748 4284 7028 4340
rect 7084 4340 7140 4350
rect 6412 3724 6692 3780
rect 6188 3442 6356 3444
rect 6188 3390 6190 3442
rect 6242 3390 6356 3442
rect 6188 3388 6356 3390
rect 6188 3378 6244 3388
rect 6636 800 6692 3724
rect 6748 3442 6804 4284
rect 7084 4246 7140 4284
rect 7644 4228 7700 4238
rect 7308 4226 7700 4228
rect 7308 4174 7646 4226
rect 7698 4174 7700 4226
rect 7308 4172 7700 4174
rect 6748 3390 6750 3442
rect 6802 3390 6804 3442
rect 6748 3378 6804 3390
rect 7084 3444 7140 3454
rect 7308 3444 7364 4172
rect 7644 4162 7700 4172
rect 7084 3442 7364 3444
rect 7084 3390 7086 3442
rect 7138 3390 7364 3442
rect 7084 3388 7364 3390
rect 7084 3378 7140 3388
rect 7308 800 7364 3388
rect 7644 3444 7700 3454
rect 7756 3444 7812 6076
rect 8092 4228 8148 4238
rect 8652 4228 8708 4238
rect 7644 3442 7812 3444
rect 7644 3390 7646 3442
rect 7698 3390 7812 3442
rect 7644 3388 7812 3390
rect 7980 4226 8148 4228
rect 7980 4174 8094 4226
rect 8146 4174 8148 4226
rect 7980 4172 8148 4174
rect 7980 3442 8036 4172
rect 8092 4162 8148 4172
rect 8540 4226 8708 4228
rect 8540 4174 8654 4226
rect 8706 4174 8708 4226
rect 8540 4172 8708 4174
rect 7980 3390 7982 3442
rect 8034 3390 8036 3442
rect 7644 3378 7700 3388
rect 7980 800 8036 3390
rect 8540 3444 8596 4172
rect 8652 4162 8708 4172
rect 8540 3350 8596 3388
rect 8876 3330 8932 8372
rect 9100 8148 9156 8158
rect 9100 8054 9156 8092
rect 9436 8036 9492 8046
rect 9436 7942 9492 7980
rect 8876 3278 8878 3330
rect 8930 3278 8932 3330
rect 8876 3266 8932 3278
rect 8988 4340 9044 4350
rect 8988 4226 9044 4284
rect 8988 4174 8990 4226
rect 9042 4174 9044 4226
rect 8988 2884 9044 4174
rect 8652 2828 9044 2884
rect 9324 3444 9380 3454
rect 8652 800 8708 2828
rect 9324 800 9380 3388
rect 9660 3332 9716 9660
rect 10556 9716 10612 9726
rect 10556 9622 10612 9660
rect 10892 9604 10948 9614
rect 10892 9510 10948 9548
rect 10220 9156 10276 9166
rect 10220 9062 10276 9100
rect 9884 9044 9940 9054
rect 9884 8950 9940 8988
rect 9772 8148 9828 8158
rect 9772 4562 9828 8092
rect 9772 4510 9774 4562
rect 9826 4510 9828 4562
rect 9772 4498 9828 4510
rect 10332 4898 10388 4910
rect 10332 4846 10334 4898
rect 10386 4846 10388 4898
rect 9996 4340 10052 4350
rect 9996 4246 10052 4284
rect 10108 3444 10164 3454
rect 10332 3444 10388 4846
rect 9996 3442 10388 3444
rect 9996 3390 10110 3442
rect 10162 3390 10388 3442
rect 9996 3388 10388 3390
rect 10668 4226 10724 4238
rect 10668 4174 10670 4226
rect 10722 4174 10724 4226
rect 10668 3442 10724 4174
rect 10668 3390 10670 3442
rect 10722 3390 10724 3442
rect 9772 3332 9828 3342
rect 9660 3330 9828 3332
rect 9660 3278 9774 3330
rect 9826 3278 9828 3330
rect 9660 3276 9828 3278
rect 9772 3266 9828 3276
rect 9996 800 10052 3388
rect 10108 3378 10164 3388
rect 10668 800 10724 3390
rect 11004 3330 11060 10556
rect 11116 10546 11172 10556
rect 11564 9716 11620 11228
rect 11676 11218 11732 11228
rect 11788 10388 11844 12124
rect 12572 12114 12628 12124
rect 12572 11282 12628 11294
rect 12572 11230 12574 11282
rect 12626 11230 12628 11282
rect 12012 11172 12068 11182
rect 12012 11078 12068 11116
rect 12236 10500 12292 10510
rect 12572 10500 12628 11230
rect 12236 10498 12628 10500
rect 12236 10446 12238 10498
rect 12290 10446 12628 10498
rect 12236 10444 12628 10446
rect 12236 10388 12292 10444
rect 11788 10332 12292 10388
rect 11900 9940 11956 10332
rect 11564 9650 11620 9660
rect 11676 9884 11956 9940
rect 11564 4338 11620 4350
rect 11564 4286 11566 4338
rect 11618 4286 11620 4338
rect 11116 4228 11172 4238
rect 11564 4228 11620 4286
rect 11116 4226 11620 4228
rect 11116 4174 11118 4226
rect 11170 4174 11620 4226
rect 11116 4172 11620 4174
rect 11116 4162 11172 4172
rect 11004 3278 11006 3330
rect 11058 3278 11060 3330
rect 11004 3266 11060 3278
rect 11340 800 11396 4172
rect 11564 3332 11620 3342
rect 11676 3332 11732 9884
rect 11900 9716 11956 9726
rect 11900 4562 11956 9660
rect 12684 8428 12740 12124
rect 13020 12180 13076 12686
rect 13580 12292 13636 12302
rect 13580 12198 13636 12236
rect 13020 12114 13076 12124
rect 13244 12180 13300 12190
rect 13244 12086 13300 12124
rect 12908 11284 12964 11294
rect 12908 11190 12964 11228
rect 12684 8372 12852 8428
rect 12124 4900 12180 4910
rect 11900 4510 11902 4562
rect 11954 4510 11956 4562
rect 11900 4498 11956 4510
rect 12012 4898 12180 4900
rect 12012 4846 12126 4898
rect 12178 4846 12180 4898
rect 12012 4844 12180 4846
rect 11900 3444 11956 3454
rect 12012 3444 12068 4844
rect 12124 4834 12180 4844
rect 12684 4226 12740 4238
rect 12684 4174 12686 4226
rect 12738 4174 12740 4226
rect 12572 3556 12628 3566
rect 12684 3556 12740 4174
rect 12572 3554 12740 3556
rect 12572 3502 12574 3554
rect 12626 3502 12740 3554
rect 12572 3500 12740 3502
rect 12572 3490 12628 3500
rect 11900 3442 12068 3444
rect 11900 3390 11902 3442
rect 11954 3390 12068 3442
rect 11900 3388 12068 3390
rect 11900 3378 11956 3388
rect 11564 3330 11732 3332
rect 11564 3278 11566 3330
rect 11618 3278 11732 3330
rect 11564 3276 11732 3278
rect 11564 3266 11620 3276
rect 12012 800 12068 3388
rect 12684 800 12740 3500
rect 12796 3330 12852 8372
rect 13580 4338 13636 4350
rect 13580 4286 13582 4338
rect 13634 4286 13636 4338
rect 13132 4228 13188 4238
rect 13580 4228 13636 4286
rect 13132 4226 13636 4228
rect 13132 4174 13134 4226
rect 13186 4174 13636 4226
rect 13132 4172 13636 4174
rect 13132 4162 13188 4172
rect 12796 3278 12798 3330
rect 12850 3278 12852 3330
rect 12796 3266 12852 3278
rect 13356 800 13412 4172
rect 13692 3330 13748 13468
rect 13916 13748 13972 13758
rect 13916 4562 13972 13692
rect 14140 13634 14196 13646
rect 14140 13582 14142 13634
rect 14194 13582 14196 13634
rect 14140 13524 14196 13582
rect 14140 13458 14196 13468
rect 14028 12180 14084 12190
rect 14028 12086 14084 12124
rect 14812 8428 14868 14364
rect 15708 9268 15764 9278
rect 14812 8372 14980 8428
rect 14252 4900 14308 4910
rect 13916 4510 13918 4562
rect 13970 4510 13972 4562
rect 13916 4498 13972 4510
rect 14028 4898 14308 4900
rect 14028 4846 14254 4898
rect 14306 4846 14308 4898
rect 14028 4844 14308 4846
rect 13692 3278 13694 3330
rect 13746 3278 13748 3330
rect 13692 3266 13748 3278
rect 14028 3442 14084 4844
rect 14252 4834 14308 4844
rect 14028 3390 14030 3442
rect 14082 3390 14084 3442
rect 14028 800 14084 3390
rect 14700 4226 14756 4238
rect 14700 4174 14702 4226
rect 14754 4174 14756 4226
rect 14700 3554 14756 4174
rect 14700 3502 14702 3554
rect 14754 3502 14756 3554
rect 14700 800 14756 3502
rect 14924 3330 14980 8372
rect 15148 4340 15204 4350
rect 15148 4246 15204 4284
rect 15372 4340 15428 4350
rect 14924 3278 14926 3330
rect 14978 3278 14980 3330
rect 14924 3266 14980 3278
rect 15372 800 15428 4284
rect 15596 4340 15652 4350
rect 15596 4246 15652 4284
rect 15596 3554 15652 3566
rect 15596 3502 15598 3554
rect 15650 3502 15652 3554
rect 15596 3108 15652 3502
rect 15708 3388 15764 9212
rect 15820 4564 15876 15092
rect 16268 9268 16324 15148
rect 16268 9202 16324 9212
rect 16380 15204 16436 15214
rect 16044 4900 16100 4910
rect 16044 4898 16324 4900
rect 16044 4846 16046 4898
rect 16098 4846 16324 4898
rect 16044 4844 16324 4846
rect 16044 4834 16100 4844
rect 15932 4564 15988 4574
rect 15820 4562 15988 4564
rect 15820 4510 15934 4562
rect 15986 4510 15988 4562
rect 15820 4508 15988 4510
rect 15932 4498 15988 4508
rect 16268 4116 16324 4844
rect 16044 4060 16324 4116
rect 15708 3332 15876 3388
rect 15820 3330 15876 3332
rect 15820 3278 15822 3330
rect 15874 3278 15876 3330
rect 15820 3266 15876 3278
rect 16044 3108 16100 4060
rect 16380 3330 16436 15148
rect 17052 15202 17108 16828
rect 18060 16884 18116 17500
rect 18060 16818 18116 16828
rect 18284 16882 18340 16894
rect 18284 16830 18286 16882
rect 18338 16830 18340 16882
rect 17724 16772 17780 16782
rect 17612 16770 17780 16772
rect 17612 16718 17726 16770
rect 17778 16718 17780 16770
rect 17612 16716 17780 16718
rect 17612 16212 17668 16716
rect 17724 16706 17780 16716
rect 17276 15876 17332 15886
rect 17276 15782 17332 15820
rect 17052 15150 17054 15202
rect 17106 15150 17108 15202
rect 17052 15148 17108 15150
rect 17612 15204 17668 16156
rect 17724 16322 17780 16334
rect 17724 16270 17726 16322
rect 17778 16270 17780 16322
rect 17724 15876 17780 16270
rect 18284 16100 18340 16830
rect 18508 16884 18564 17500
rect 18620 17490 18676 17500
rect 18956 17554 19012 17836
rect 18956 17502 18958 17554
rect 19010 17502 19012 17554
rect 18956 17490 19012 17502
rect 18620 16996 18676 17006
rect 19068 16996 19124 18396
rect 19628 18340 19684 18350
rect 19516 18338 19684 18340
rect 19516 18286 19630 18338
rect 19682 18286 19684 18338
rect 19516 18284 19684 18286
rect 19404 17444 19460 17454
rect 19516 17444 19572 18284
rect 19628 18274 19684 18284
rect 20076 18338 20132 18508
rect 20076 18286 20078 18338
rect 20130 18286 20132 18338
rect 19404 17442 19572 17444
rect 19404 17390 19406 17442
rect 19458 17390 19572 17442
rect 19404 17388 19572 17390
rect 19628 17780 19684 17790
rect 19404 17108 19460 17388
rect 19628 17108 19684 17724
rect 20076 17666 20132 18286
rect 20300 17668 20356 19964
rect 20636 20020 20692 20526
rect 21532 20580 21588 21644
rect 21644 21634 21700 21644
rect 21868 21586 21924 21598
rect 21868 21534 21870 21586
rect 21922 21534 21924 21586
rect 21644 20692 21700 20702
rect 21644 20598 21700 20636
rect 21532 20514 21588 20524
rect 21868 20580 21924 21534
rect 22428 21476 22484 22204
rect 22988 22260 23044 22270
rect 22988 22166 23044 22204
rect 23324 22148 23380 22158
rect 23324 22054 23380 22092
rect 23660 21586 23716 21598
rect 23660 21534 23662 21586
rect 23714 21534 23716 21586
rect 22652 21476 22708 21486
rect 22428 21474 22708 21476
rect 22428 21422 22654 21474
rect 22706 21422 22708 21474
rect 22428 21420 22708 21422
rect 21196 20130 21252 20142
rect 21196 20078 21198 20130
rect 21250 20078 21252 20130
rect 20636 19954 20692 19964
rect 20860 20020 20916 20030
rect 20860 19926 20916 19964
rect 21196 20020 21252 20078
rect 21196 19954 21252 19964
rect 21756 19906 21812 19918
rect 21756 19854 21758 19906
rect 21810 19854 21812 19906
rect 20524 19234 20580 19246
rect 20524 19182 20526 19234
rect 20578 19182 20580 19234
rect 20524 19124 20580 19182
rect 20524 18900 20580 19068
rect 21644 19122 21700 19134
rect 21644 19070 21646 19122
rect 21698 19070 21700 19122
rect 20748 19012 20804 19022
rect 20748 18918 20804 18956
rect 20412 18564 20468 18574
rect 20524 18564 20580 18844
rect 20468 18508 20580 18564
rect 20860 18676 20916 18686
rect 20412 18498 20468 18508
rect 20748 18452 20804 18462
rect 20524 18450 20804 18452
rect 20524 18398 20750 18450
rect 20802 18398 20804 18450
rect 20524 18396 20804 18398
rect 20524 17892 20580 18396
rect 20748 18386 20804 18396
rect 20076 17614 20078 17666
rect 20130 17614 20132 17666
rect 20076 17444 20132 17614
rect 20076 17378 20132 17388
rect 20188 17666 20356 17668
rect 20188 17614 20302 17666
rect 20354 17614 20356 17666
rect 20188 17612 20356 17614
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19852 17108 19908 17118
rect 19628 17106 19908 17108
rect 19628 17054 19854 17106
rect 19906 17054 19908 17106
rect 19628 17052 19908 17054
rect 19404 16996 19460 17052
rect 19852 17042 19908 17052
rect 19068 16940 19460 16996
rect 18620 16902 18676 16940
rect 18508 16322 18564 16828
rect 18508 16270 18510 16322
rect 18562 16270 18564 16322
rect 18508 16258 18564 16270
rect 18956 16212 19012 16222
rect 18956 16118 19012 16156
rect 18172 16098 18340 16100
rect 18172 16046 18286 16098
rect 18338 16046 18340 16098
rect 18172 16044 18340 16046
rect 17724 15874 17892 15876
rect 17724 15822 17726 15874
rect 17778 15822 17892 15874
rect 17724 15820 17892 15822
rect 17724 15810 17780 15820
rect 17724 15204 17780 15214
rect 17612 15148 17724 15204
rect 17836 15204 17892 15820
rect 18172 15204 18228 16044
rect 18284 16034 18340 16044
rect 18732 16098 18788 16110
rect 18732 16046 18734 16098
rect 18786 16046 18788 16098
rect 18732 15876 18788 16046
rect 19068 16100 19124 16110
rect 19068 16006 19124 16044
rect 18732 15810 18788 15820
rect 17836 15202 18228 15204
rect 17836 15150 18174 15202
rect 18226 15150 18228 15202
rect 17836 15148 18228 15150
rect 17052 15092 17556 15148
rect 17724 15110 17780 15148
rect 17052 4340 17108 4350
rect 17052 4246 17108 4284
rect 17388 4340 17444 4350
rect 16604 4226 16660 4238
rect 16604 4174 16606 4226
rect 16658 4174 16660 4226
rect 16604 3554 16660 4174
rect 16604 3502 16606 3554
rect 16658 3502 16660 3554
rect 16604 3388 16660 3502
rect 16604 3332 16772 3388
rect 16380 3278 16382 3330
rect 16434 3278 16436 3330
rect 16380 3266 16436 3278
rect 15596 3052 16100 3108
rect 16044 800 16100 3052
rect 16716 800 16772 3332
rect 17388 800 17444 4284
rect 17500 3388 17556 15092
rect 18060 4562 18116 15148
rect 18172 15138 18228 15148
rect 18060 4510 18062 4562
rect 18114 4510 18116 4562
rect 18060 4498 18116 4510
rect 18172 4898 18228 4910
rect 18172 4846 18174 4898
rect 18226 4846 18228 4898
rect 17724 4340 17780 4350
rect 17724 4246 17780 4284
rect 17948 3556 18004 3566
rect 18172 3556 18228 4846
rect 18844 4228 18900 4238
rect 17948 3554 18228 3556
rect 17948 3502 17950 3554
rect 18002 3502 18228 3554
rect 17948 3500 18228 3502
rect 18620 4226 18900 4228
rect 18620 4174 18846 4226
rect 18898 4174 18900 4226
rect 18620 4172 18900 4174
rect 18620 3554 18676 4172
rect 18844 4162 18900 4172
rect 18620 3502 18622 3554
rect 18674 3502 18676 3554
rect 17948 3490 18004 3500
rect 17500 3332 17668 3388
rect 17612 3330 17668 3332
rect 17612 3278 17614 3330
rect 17666 3278 17668 3330
rect 17612 3266 17668 3278
rect 18060 800 18116 3500
rect 18620 3388 18676 3502
rect 19180 3388 19236 16940
rect 19516 16884 19572 16894
rect 19404 16882 19572 16884
rect 19404 16830 19518 16882
rect 19570 16830 19572 16882
rect 19404 16828 19572 16830
rect 19404 16212 19460 16828
rect 19516 16818 19572 16828
rect 19628 16772 19684 16782
rect 19628 16212 19684 16716
rect 19404 16146 19460 16156
rect 19516 16156 19684 16212
rect 19292 15876 19348 15886
rect 19292 15538 19348 15820
rect 19292 15486 19294 15538
rect 19346 15486 19348 15538
rect 19292 15474 19348 15486
rect 18620 3332 18788 3388
rect 18732 800 18788 3332
rect 18844 3332 18900 3342
rect 18956 3332 19236 3388
rect 19404 4226 19460 4238
rect 19404 4174 19406 4226
rect 19458 4174 19460 4226
rect 19404 3554 19460 4174
rect 19404 3502 19406 3554
rect 19458 3502 19460 3554
rect 18844 3330 19012 3332
rect 18844 3278 18846 3330
rect 18898 3278 19012 3330
rect 18844 3276 19012 3278
rect 18844 3266 18900 3276
rect 19404 800 19460 3502
rect 19516 3332 19572 16156
rect 19628 15986 19684 15998
rect 19628 15934 19630 15986
rect 19682 15934 19684 15986
rect 19628 15876 19684 15934
rect 19628 15810 19684 15820
rect 19964 15876 20020 15914
rect 19964 15810 20020 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15148 20244 17612
rect 20300 17556 20356 17612
rect 20300 17490 20356 17500
rect 20412 17890 20580 17892
rect 20412 17838 20526 17890
rect 20578 17838 20580 17890
rect 20412 17836 20580 17838
rect 20300 17108 20356 17118
rect 20412 17108 20468 17836
rect 20524 17826 20580 17836
rect 20748 17892 20804 17902
rect 20860 17892 20916 18620
rect 21532 18676 21588 18686
rect 21644 18676 21700 19070
rect 21756 18900 21812 19854
rect 21756 18834 21812 18844
rect 21588 18620 21700 18676
rect 20748 17890 20916 17892
rect 20748 17838 20750 17890
rect 20802 17838 20916 17890
rect 20748 17836 20916 17838
rect 21084 18562 21140 18574
rect 21084 18510 21086 18562
rect 21138 18510 21140 18562
rect 21532 18544 21588 18620
rect 20356 17052 20468 17108
rect 20636 17444 20692 17454
rect 20300 16976 20356 17052
rect 20188 15092 20580 15148
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19852 4340 19908 4350
rect 20300 4340 20356 4350
rect 19852 4246 19908 4284
rect 20188 4284 20300 4340
rect 19740 3332 19796 3342
rect 19516 3330 19796 3332
rect 19516 3278 19742 3330
rect 19794 3278 19796 3330
rect 19516 3276 19796 3278
rect 19740 3266 19796 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 2996 20244 4284
rect 20300 4246 20356 4284
rect 20300 3332 20356 3342
rect 20524 3332 20580 15092
rect 20636 4562 20692 17388
rect 20748 17106 20804 17836
rect 21084 17668 21140 18510
rect 21084 17602 21140 17612
rect 20860 17554 20916 17566
rect 20860 17502 20862 17554
rect 20914 17502 20916 17554
rect 20860 17220 20916 17502
rect 21532 17556 21588 17566
rect 21532 17462 21588 17500
rect 20860 17154 20916 17164
rect 20748 17054 20750 17106
rect 20802 17054 20804 17106
rect 20748 16772 20804 17054
rect 21532 16884 21588 16894
rect 21532 16790 21588 16828
rect 21868 16882 21924 20524
rect 21980 20690 22036 20702
rect 21980 20638 21982 20690
rect 22034 20638 22036 20690
rect 21980 20188 22036 20638
rect 22428 20580 22484 20590
rect 22428 20486 22484 20524
rect 21980 20132 22260 20188
rect 22204 19908 22260 20132
rect 21980 19124 22036 19134
rect 21980 19030 22036 19068
rect 21980 18900 22036 18910
rect 21980 17778 22036 18844
rect 21980 17726 21982 17778
rect 22034 17726 22036 17778
rect 21980 17714 22036 17726
rect 21868 16830 21870 16882
rect 21922 16830 21924 16882
rect 20748 16706 20804 16716
rect 20860 4900 20916 4910
rect 20636 4510 20638 4562
rect 20690 4510 20692 4562
rect 20636 4498 20692 4510
rect 20748 4898 20916 4900
rect 20748 4846 20862 4898
rect 20914 4846 20916 4898
rect 20748 4844 20916 4846
rect 20636 3556 20692 3566
rect 20748 3556 20804 4844
rect 20860 4834 20916 4844
rect 21196 4340 21252 4350
rect 21196 4246 21252 4284
rect 21420 4340 21476 4350
rect 20636 3554 20804 3556
rect 20636 3502 20638 3554
rect 20690 3502 20804 3554
rect 20636 3500 20804 3502
rect 20636 3490 20692 3500
rect 20300 3330 20580 3332
rect 20300 3278 20302 3330
rect 20354 3278 20580 3330
rect 20300 3276 20580 3278
rect 20300 3266 20356 3276
rect 20076 2940 20244 2996
rect 20076 800 20132 2940
rect 20748 800 20804 3500
rect 21420 800 21476 4284
rect 21644 4340 21700 4350
rect 21644 4246 21700 4284
rect 21644 3556 21700 3566
rect 21644 3462 21700 3500
rect 21868 3330 21924 16830
rect 22204 16772 22260 19852
rect 22428 16884 22484 16894
rect 22316 16772 22372 16782
rect 21980 16716 22316 16772
rect 21980 4562 22036 16716
rect 22316 16640 22372 16716
rect 22428 15148 22484 16828
rect 22652 16884 22708 21420
rect 23100 21474 23156 21486
rect 23100 21422 23102 21474
rect 23154 21422 23156 21474
rect 23100 20580 23156 21422
rect 23100 20514 23156 20524
rect 23212 20690 23268 20702
rect 23212 20638 23214 20690
rect 23266 20638 23268 20690
rect 22876 19908 22932 19918
rect 23212 19908 23268 20638
rect 23548 20580 23604 20590
rect 23548 20486 23604 20524
rect 23660 20468 23716 21534
rect 23660 20188 23716 20412
rect 22932 19852 23268 19908
rect 23548 20132 23716 20188
rect 23772 20188 23828 23100
rect 23996 23044 24052 23548
rect 24780 23156 24836 23166
rect 24780 23062 24836 23100
rect 24332 23044 24388 23054
rect 23996 23042 24388 23044
rect 23996 22990 24334 23042
rect 24386 22990 24388 23042
rect 23996 22988 24388 22990
rect 23996 21700 24052 21710
rect 23996 21606 24052 21644
rect 23772 20132 23940 20188
rect 22876 19814 22932 19852
rect 23212 17332 23268 17342
rect 22988 17108 23044 17118
rect 22652 16818 22708 16828
rect 22876 17106 23044 17108
rect 22876 17054 22990 17106
rect 23042 17054 23044 17106
rect 22876 17052 23044 17054
rect 22876 16322 22932 17052
rect 22988 17042 23044 17052
rect 22988 16884 23044 16894
rect 22988 16790 23044 16828
rect 23100 16660 23156 16670
rect 23100 16566 23156 16604
rect 22876 16270 22878 16322
rect 22930 16270 22932 16322
rect 22876 16258 22932 16270
rect 23212 16322 23268 17276
rect 23324 16772 23380 16782
rect 23324 16678 23380 16716
rect 23548 16770 23604 20132
rect 23548 16718 23550 16770
rect 23602 16718 23604 16770
rect 23548 16706 23604 16718
rect 23212 16270 23214 16322
rect 23266 16270 23268 16322
rect 23212 16258 23268 16270
rect 23884 16660 23940 20132
rect 24332 17108 24388 22988
rect 25564 23044 25620 23660
rect 25788 23716 25844 23726
rect 25788 23622 25844 23660
rect 25900 23492 25956 24556
rect 26348 24500 26404 25342
rect 26236 24498 26404 24500
rect 26236 24446 26350 24498
rect 26402 24446 26404 24498
rect 26236 24444 26404 24446
rect 25788 23436 25956 23492
rect 26012 23604 26068 23614
rect 25564 23042 25732 23044
rect 25564 22990 25566 23042
rect 25618 22990 25732 23042
rect 25564 22988 25732 22990
rect 25564 22978 25620 22988
rect 25452 17556 25508 17566
rect 24332 17042 24388 17052
rect 24892 17108 24948 17118
rect 22652 16100 22708 16110
rect 22652 16006 22708 16044
rect 23884 15874 23940 16604
rect 23884 15822 23886 15874
rect 23938 15822 23940 15874
rect 23884 15148 23940 15822
rect 21980 4510 21982 4562
rect 22034 4510 22036 4562
rect 21980 4498 22036 4510
rect 22316 15092 22484 15148
rect 23660 15092 23940 15148
rect 24444 16884 24500 16894
rect 24892 16884 24948 17052
rect 21868 3278 21870 3330
rect 21922 3278 21924 3330
rect 21868 3266 21924 3278
rect 22092 3556 22148 3566
rect 22092 800 22148 3500
rect 22316 3332 22372 15092
rect 22428 4226 22484 4238
rect 22428 4174 22430 4226
rect 22482 4174 22484 4226
rect 22428 3556 22484 4174
rect 22876 4226 22932 4238
rect 22876 4174 22878 4226
rect 22930 4174 22932 4226
rect 22428 3490 22484 3500
rect 22764 3556 22820 3566
rect 22876 3556 22932 4174
rect 22764 3554 22932 3556
rect 22764 3502 22766 3554
rect 22818 3502 22932 3554
rect 22764 3500 22932 3502
rect 23436 4226 23492 4238
rect 23436 4174 23438 4226
rect 23490 4174 23492 4226
rect 23436 3554 23492 4174
rect 23436 3502 23438 3554
rect 23490 3502 23492 3554
rect 22428 3332 22484 3342
rect 22316 3330 22484 3332
rect 22316 3278 22430 3330
rect 22482 3278 22484 3330
rect 22316 3276 22484 3278
rect 22428 3266 22484 3276
rect 22764 800 22820 3500
rect 23436 800 23492 3502
rect 23660 3330 23716 15092
rect 23884 4340 23940 4350
rect 23884 4246 23940 4284
rect 24108 4340 24164 4350
rect 23660 3278 23662 3330
rect 23714 3278 23716 3330
rect 23660 3266 23716 3278
rect 24108 800 24164 4284
rect 24332 4340 24388 4350
rect 24332 4246 24388 4284
rect 24444 3388 24500 16828
rect 24668 16882 24948 16884
rect 24668 16830 24894 16882
rect 24946 16830 24948 16882
rect 24668 16828 24948 16830
rect 24668 4562 24724 16828
rect 24892 16818 24948 16828
rect 24668 4510 24670 4562
rect 24722 4510 24724 4562
rect 24668 4498 24724 4510
rect 24780 4898 24836 4910
rect 24780 4846 24782 4898
rect 24834 4846 24836 4898
rect 24556 3556 24612 3566
rect 24780 3556 24836 4846
rect 24556 3554 24836 3556
rect 24556 3502 24558 3554
rect 24610 3502 24836 3554
rect 24556 3500 24836 3502
rect 24556 3490 24612 3500
rect 24220 3332 24500 3388
rect 24220 3330 24276 3332
rect 24220 3278 24222 3330
rect 24274 3278 24276 3330
rect 24220 3266 24276 3278
rect 24780 800 24836 3500
rect 25452 3330 25508 17500
rect 25676 16884 25732 22988
rect 25788 17556 25844 23436
rect 26012 23378 26068 23548
rect 26012 23326 26014 23378
rect 26066 23326 26068 23378
rect 26012 23314 26068 23326
rect 25788 17462 25844 17500
rect 26124 17778 26180 17790
rect 26124 17726 26126 17778
rect 26178 17726 26180 17778
rect 26012 17444 26068 17482
rect 26012 17378 26068 17388
rect 26012 17220 26068 17230
rect 25788 17108 25844 17118
rect 25788 16994 25844 17052
rect 25788 16942 25790 16994
rect 25842 16942 25844 16994
rect 25788 16930 25844 16942
rect 26012 16994 26068 17164
rect 26012 16942 26014 16994
rect 26066 16942 26068 16994
rect 26012 16930 26068 16942
rect 26124 16884 26180 17726
rect 26236 17444 26292 24444
rect 26348 24434 26404 24444
rect 26460 25396 26516 26124
rect 26348 23826 26404 23838
rect 26348 23774 26350 23826
rect 26402 23774 26404 23826
rect 26348 23604 26404 23774
rect 26348 23538 26404 23548
rect 26236 17378 26292 17388
rect 26236 16884 26292 16894
rect 26124 16882 26292 16884
rect 26124 16830 26238 16882
rect 26290 16830 26292 16882
rect 26124 16828 26292 16830
rect 25676 16790 25732 16828
rect 26236 16818 26292 16828
rect 26012 4898 26068 4910
rect 26012 4846 26014 4898
rect 26066 4846 26068 4898
rect 25900 4340 25956 4350
rect 25900 4246 25956 4284
rect 25788 3556 25844 3566
rect 26012 3556 26068 4846
rect 25788 3554 26068 3556
rect 25788 3502 25790 3554
rect 25842 3502 26068 3554
rect 25788 3500 26068 3502
rect 26124 4340 26180 4350
rect 25788 3388 25844 3500
rect 25452 3278 25454 3330
rect 25506 3278 25508 3330
rect 25452 3266 25508 3278
rect 25676 3332 25844 3388
rect 25676 980 25732 3332
rect 25452 924 25732 980
rect 25452 800 25508 924
rect 26124 800 26180 4284
rect 26348 4340 26404 4350
rect 26348 4246 26404 4284
rect 26460 3388 26516 25340
rect 27132 25396 27188 25406
rect 27132 25302 27188 25340
rect 26684 25284 26740 25294
rect 26684 25190 26740 25228
rect 26572 24610 26628 24622
rect 26572 24558 26574 24610
rect 26626 24558 26628 24610
rect 26572 24498 26628 24558
rect 27020 24612 27076 24622
rect 27020 24518 27076 24556
rect 26572 24446 26574 24498
rect 26626 24446 26628 24498
rect 26572 24434 26628 24446
rect 26684 23828 26740 23838
rect 26684 23734 26740 23772
rect 27020 17556 27076 17566
rect 27020 17462 27076 17500
rect 26572 17444 26628 17454
rect 26572 4564 26628 17388
rect 26684 16884 26740 16894
rect 26684 16790 26740 16828
rect 26684 4564 26740 4574
rect 26572 4562 26740 4564
rect 26572 4510 26686 4562
rect 26738 4510 26740 4562
rect 26572 4508 26740 4510
rect 26684 4498 26740 4508
rect 27132 4228 27188 4238
rect 26796 4226 27188 4228
rect 26796 4174 27134 4226
rect 27186 4174 27188 4226
rect 26796 4172 27188 4174
rect 26684 3556 26740 3566
rect 26796 3556 26852 4172
rect 27132 4162 27188 4172
rect 26684 3554 26852 3556
rect 26684 3502 26686 3554
rect 26738 3502 26852 3554
rect 26684 3500 26852 3502
rect 26684 3490 26740 3500
rect 26236 3332 26516 3388
rect 26236 3330 26404 3332
rect 26236 3278 26350 3330
rect 26402 3278 26404 3330
rect 26236 3276 26404 3278
rect 26348 3266 26404 3276
rect 26796 800 26852 3500
rect 27244 3330 27300 26908
rect 28028 26964 28084 26974
rect 28028 26870 28084 26908
rect 28364 26852 28420 26862
rect 28364 26758 28420 26796
rect 27692 26404 27748 26414
rect 27692 26310 27748 26348
rect 27356 26290 27412 26302
rect 27356 26238 27358 26290
rect 27410 26238 27412 26290
rect 27356 25396 27412 26238
rect 27580 25508 27636 25518
rect 27580 25414 27636 25452
rect 27356 25330 27412 25340
rect 27580 4228 27636 4238
rect 27244 3278 27246 3330
rect 27298 3278 27300 3330
rect 27244 3266 27300 3278
rect 27468 4226 27636 4228
rect 27468 4174 27582 4226
rect 27634 4174 27636 4226
rect 27468 4172 27636 4174
rect 27468 3554 27524 4172
rect 27580 4162 27636 4172
rect 28140 4226 28196 4238
rect 28140 4174 28142 4226
rect 28194 4174 28196 4226
rect 27468 3502 27470 3554
rect 27522 3502 27524 3554
rect 27468 800 27524 3502
rect 28140 3442 28196 4174
rect 28140 3390 28142 3442
rect 28194 3390 28196 3442
rect 28140 800 28196 3390
rect 28476 3330 28532 27804
rect 28588 27794 28644 27804
rect 29372 27748 29428 28476
rect 29596 28466 29652 28476
rect 29260 27746 29428 27748
rect 29260 27694 29374 27746
rect 29426 27694 29428 27746
rect 29260 27692 29428 27694
rect 28812 26964 28868 26974
rect 28812 26870 28868 26908
rect 29260 4564 29316 27692
rect 29372 27682 29428 27692
rect 29708 8428 29764 28588
rect 29932 28420 29988 28430
rect 29932 28326 29988 28364
rect 29820 27860 29876 27870
rect 29820 27766 29876 27804
rect 29484 8372 29764 8428
rect 29372 4564 29428 4574
rect 29260 4562 29428 4564
rect 29260 4510 29374 4562
rect 29426 4510 29428 4562
rect 29260 4508 29428 4510
rect 29372 4498 29428 4508
rect 29036 4338 29092 4350
rect 29036 4286 29038 4338
rect 29090 4286 29092 4338
rect 28588 4228 28644 4238
rect 29036 4228 29092 4286
rect 28588 4226 29092 4228
rect 28588 4174 28590 4226
rect 28642 4174 29092 4226
rect 28588 4172 29092 4174
rect 28588 4162 28644 4172
rect 28476 3278 28478 3330
rect 28530 3278 28532 3330
rect 28476 3266 28532 3278
rect 28812 800 28868 4172
rect 29372 3332 29428 3342
rect 29484 3332 29540 8372
rect 29932 4900 29988 4910
rect 29820 4898 29988 4900
rect 29820 4846 29934 4898
rect 29986 4846 29988 4898
rect 29820 4844 29988 4846
rect 29372 3330 29540 3332
rect 29372 3278 29374 3330
rect 29426 3278 29540 3330
rect 29372 3276 29540 3278
rect 29596 3556 29652 3566
rect 29820 3556 29876 4844
rect 29932 4834 29988 4844
rect 30156 4340 30212 4350
rect 29932 4228 29988 4238
rect 30156 4228 30212 4284
rect 29932 4226 30212 4228
rect 29932 4174 29934 4226
rect 29986 4174 30212 4226
rect 29932 4172 30212 4174
rect 29932 4162 29988 4172
rect 29596 3554 29876 3556
rect 29596 3502 29598 3554
rect 29650 3502 29876 3554
rect 29596 3500 29876 3502
rect 29372 3266 29428 3276
rect 29596 2772 29652 3500
rect 29484 2716 29652 2772
rect 29484 800 29540 2716
rect 30156 800 30212 4172
rect 30268 3330 30324 28814
rect 30380 28644 30436 28654
rect 30492 28644 30548 29374
rect 30436 28588 30548 28644
rect 30604 29428 30660 29438
rect 30604 28644 30660 29372
rect 31276 29316 31332 30046
rect 31612 30100 31668 30110
rect 31612 30006 31668 30044
rect 32060 29988 32116 30270
rect 30940 29314 31332 29316
rect 30940 29262 31278 29314
rect 31330 29262 31332 29314
rect 30940 29260 31332 29262
rect 30940 28866 30996 29260
rect 31276 29250 31332 29260
rect 31724 29932 32116 29988
rect 30940 28814 30942 28866
rect 30994 28814 30996 28866
rect 30940 28802 30996 28814
rect 30828 28644 30884 28654
rect 30604 28642 30884 28644
rect 30604 28590 30830 28642
rect 30882 28590 30884 28642
rect 30604 28588 30884 28590
rect 30380 28550 30436 28588
rect 30604 4564 30660 28588
rect 30828 28578 30884 28588
rect 31724 8428 31780 29932
rect 32172 8428 32228 31892
rect 32620 31668 32676 31678
rect 32284 31108 32340 31118
rect 32284 31014 32340 31052
rect 32620 20188 32676 31612
rect 32956 31556 33012 31566
rect 32956 31462 33012 31500
rect 32732 30996 32788 31006
rect 32732 30902 32788 30940
rect 32620 20132 32900 20188
rect 31164 8372 31780 8428
rect 32060 8372 32228 8428
rect 30828 4898 30884 4910
rect 30828 4846 30830 4898
rect 30882 4846 30884 4898
rect 30716 4564 30772 4574
rect 30604 4562 30772 4564
rect 30604 4510 30718 4562
rect 30770 4510 30772 4562
rect 30604 4508 30772 4510
rect 30716 4498 30772 4508
rect 30380 4340 30436 4350
rect 30380 4246 30436 4284
rect 30604 3444 30660 3454
rect 30828 3444 30884 4846
rect 30604 3442 30884 3444
rect 30604 3390 30606 3442
rect 30658 3390 30884 3442
rect 30604 3388 30884 3390
rect 30604 3378 30660 3388
rect 30268 3278 30270 3330
rect 30322 3278 30324 3330
rect 30268 3266 30324 3278
rect 30828 800 30884 3388
rect 31164 3330 31220 8372
rect 31948 4340 32004 4350
rect 31164 3278 31166 3330
rect 31218 3278 31220 3330
rect 31164 3266 31220 3278
rect 31500 4226 31556 4238
rect 31500 4174 31502 4226
rect 31554 4174 31556 4226
rect 31500 3442 31556 4174
rect 31500 3390 31502 3442
rect 31554 3390 31556 3442
rect 31500 800 31556 3390
rect 31948 4226 32004 4284
rect 31948 4174 31950 4226
rect 32002 4174 32004 4226
rect 31948 2884 32004 4174
rect 32060 3330 32116 8372
rect 32732 4900 32788 4910
rect 32620 4898 32788 4900
rect 32620 4846 32734 4898
rect 32786 4846 32788 4898
rect 32620 4844 32788 4846
rect 32396 4340 32452 4350
rect 32396 4246 32452 4284
rect 32060 3278 32062 3330
rect 32114 3278 32116 3330
rect 32060 3266 32116 3278
rect 32396 3442 32452 3454
rect 32396 3390 32398 3442
rect 32450 3390 32452 3442
rect 31948 2828 32228 2884
rect 32172 800 32228 2828
rect 32396 2772 32452 3390
rect 32620 2772 32676 4844
rect 32732 4834 32788 4844
rect 32732 4564 32788 4574
rect 32844 4564 32900 20132
rect 32732 4562 32900 4564
rect 32732 4510 32734 4562
rect 32786 4510 32900 4562
rect 32732 4508 32900 4510
rect 32732 4498 32788 4508
rect 33292 3330 33348 31892
rect 33404 31890 33460 32508
rect 33628 32564 33684 32574
rect 33628 32470 33684 32508
rect 33404 31838 33406 31890
rect 33458 31838 33460 31890
rect 33404 31826 33460 31838
rect 33852 31668 33908 31678
rect 33852 31574 33908 31612
rect 34860 8428 34916 33070
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 34524 8372 34916 8428
rect 33628 4226 33684 4238
rect 33628 4174 33630 4226
rect 33682 4174 33684 4226
rect 33628 3444 33684 4174
rect 33292 3278 33294 3330
rect 33346 3278 33348 3330
rect 33292 3266 33348 3278
rect 33516 3442 33684 3444
rect 33516 3390 33630 3442
rect 33682 3390 33684 3442
rect 33516 3388 33684 3390
rect 32396 2716 32900 2772
rect 32844 800 32900 2716
rect 33516 800 33572 3388
rect 33628 3378 33684 3388
rect 34188 4226 34244 4238
rect 34188 4174 34190 4226
rect 34242 4174 34244 4226
rect 34188 3442 34244 4174
rect 34188 3390 34190 3442
rect 34242 3390 34244 3442
rect 34188 800 34244 3390
rect 34524 3330 34580 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35420 4564 35476 4574
rect 35532 4564 35588 33964
rect 35644 33954 35700 33964
rect 36092 34018 36148 34862
rect 36764 35698 36820 35756
rect 36988 35812 37044 35822
rect 36988 35718 37044 35756
rect 36764 35646 36766 35698
rect 36818 35646 36820 35698
rect 36316 34804 36372 34814
rect 36316 34710 36372 34748
rect 36092 33966 36094 34018
rect 36146 33966 36148 34018
rect 35980 33906 36036 33918
rect 35980 33854 35982 33906
rect 36034 33854 36036 33906
rect 35420 4562 35588 4564
rect 35420 4510 35422 4562
rect 35474 4510 35588 4562
rect 35420 4508 35588 4510
rect 35644 4898 35700 4910
rect 35644 4846 35646 4898
rect 35698 4846 35700 4898
rect 35420 4498 35476 4508
rect 35084 4338 35140 4350
rect 35084 4286 35086 4338
rect 35138 4286 35140 4338
rect 34636 4228 34692 4238
rect 35084 4228 35140 4286
rect 34636 4226 35140 4228
rect 34636 4174 34638 4226
rect 34690 4174 35140 4226
rect 34636 4172 35140 4174
rect 34636 4162 34692 4172
rect 34524 3278 34526 3330
rect 34578 3278 34580 3330
rect 34524 3266 34580 3278
rect 34860 800 34916 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35420 3444 35476 3454
rect 35644 3444 35700 4846
rect 35420 3442 35700 3444
rect 35420 3390 35422 3442
rect 35474 3390 35700 3442
rect 35420 3388 35700 3390
rect 35420 3378 35476 3388
rect 35084 3332 35140 3342
rect 35084 3238 35140 3276
rect 35532 800 35588 3388
rect 35980 3330 36036 33854
rect 35980 3278 35982 3330
rect 36034 3278 36036 3330
rect 35980 3266 36036 3278
rect 36092 3332 36148 33966
rect 36764 34690 36820 35646
rect 36764 34638 36766 34690
rect 36818 34638 36820 34690
rect 36204 33908 36260 33918
rect 36764 33908 36820 34638
rect 36204 33906 36820 33908
rect 36204 33854 36206 33906
rect 36258 33854 36820 33906
rect 36204 33852 36820 33854
rect 36204 33842 36260 33852
rect 37100 4338 37156 4350
rect 37100 4286 37102 4338
rect 37154 4286 37156 4338
rect 36092 3266 36148 3276
rect 36204 4226 36260 4238
rect 36204 4174 36206 4226
rect 36258 4174 36260 4226
rect 36204 3554 36260 4174
rect 36652 4228 36708 4238
rect 37100 4228 37156 4286
rect 36652 4226 37156 4228
rect 36652 4174 36654 4226
rect 36706 4174 37156 4226
rect 36652 4172 37156 4174
rect 36652 4162 36708 4172
rect 36204 3502 36206 3554
rect 36258 3502 36260 3554
rect 36204 800 36260 3502
rect 36876 800 36932 4172
rect 37212 3330 37268 37100
rect 37996 37266 38052 37278
rect 37996 37214 37998 37266
rect 38050 37214 38052 37266
rect 37996 37156 38052 37214
rect 37996 37090 38052 37100
rect 38332 37156 38388 37166
rect 38668 37156 38724 37884
rect 39004 37828 39060 37838
rect 39004 37734 39060 37772
rect 38780 37156 38836 37166
rect 38332 36594 38388 37100
rect 38332 36542 38334 36594
rect 38386 36542 38388 36594
rect 38332 36530 38388 36542
rect 38444 37154 38836 37156
rect 38444 37102 38782 37154
rect 38834 37102 38836 37154
rect 38444 37100 38836 37102
rect 37548 36372 37604 36382
rect 37436 35700 37492 35710
rect 37436 35606 37492 35644
rect 37548 31948 37604 36316
rect 37884 36260 37940 36270
rect 37884 36166 37940 36204
rect 37436 31892 37604 31948
rect 37436 4562 37492 31892
rect 37436 4510 37438 4562
rect 37490 4510 37492 4562
rect 37436 4498 37492 4510
rect 37772 4898 37828 4910
rect 37772 4846 37774 4898
rect 37826 4846 37828 4898
rect 37212 3278 37214 3330
rect 37266 3278 37268 3330
rect 37212 3266 37268 3278
rect 37548 3444 37604 3454
rect 37772 3444 37828 4846
rect 37548 3442 37828 3444
rect 37548 3390 37550 3442
rect 37602 3390 37828 3442
rect 37548 3388 37828 3390
rect 38220 4226 38276 4238
rect 38220 4174 38222 4226
rect 38274 4174 38276 4226
rect 38220 3554 38276 4174
rect 38220 3502 38222 3554
rect 38274 3502 38276 3554
rect 37548 800 37604 3388
rect 38220 800 38276 3502
rect 38444 3330 38500 37100
rect 38780 37090 38836 37100
rect 38780 36372 38836 36382
rect 38780 36278 38836 36316
rect 39116 15148 39172 39452
rect 39676 39508 39732 39518
rect 39676 39414 39732 39452
rect 39788 38948 39844 38958
rect 39788 38854 39844 38892
rect 39564 38836 39620 38846
rect 39452 37940 39508 37950
rect 39452 37846 39508 37884
rect 39564 31948 39620 38780
rect 39004 15092 39172 15148
rect 39452 31892 39620 31948
rect 39900 38724 39956 40348
rect 40572 40404 40628 40414
rect 40572 40310 40628 40348
rect 41580 40404 41636 40414
rect 40572 39506 40628 39518
rect 40572 39454 40574 39506
rect 40626 39454 40628 39506
rect 40012 39396 40068 39406
rect 40012 39302 40068 39340
rect 40236 38724 40292 38734
rect 40572 38724 40628 39454
rect 40908 39508 40964 39518
rect 40908 39414 40964 39452
rect 41356 39396 41412 39406
rect 41580 39396 41636 40348
rect 41356 39394 41636 39396
rect 41356 39342 41358 39394
rect 41410 39342 41636 39394
rect 41356 39340 41636 39342
rect 40684 38836 40740 38846
rect 40684 38742 40740 38780
rect 39900 38722 40628 38724
rect 39900 38670 40238 38722
rect 40290 38670 40628 38722
rect 39900 38668 40628 38670
rect 38668 4340 38724 4350
rect 38668 4246 38724 4284
rect 38892 4340 38948 4350
rect 38444 3278 38446 3330
rect 38498 3278 38500 3330
rect 38444 3266 38500 3278
rect 38892 800 38948 4284
rect 39004 3330 39060 15092
rect 39452 4562 39508 31892
rect 39900 20188 39956 38668
rect 40236 38658 40292 38668
rect 41356 31948 41412 39340
rect 41356 31892 41972 31948
rect 39900 20132 40068 20188
rect 39452 4510 39454 4562
rect 39506 4510 39508 4562
rect 39452 4498 39508 4510
rect 39116 4340 39172 4350
rect 39116 4246 39172 4284
rect 39900 4228 39956 4238
rect 39564 4226 39956 4228
rect 39564 4174 39902 4226
rect 39954 4174 39956 4226
rect 39564 4172 39956 4174
rect 39340 3556 39396 3566
rect 39564 3556 39620 4172
rect 39900 4162 39956 4172
rect 39340 3554 39620 3556
rect 39340 3502 39342 3554
rect 39394 3502 39620 3554
rect 39340 3500 39620 3502
rect 39340 3490 39396 3500
rect 39004 3278 39006 3330
rect 39058 3278 39060 3330
rect 39004 3266 39060 3278
rect 39564 800 39620 3500
rect 39900 3332 39956 3342
rect 40012 3332 40068 20132
rect 41916 4562 41972 31892
rect 41916 4510 41918 4562
rect 41970 4510 41972 4562
rect 41916 4498 41972 4510
rect 40908 4340 40964 4350
rect 40348 4226 40404 4238
rect 40348 4174 40350 4226
rect 40402 4174 40404 4226
rect 39900 3330 40068 3332
rect 39900 3278 39902 3330
rect 39954 3278 40068 3330
rect 39900 3276 40068 3278
rect 40236 3556 40292 3566
rect 40348 3556 40404 4174
rect 40236 3554 40404 3556
rect 40236 3502 40238 3554
rect 40290 3502 40404 3554
rect 40236 3500 40404 3502
rect 40908 4226 40964 4284
rect 41580 4340 41636 4350
rect 41580 4246 41636 4284
rect 40908 4174 40910 4226
rect 40962 4174 40964 4226
rect 39900 3266 39956 3276
rect 40236 800 40292 3500
rect 40908 800 40964 4174
rect 41356 3442 41412 3454
rect 41356 3390 41358 3442
rect 41410 3390 41412 3442
rect 41356 3388 41412 3390
rect 41804 3442 41860 3454
rect 41804 3390 41806 3442
rect 41858 3390 41860 3442
rect 41804 3388 41860 3390
rect 41356 3332 41860 3388
rect 41580 800 41636 3332
rect 42140 3330 42196 40908
rect 42812 40964 42868 40974
rect 42812 40870 42868 40908
rect 42364 40404 42420 40414
rect 42364 40310 42420 40348
rect 42924 31948 42980 41804
rect 43036 40964 43092 42030
rect 43484 41860 43540 41870
rect 43484 41766 43540 41804
rect 43932 41860 43988 41870
rect 43932 41766 43988 41804
rect 43036 40898 43092 40908
rect 42924 31892 43092 31948
rect 42476 4228 42532 4238
rect 42476 4226 42756 4228
rect 42476 4174 42478 4226
rect 42530 4174 42756 4226
rect 42476 4172 42756 4174
rect 42476 4162 42532 4172
rect 42700 3554 42756 4172
rect 42700 3502 42702 3554
rect 42754 3502 42756 3554
rect 42700 3388 42756 3502
rect 42140 3278 42142 3330
rect 42194 3278 42196 3330
rect 42140 3266 42196 3278
rect 42252 3332 42756 3388
rect 42924 4226 42980 4238
rect 42924 4174 42926 4226
rect 42978 4174 42980 4226
rect 42924 3556 42980 4174
rect 42252 800 42308 3332
rect 42924 800 42980 3500
rect 43036 3330 43092 31892
rect 43820 4338 43876 4350
rect 43820 4286 43822 4338
rect 43874 4286 43876 4338
rect 43372 4228 43428 4238
rect 43820 4228 43876 4286
rect 43372 4226 43876 4228
rect 43372 4174 43374 4226
rect 43426 4174 43876 4226
rect 43372 4172 43876 4174
rect 43372 4162 43428 4172
rect 43036 3278 43038 3330
rect 43090 3278 43092 3330
rect 43036 3266 43092 3278
rect 43484 3220 43540 4172
rect 43596 3556 43652 3566
rect 43596 3462 43652 3500
rect 44044 3388 44100 42476
rect 44156 42466 44212 42476
rect 44268 31948 44324 43372
rect 44828 43428 44884 43438
rect 44828 43334 44884 43372
rect 45276 43426 45332 44156
rect 45500 44212 45556 44222
rect 45500 44118 45556 44156
rect 45836 44212 45892 44222
rect 45836 44118 45892 44156
rect 46396 43708 46452 44270
rect 46732 44100 46788 44110
rect 46732 44006 46788 44044
rect 46172 43652 46452 43708
rect 45276 43374 45278 43426
rect 45330 43374 45332 43426
rect 44156 31892 44324 31948
rect 44156 4562 44212 31892
rect 44156 4510 44158 4562
rect 44210 4510 44212 4562
rect 44156 4498 44212 4510
rect 44716 4228 44772 4238
rect 44716 4226 44996 4228
rect 44716 4174 44718 4226
rect 44770 4174 44996 4226
rect 44716 4172 44996 4174
rect 44716 4162 44772 4172
rect 43932 3332 44100 3388
rect 44268 3556 44324 3566
rect 43932 3330 43988 3332
rect 43932 3278 43934 3330
rect 43986 3278 43988 3330
rect 43932 3266 43988 3278
rect 43484 3164 43652 3220
rect 43596 800 43652 3164
rect 44268 800 44324 3500
rect 44940 3556 44996 4172
rect 44940 3424 44996 3500
rect 45052 3444 45108 3454
rect 45052 2884 45108 3388
rect 45276 3330 45332 43374
rect 46060 43428 46116 43438
rect 46172 43428 46228 43652
rect 46060 43426 46228 43428
rect 46060 43374 46062 43426
rect 46114 43374 46228 43426
rect 46060 43372 46228 43374
rect 46060 43362 46116 43372
rect 46060 4340 46116 4350
rect 45612 4226 45668 4238
rect 45612 4174 45614 4226
rect 45666 4174 45668 4226
rect 45612 3556 45668 4174
rect 46060 4226 46116 4284
rect 46060 4174 46062 4226
rect 46114 4174 46116 4226
rect 45836 3556 45892 3566
rect 45612 3554 45892 3556
rect 45612 3502 45838 3554
rect 45890 3502 45892 3554
rect 45612 3500 45892 3502
rect 45612 3444 45668 3500
rect 45836 3490 45892 3500
rect 45948 3444 46004 3454
rect 45612 3378 45668 3388
rect 45276 3278 45278 3330
rect 45330 3278 45332 3330
rect 45276 3266 45332 3278
rect 45724 3332 46004 3388
rect 44940 2828 45108 2884
rect 44940 800 44996 2828
rect 45724 2772 45780 3332
rect 46060 2884 46116 4174
rect 46172 3330 46228 43372
rect 46844 4562 46900 45724
rect 47180 45780 47236 45790
rect 47180 45686 47236 45724
rect 46844 4510 46846 4562
rect 46898 4510 46900 4562
rect 46844 4498 46900 4510
rect 46956 45108 47012 45118
rect 46956 44996 47012 45052
rect 47404 44996 47460 45006
rect 46956 44994 47460 44996
rect 46956 44942 46958 44994
rect 47010 44942 47406 44994
rect 47458 44942 47460 44994
rect 46956 44940 47460 44942
rect 46508 4340 46564 4350
rect 46956 4340 47012 44940
rect 47404 44930 47460 44940
rect 47628 15148 47684 46508
rect 47740 45892 47796 45902
rect 47740 45798 47796 45836
rect 48076 45892 48132 45902
rect 48076 45798 48132 45836
rect 46508 4246 46564 4284
rect 46732 4284 47012 4340
rect 47516 15092 47684 15148
rect 46172 3278 46174 3330
rect 46226 3278 46228 3330
rect 46172 3266 46228 3278
rect 46732 3330 46788 4284
rect 47292 4228 47348 4238
rect 47068 4226 47348 4228
rect 47068 4174 47294 4226
rect 47346 4174 47348 4226
rect 47068 4172 47348 4174
rect 46732 3278 46734 3330
rect 46786 3278 46788 3330
rect 46732 3266 46788 3278
rect 46956 3556 47012 3566
rect 46060 2828 46340 2884
rect 45612 2716 45780 2772
rect 45612 800 45668 2716
rect 46284 800 46340 2828
rect 46956 800 47012 3500
rect 47068 3554 47124 4172
rect 47292 4162 47348 4172
rect 47068 3502 47070 3554
rect 47122 3502 47124 3554
rect 47068 3444 47124 3502
rect 47068 3378 47124 3388
rect 47516 3332 47572 15092
rect 47628 4900 47684 4910
rect 47628 4898 47908 4900
rect 47628 4846 47630 4898
rect 47682 4846 47908 4898
rect 47628 4844 47908 4846
rect 47628 4834 47684 4844
rect 47852 4450 47908 4844
rect 48188 4562 48244 47292
rect 48972 47348 49028 47358
rect 48972 47254 49028 47292
rect 48524 47236 48580 47246
rect 48524 47142 48580 47180
rect 48300 46564 48356 46574
rect 48300 46470 48356 46508
rect 49308 31948 49364 48750
rect 49420 48804 49476 48814
rect 49420 48710 49476 48748
rect 49532 48468 49588 49534
rect 49644 49138 49700 49644
rect 49756 49568 49812 49644
rect 49980 49252 50036 49758
rect 49980 49186 50036 49196
rect 50092 49698 50148 49710
rect 50092 49646 50094 49698
rect 50146 49646 50148 49698
rect 49644 49086 49646 49138
rect 49698 49086 49700 49138
rect 49644 49074 49700 49086
rect 49868 49028 49924 49038
rect 49868 48934 49924 48972
rect 49868 48804 49924 48814
rect 49756 48468 49812 48478
rect 49532 48466 49812 48468
rect 49532 48414 49758 48466
rect 49810 48414 49812 48466
rect 49532 48412 49812 48414
rect 49756 48402 49812 48412
rect 49868 48354 49924 48748
rect 49868 48302 49870 48354
rect 49922 48302 49924 48354
rect 49868 48290 49924 48302
rect 50092 31948 50148 49646
rect 50428 49588 50484 49980
rect 50876 49700 50932 50372
rect 51772 50372 51828 50382
rect 50876 49634 50932 49644
rect 50988 50148 51044 50158
rect 50988 50034 51044 50092
rect 50988 49982 50990 50034
rect 51042 49982 51044 50034
rect 50428 49522 50484 49532
rect 50988 49588 51044 49982
rect 51212 50036 51268 50046
rect 51212 49942 51268 49980
rect 50988 49522 51044 49532
rect 51100 49698 51156 49710
rect 51100 49646 51102 49698
rect 51154 49646 51156 49698
rect 50316 49476 50372 49486
rect 50316 48804 50372 49420
rect 50428 49028 50484 49038
rect 51100 49028 51156 49646
rect 51436 49700 51492 49710
rect 51436 49606 51492 49644
rect 51660 49588 51716 49598
rect 51660 49494 51716 49532
rect 51100 48972 51268 49028
rect 50428 48934 50484 48972
rect 50316 48466 50372 48748
rect 50540 48914 50596 48926
rect 50540 48862 50542 48914
rect 50594 48862 50596 48914
rect 50540 48804 50596 48862
rect 50540 48738 50596 48748
rect 51100 48804 51156 48814
rect 51100 48710 51156 48748
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50316 48414 50318 48466
rect 50370 48414 50372 48466
rect 50316 48402 50372 48414
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 51212 31948 51268 48972
rect 49196 31892 49364 31948
rect 49980 31892 50148 31948
rect 51100 31892 51268 31948
rect 49196 5236 49252 31892
rect 49308 5236 49364 5246
rect 49196 5234 49364 5236
rect 49196 5182 49310 5234
rect 49362 5182 49364 5234
rect 49196 5180 49364 5182
rect 48188 4510 48190 4562
rect 48242 4510 48244 4562
rect 48188 4498 48244 4510
rect 47852 4398 47854 4450
rect 47906 4398 47908 4450
rect 47628 3332 47684 3342
rect 47516 3330 47684 3332
rect 47516 3278 47630 3330
rect 47682 3278 47684 3330
rect 47516 3276 47684 3278
rect 47628 3266 47684 3276
rect 47852 3108 47908 4398
rect 49308 4340 49364 5180
rect 49980 5236 50036 31892
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50316 5908 50372 5918
rect 50316 5236 50372 5852
rect 49980 5104 50036 5180
rect 50092 5234 50372 5236
rect 50092 5182 50318 5234
rect 50370 5182 50372 5234
rect 50092 5180 50372 5182
rect 49532 4340 49588 4350
rect 49308 4338 49588 4340
rect 49308 4286 49534 4338
rect 49586 4286 49588 4338
rect 49308 4284 49588 4286
rect 49532 4274 49588 4284
rect 47964 4228 48020 4238
rect 47964 3556 48020 4172
rect 48636 4228 48692 4238
rect 48636 4134 48692 4172
rect 48972 4228 49028 4238
rect 47964 3424 48020 3500
rect 48300 3444 48356 3454
rect 47628 3052 47908 3108
rect 47628 800 47684 3052
rect 48300 800 48356 3388
rect 48972 800 49028 4172
rect 50092 3554 50148 5180
rect 50316 5170 50372 5180
rect 50876 5236 50932 5246
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 50204 4228 50260 4238
rect 50204 4134 50260 4172
rect 50092 3502 50094 3554
rect 50146 3502 50148 3554
rect 50092 3490 50148 3502
rect 50316 3556 50372 3566
rect 49196 3444 49252 3482
rect 49196 3378 49252 3388
rect 49644 3444 49700 3454
rect 49644 800 49700 3388
rect 50316 800 50372 3500
rect 50876 3554 50932 5180
rect 51100 5234 51156 31892
rect 51100 5182 51102 5234
rect 51154 5182 51156 5234
rect 51100 4340 51156 5182
rect 51772 5236 51828 50316
rect 51996 5236 52052 51214
rect 52220 49812 52276 51660
rect 52332 51378 52388 52220
rect 52444 52210 52500 52220
rect 52556 52276 52612 52286
rect 52332 51326 52334 51378
rect 52386 51326 52388 51378
rect 52332 51314 52388 51326
rect 52556 51378 52612 52220
rect 52556 51326 52558 51378
rect 52610 51326 52612 51378
rect 52556 51314 52612 51326
rect 52668 51492 52724 51502
rect 52332 50596 52388 50606
rect 52332 50502 52388 50540
rect 52332 49924 52388 49934
rect 52668 49924 52724 51436
rect 52332 49922 52724 49924
rect 52332 49870 52334 49922
rect 52386 49870 52724 49922
rect 52332 49868 52724 49870
rect 52780 49924 52836 52782
rect 53116 52836 53172 52846
rect 53116 52742 53172 52780
rect 53228 51940 53284 53116
rect 53900 52946 53956 53452
rect 54460 53172 54516 53182
rect 54572 53172 54628 54124
rect 54684 53732 54740 53742
rect 54684 53638 54740 53676
rect 54908 53732 54964 54796
rect 55020 54516 55076 54526
rect 55244 54516 55300 55022
rect 55356 55076 55412 55086
rect 55356 54982 55412 55020
rect 55020 54422 55076 54460
rect 55132 54460 55300 54516
rect 55132 54180 55188 54460
rect 55356 54404 55412 54414
rect 55244 54292 55300 54302
rect 55244 54198 55300 54236
rect 55132 54114 55188 54124
rect 54908 53600 54964 53676
rect 54796 53506 54852 53518
rect 54796 53454 54798 53506
rect 54850 53454 54852 53506
rect 54572 53116 54740 53172
rect 54348 53060 54404 53070
rect 54460 53060 54516 53116
rect 54460 53004 54628 53060
rect 54348 52966 54404 53004
rect 53900 52894 53902 52946
rect 53954 52894 53956 52946
rect 53900 52882 53956 52894
rect 54572 52946 54628 53004
rect 54572 52894 54574 52946
rect 54626 52894 54628 52946
rect 54572 52882 54628 52894
rect 54124 52836 54180 52846
rect 54124 52742 54180 52780
rect 54460 52834 54516 52846
rect 54460 52782 54462 52834
rect 54514 52782 54516 52834
rect 53340 52724 53396 52734
rect 53340 52630 53396 52668
rect 53228 51604 53284 51884
rect 53340 51604 53396 51614
rect 53228 51602 53396 51604
rect 53228 51550 53342 51602
rect 53394 51550 53396 51602
rect 53228 51548 53396 51550
rect 53340 51538 53396 51548
rect 53676 51604 53732 51614
rect 53676 51490 53732 51548
rect 53676 51438 53678 51490
rect 53730 51438 53732 51490
rect 53676 50594 53732 51438
rect 53676 50542 53678 50594
rect 53730 50542 53732 50594
rect 53676 50530 53732 50542
rect 53452 50370 53508 50382
rect 53452 50318 53454 50370
rect 53506 50318 53508 50370
rect 53452 50148 53508 50318
rect 53452 50082 53508 50092
rect 52780 49868 52948 49924
rect 52332 49858 52388 49868
rect 52108 49756 52276 49812
rect 52108 43708 52164 49756
rect 52668 49700 52724 49868
rect 52780 49700 52836 49710
rect 52668 49698 52836 49700
rect 52668 49646 52782 49698
rect 52834 49646 52836 49698
rect 52668 49644 52836 49646
rect 52780 49634 52836 49644
rect 52220 49588 52276 49598
rect 52220 49494 52276 49532
rect 52108 43652 52724 43708
rect 52668 6132 52724 43652
rect 52892 31948 52948 49868
rect 52668 6066 52724 6076
rect 52780 31892 52948 31948
rect 52780 5572 52836 31892
rect 54460 20188 54516 52782
rect 54348 20132 54516 20188
rect 53564 17442 53620 17454
rect 53564 17390 53566 17442
rect 53618 17390 53620 17442
rect 53564 17108 53620 17390
rect 54012 17444 54068 17454
rect 54012 17350 54068 17388
rect 53564 17042 53620 17052
rect 53900 15316 53956 15326
rect 53900 14642 53956 15260
rect 53900 14590 53902 14642
rect 53954 14590 53956 14642
rect 53900 14578 53956 14590
rect 53452 14420 53508 14430
rect 53452 14326 53508 14364
rect 54348 14308 54404 20132
rect 54572 18452 54628 18462
rect 54572 18340 54628 18396
rect 54460 18338 54628 18340
rect 54460 18286 54574 18338
rect 54626 18286 54628 18338
rect 54460 18284 54628 18286
rect 54460 16884 54516 18284
rect 54572 18274 54628 18284
rect 54460 16790 54516 16828
rect 54572 17220 54628 17230
rect 54572 14756 54628 17164
rect 54460 14700 54628 14756
rect 54460 14420 54516 14700
rect 54684 14532 54740 53116
rect 54796 43708 54852 53454
rect 54796 43652 55188 43708
rect 54796 18564 54852 18574
rect 54796 17554 54852 18508
rect 54796 17502 54798 17554
rect 54850 17502 54852 17554
rect 54796 16212 54852 17502
rect 55020 18340 55076 18350
rect 55020 17442 55076 18284
rect 55020 17390 55022 17442
rect 55074 17390 55076 17442
rect 55020 17108 55076 17390
rect 55132 17220 55188 43652
rect 55132 17154 55188 17164
rect 55244 17442 55300 17454
rect 55244 17390 55246 17442
rect 55298 17390 55300 17442
rect 55020 17042 55076 17052
rect 55244 16884 55300 17390
rect 55244 16818 55300 16828
rect 54796 16156 55188 16212
rect 54796 15316 54852 15326
rect 54796 14754 54852 15260
rect 55020 15316 55076 15326
rect 55020 15222 55076 15260
rect 54796 14702 54798 14754
rect 54850 14702 54852 14754
rect 54796 14690 54852 14702
rect 54684 14476 54852 14532
rect 54460 14364 54740 14420
rect 54348 14252 54516 14308
rect 54348 13634 54404 13646
rect 54348 13582 54350 13634
rect 54402 13582 54404 13634
rect 54348 13524 54404 13582
rect 54348 13458 54404 13468
rect 54236 6132 54292 6142
rect 54236 6038 54292 6076
rect 52780 5516 53508 5572
rect 52332 5348 52388 5358
rect 52332 5236 52388 5292
rect 51996 5234 52388 5236
rect 51996 5182 52334 5234
rect 52386 5182 52388 5234
rect 51996 5180 52388 5182
rect 51772 5104 51828 5180
rect 52332 5170 52388 5180
rect 52668 5236 52724 5246
rect 51324 4340 51380 4350
rect 51100 4338 51380 4340
rect 51100 4286 51326 4338
rect 51378 4286 51380 4338
rect 51100 4284 51380 4286
rect 51324 4274 51380 4284
rect 52108 4226 52164 4238
rect 52108 4174 52110 4226
rect 52162 4174 52164 4226
rect 51660 3780 51716 3790
rect 50876 3502 50878 3554
rect 50930 3502 50932 3554
rect 50876 3490 50932 3502
rect 50988 3668 51044 3678
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 50988 800 51044 3612
rect 51548 3444 51604 3454
rect 51548 3350 51604 3388
rect 51660 800 51716 3724
rect 52108 3556 52164 4174
rect 52668 3556 52724 5180
rect 52780 5234 52836 5516
rect 52780 5182 52782 5234
rect 52834 5182 52836 5234
rect 52780 5170 52836 5182
rect 53116 5348 53172 5358
rect 53116 4338 53172 5292
rect 53452 5122 53508 5516
rect 53452 5070 53454 5122
rect 53506 5070 53508 5122
rect 53452 5058 53508 5070
rect 53564 5236 53620 5246
rect 53116 4286 53118 4338
rect 53170 4286 53172 4338
rect 53116 4274 53172 4286
rect 53452 3668 53508 3678
rect 53452 3574 53508 3612
rect 52780 3556 52836 3566
rect 52668 3554 52836 3556
rect 52668 3502 52782 3554
rect 52834 3502 52836 3554
rect 52668 3500 52836 3502
rect 52108 3490 52164 3500
rect 52780 3490 52836 3500
rect 52332 3444 52388 3454
rect 52332 800 52388 3388
rect 53564 2660 53620 5180
rect 54124 5236 54180 5246
rect 54124 5142 54180 5180
rect 54460 4340 54516 14252
rect 54572 14196 54628 14206
rect 54572 6244 54628 14140
rect 54684 8428 54740 14364
rect 54796 14308 54852 14476
rect 55020 14530 55076 14542
rect 55020 14478 55022 14530
rect 55074 14478 55076 14530
rect 55020 14420 55076 14478
rect 55020 14354 55076 14364
rect 54796 14242 54852 14252
rect 55132 14306 55188 16156
rect 55132 14254 55134 14306
rect 55186 14254 55188 14306
rect 55132 14242 55188 14254
rect 55244 14530 55300 14542
rect 55244 14478 55246 14530
rect 55298 14478 55300 14530
rect 55244 13746 55300 14478
rect 55244 13694 55246 13746
rect 55298 13694 55300 13746
rect 54908 13524 54964 13534
rect 54908 13074 54964 13468
rect 55244 13524 55300 13694
rect 55244 13458 55300 13468
rect 54908 13022 54910 13074
rect 54962 13022 54964 13074
rect 54908 13010 54964 13022
rect 55356 8428 55412 54348
rect 55468 53956 55524 55918
rect 55580 55412 55636 55422
rect 55692 55412 55748 56030
rect 56028 56082 56084 56364
rect 56588 56306 56644 56364
rect 56588 56254 56590 56306
rect 56642 56254 56644 56306
rect 56588 56242 56644 56254
rect 56812 56308 56868 56590
rect 56812 56242 56868 56252
rect 56028 56030 56030 56082
rect 56082 56030 56084 56082
rect 56028 56018 56084 56030
rect 56252 56196 56308 56206
rect 55580 55410 55748 55412
rect 55580 55358 55582 55410
rect 55634 55358 55748 55410
rect 55580 55356 55748 55358
rect 55580 55188 55636 55356
rect 55580 54516 55636 55132
rect 55804 55298 55860 55310
rect 55804 55246 55806 55298
rect 55858 55246 55860 55298
rect 55804 54964 55860 55246
rect 56252 55076 56308 56140
rect 56700 55972 56756 55982
rect 56700 55878 56756 55916
rect 56924 55300 56980 55310
rect 56924 55186 56980 55244
rect 56924 55134 56926 55186
rect 56978 55134 56980 55186
rect 56924 55076 56980 55134
rect 57260 55188 57316 55198
rect 57260 55094 57316 55132
rect 55804 54898 55860 54908
rect 55916 55074 56308 55076
rect 55916 55022 56254 55074
rect 56306 55022 56308 55074
rect 55916 55020 56308 55022
rect 55916 54626 55972 55020
rect 56252 55010 56308 55020
rect 56700 55020 56924 55076
rect 56476 54964 56532 54974
rect 56476 54738 56532 54908
rect 56476 54686 56478 54738
rect 56530 54686 56532 54738
rect 56476 54674 56532 54686
rect 56588 54852 56644 54862
rect 55916 54574 55918 54626
rect 55970 54574 55972 54626
rect 55916 54562 55972 54574
rect 56588 54626 56644 54796
rect 56588 54574 56590 54626
rect 56642 54574 56644 54626
rect 56588 54562 56644 54574
rect 55580 54450 55636 54460
rect 55804 54292 55860 54302
rect 55804 54198 55860 54236
rect 55468 53900 56532 53956
rect 55580 53732 55636 53742
rect 55580 53618 55636 53676
rect 55916 53732 55972 53742
rect 55916 53638 55972 53676
rect 56140 53732 56196 53742
rect 55580 53566 55582 53618
rect 55634 53566 55636 53618
rect 55580 53554 55636 53566
rect 56028 52948 56084 52958
rect 56028 52050 56084 52892
rect 56028 51998 56030 52050
rect 56082 51998 56084 52050
rect 56028 51986 56084 51998
rect 56140 51604 56196 53676
rect 56140 51472 56196 51548
rect 56252 52164 56308 52174
rect 55692 51380 55748 51390
rect 55580 51268 55636 51278
rect 55692 51268 55748 51324
rect 55580 51266 55748 51268
rect 55580 51214 55582 51266
rect 55634 51214 55748 51266
rect 55580 51212 55748 51214
rect 55580 51202 55636 51212
rect 55580 18564 55636 18574
rect 55580 18470 55636 18508
rect 55580 17780 55636 17790
rect 55692 17780 55748 51212
rect 56252 18674 56308 52108
rect 56364 51380 56420 51390
rect 56364 51286 56420 51324
rect 56252 18622 56254 18674
rect 56306 18622 56308 18674
rect 56252 18610 56308 18622
rect 55804 18450 55860 18462
rect 55804 18398 55806 18450
rect 55858 18398 55860 18450
rect 55804 18340 55860 18398
rect 56028 18452 56084 18462
rect 56028 18358 56084 18396
rect 56252 18450 56308 18462
rect 56252 18398 56254 18450
rect 56306 18398 56308 18450
rect 55804 18274 55860 18284
rect 56140 17892 56196 17902
rect 56252 17892 56308 18398
rect 56140 17890 56308 17892
rect 56140 17838 56142 17890
rect 56194 17838 56308 17890
rect 56140 17836 56308 17838
rect 56140 17826 56196 17836
rect 55580 17778 55748 17780
rect 55580 17726 55582 17778
rect 55634 17726 55748 17778
rect 55580 17724 55748 17726
rect 55580 17714 55636 17724
rect 55468 17554 55524 17566
rect 55468 17502 55470 17554
rect 55522 17502 55524 17554
rect 55468 17444 55524 17502
rect 55468 13748 55524 17388
rect 56028 17554 56084 17566
rect 56028 17502 56030 17554
rect 56082 17502 56084 17554
rect 56028 17444 56084 17502
rect 56028 17378 56084 17388
rect 55916 15428 55972 15438
rect 55916 15334 55972 15372
rect 55580 15316 55636 15326
rect 55580 15222 55636 15260
rect 56140 15204 56196 15214
rect 55916 14532 55972 14542
rect 55916 14438 55972 14476
rect 56140 14418 56196 15148
rect 56140 14366 56142 14418
rect 56194 14366 56196 14418
rect 56140 14354 56196 14366
rect 55580 13860 55636 13870
rect 55580 13766 55636 13804
rect 55468 13682 55524 13692
rect 54684 8372 54964 8428
rect 54572 6178 54628 6188
rect 54460 4274 54516 4284
rect 54684 6132 54740 6142
rect 53004 2604 53620 2660
rect 53676 4228 53732 4238
rect 53004 800 53060 2604
rect 53676 800 53732 4172
rect 53788 4226 53844 4238
rect 53788 4174 53790 4226
rect 53842 4174 53844 4226
rect 53788 3780 53844 4174
rect 53788 3714 53844 3724
rect 54348 3668 54404 3678
rect 54348 800 54404 3612
rect 54684 3554 54740 6076
rect 54908 6132 54964 8372
rect 55244 8372 55412 8428
rect 54908 6066 54964 6076
rect 55020 6132 55076 6142
rect 55244 6132 55300 8372
rect 56476 6356 56532 53900
rect 56700 53620 56756 55020
rect 56924 55010 56980 55020
rect 56588 53564 56756 53620
rect 56924 54628 56980 54638
rect 56924 53730 56980 54572
rect 56924 53678 56926 53730
rect 56978 53678 56980 53730
rect 56588 52948 56644 53564
rect 56700 53060 56756 53070
rect 56924 53060 56980 53678
rect 57148 53954 57204 53966
rect 57148 53902 57150 53954
rect 57202 53902 57204 53954
rect 57148 53732 57204 53902
rect 57148 53666 57204 53676
rect 56700 53058 56980 53060
rect 56700 53006 56702 53058
rect 56754 53006 56980 53058
rect 56700 53004 56980 53006
rect 56700 52994 56756 53004
rect 56588 52882 56644 52892
rect 56588 52724 56644 52734
rect 56588 52630 56644 52668
rect 56812 52164 56868 52174
rect 56812 52070 56868 52108
rect 57260 52164 57316 52174
rect 57260 52070 57316 52108
rect 57148 51380 57204 51390
rect 57148 50706 57204 51324
rect 57148 50654 57150 50706
rect 57202 50654 57204 50706
rect 57148 50642 57204 50654
rect 57372 43708 57428 56924
rect 57820 56868 57876 56878
rect 57932 56868 57988 57932
rect 58044 57540 58100 57550
rect 58156 57540 58212 57550
rect 58044 57538 58156 57540
rect 58044 57486 58046 57538
rect 58098 57486 58156 57538
rect 58044 57484 58156 57486
rect 58044 57474 58100 57484
rect 57708 56866 57988 56868
rect 57708 56814 57822 56866
rect 57874 56814 57988 56866
rect 57708 56812 57988 56814
rect 58044 56980 58100 56990
rect 58044 56866 58100 56924
rect 58044 56814 58046 56866
rect 58098 56814 58100 56866
rect 57596 56196 57652 56206
rect 57708 56196 57764 56812
rect 57820 56802 57876 56812
rect 58044 56802 58100 56814
rect 58156 56866 58212 57484
rect 58268 57428 58324 57438
rect 58268 57334 58324 57372
rect 58156 56814 58158 56866
rect 58210 56814 58212 56866
rect 57932 56642 57988 56654
rect 57932 56590 57934 56642
rect 57986 56590 57988 56642
rect 57820 56308 57876 56318
rect 57820 56214 57876 56252
rect 57596 56194 57764 56196
rect 57596 56142 57598 56194
rect 57650 56142 57764 56194
rect 57596 56140 57764 56142
rect 57596 55522 57652 56140
rect 57596 55470 57598 55522
rect 57650 55470 57652 55522
rect 57596 55458 57652 55470
rect 57708 55970 57764 55982
rect 57708 55918 57710 55970
rect 57762 55918 57764 55970
rect 57708 55300 57764 55918
rect 57708 55234 57764 55244
rect 57820 55522 57876 55534
rect 57820 55470 57822 55522
rect 57874 55470 57876 55522
rect 57708 55076 57764 55086
rect 57708 54982 57764 55020
rect 57596 54852 57652 54862
rect 57484 54514 57540 54526
rect 57484 54462 57486 54514
rect 57538 54462 57540 54514
rect 57484 53954 57540 54462
rect 57484 53902 57486 53954
rect 57538 53902 57540 53954
rect 57484 53890 57540 53902
rect 57484 53732 57540 53742
rect 57596 53732 57652 54796
rect 57820 54738 57876 55470
rect 57820 54686 57822 54738
rect 57874 54686 57876 54738
rect 57820 54674 57876 54686
rect 57484 53730 57652 53732
rect 57484 53678 57486 53730
rect 57538 53678 57652 53730
rect 57484 53676 57652 53678
rect 57484 53666 57540 53676
rect 57820 53172 57876 53182
rect 57820 53078 57876 53116
rect 57484 52946 57540 52958
rect 57484 52894 57486 52946
rect 57538 52894 57540 52946
rect 57484 52164 57540 52894
rect 57484 52098 57540 52108
rect 57820 51604 57876 51614
rect 57820 51510 57876 51548
rect 57484 51380 57540 51390
rect 57484 51286 57540 51324
rect 57372 43652 57764 43708
rect 56588 17444 56644 17454
rect 56588 17350 56644 17388
rect 56588 14532 56644 14542
rect 56588 14438 56644 14476
rect 56700 13748 56756 13758
rect 56700 13654 56756 13692
rect 57484 13748 57540 13758
rect 57484 13654 57540 13692
rect 56476 6290 56532 6300
rect 57372 6244 57428 6254
rect 55020 6130 55300 6132
rect 55020 6078 55022 6130
rect 55074 6078 55300 6130
rect 55020 6076 55300 6078
rect 55020 6066 55076 6076
rect 54684 3502 54686 3554
rect 54738 3502 54740 3554
rect 54684 3490 54740 3502
rect 55020 5236 55076 5246
rect 55020 800 55076 5180
rect 55244 5122 55300 6076
rect 56364 6132 56420 6142
rect 56364 5796 56420 6076
rect 57372 6132 57428 6188
rect 57708 6132 57764 43652
rect 57820 13858 57876 13870
rect 57820 13806 57822 13858
rect 57874 13806 57876 13858
rect 57820 13748 57876 13806
rect 57820 13682 57876 13692
rect 57932 6692 57988 56590
rect 58044 55972 58100 55982
rect 58156 55972 58212 56814
rect 58268 56084 58324 56094
rect 58268 55990 58324 56028
rect 58044 55970 58212 55972
rect 58044 55918 58046 55970
rect 58098 55918 58212 55970
rect 58044 55916 58212 55918
rect 58044 55188 58100 55916
rect 58044 55122 58100 55132
rect 58380 53172 58436 60620
rect 58828 60676 58884 60686
rect 58828 60582 58884 60620
rect 59388 60676 59444 60734
rect 59388 60610 59444 60620
rect 59724 60898 59780 60910
rect 59724 60846 59726 60898
rect 59778 60846 59780 60898
rect 59724 60676 59780 60846
rect 60620 60900 60676 60910
rect 60620 60806 60676 60844
rect 60956 60900 61012 60910
rect 60844 60788 60900 60798
rect 60844 60694 60900 60732
rect 59724 60610 59780 60620
rect 60396 60676 60452 60686
rect 59948 60116 60004 60126
rect 59948 60002 60004 60060
rect 59948 59950 59950 60002
rect 60002 59950 60004 60002
rect 58716 59890 58772 59902
rect 58716 59838 58718 59890
rect 58770 59838 58772 59890
rect 58716 59780 58772 59838
rect 58716 59714 58772 59724
rect 58828 59780 58884 59790
rect 59276 59780 59332 59790
rect 58828 59778 59220 59780
rect 58828 59726 58830 59778
rect 58882 59726 59220 59778
rect 58828 59724 59220 59726
rect 58828 59714 58884 59724
rect 59164 59556 59220 59724
rect 59276 59686 59332 59724
rect 59164 59500 59892 59556
rect 59836 59442 59892 59500
rect 59836 59390 59838 59442
rect 59890 59390 59892 59442
rect 59836 59378 59892 59390
rect 59612 59332 59668 59342
rect 59612 59238 59668 59276
rect 59948 59332 60004 59950
rect 60396 60114 60452 60620
rect 60396 60062 60398 60114
rect 60450 60062 60452 60114
rect 60172 59892 60228 59902
rect 60172 59798 60228 59836
rect 60060 59778 60116 59790
rect 60060 59726 60062 59778
rect 60114 59726 60116 59778
rect 60060 59332 60116 59726
rect 60284 59780 60340 59790
rect 60060 59276 60228 59332
rect 59948 59266 60004 59276
rect 59724 59106 59780 59118
rect 59724 59054 59726 59106
rect 59778 59054 59780 59106
rect 59388 58548 59444 58558
rect 59388 58454 59444 58492
rect 58492 58436 58548 58446
rect 58492 58342 58548 58380
rect 58604 58210 58660 58222
rect 58604 58158 58606 58210
rect 58658 58158 58660 58210
rect 58492 57876 58548 57886
rect 58492 57090 58548 57820
rect 58604 57652 58660 58158
rect 59276 58210 59332 58222
rect 59276 58158 59278 58210
rect 59330 58158 59332 58210
rect 59276 57876 59332 58158
rect 59276 57810 59332 57820
rect 59500 57988 59556 57998
rect 59500 57874 59556 57932
rect 59500 57822 59502 57874
rect 59554 57822 59556 57874
rect 59500 57810 59556 57822
rect 58828 57652 58884 57662
rect 58604 57650 58884 57652
rect 58604 57598 58830 57650
rect 58882 57598 58884 57650
rect 58604 57596 58884 57598
rect 58828 57586 58884 57596
rect 59276 57652 59332 57662
rect 59276 57558 59332 57596
rect 59052 57540 59108 57550
rect 59052 57446 59108 57484
rect 59388 57538 59444 57550
rect 59388 57486 59390 57538
rect 59442 57486 59444 57538
rect 58492 57038 58494 57090
rect 58546 57038 58548 57090
rect 58492 57026 58548 57038
rect 58604 57316 58660 57326
rect 58380 53106 58436 53116
rect 58492 55300 58548 55310
rect 58492 43708 58548 55244
rect 58604 51604 58660 57260
rect 59164 57204 59220 57214
rect 59164 56978 59220 57148
rect 59164 56926 59166 56978
rect 59218 56926 59220 56978
rect 59164 56914 59220 56926
rect 59052 56642 59108 56654
rect 59052 56590 59054 56642
rect 59106 56590 59108 56642
rect 59052 56084 59108 56590
rect 59052 56018 59108 56028
rect 58716 55972 58772 55982
rect 58716 55878 58772 55916
rect 59164 52276 59220 52286
rect 59164 52182 59220 52220
rect 59276 52164 59332 52174
rect 59276 52070 59332 52108
rect 58604 51538 58660 51548
rect 59388 51156 59444 57486
rect 59724 56868 59780 59054
rect 60060 59108 60116 59118
rect 60060 59014 60116 59052
rect 59948 58436 60004 58446
rect 59948 58342 60004 58380
rect 59388 51090 59444 51100
rect 59612 56812 59780 56868
rect 59836 58212 59892 58222
rect 59836 57204 59892 58156
rect 58492 43652 58772 43708
rect 57932 6626 57988 6636
rect 57372 6130 57652 6132
rect 57372 6078 57374 6130
rect 57426 6078 57652 6130
rect 57372 6076 57652 6078
rect 57372 6066 57428 6076
rect 56364 5794 56532 5796
rect 56364 5742 56366 5794
rect 56418 5742 56532 5794
rect 56364 5740 56532 5742
rect 56364 5730 56420 5740
rect 55916 5236 55972 5246
rect 55916 5142 55972 5180
rect 55244 5070 55246 5122
rect 55298 5070 55300 5122
rect 55244 5058 55300 5070
rect 55916 4340 55972 4350
rect 55916 4246 55972 4284
rect 55132 4228 55188 4238
rect 55132 4134 55188 4172
rect 55244 3666 55300 3678
rect 55244 3614 55246 3666
rect 55298 3614 55300 3666
rect 55244 3444 55300 3614
rect 55244 3378 55300 3388
rect 55692 3556 55748 3566
rect 56476 3556 56532 5740
rect 57484 5236 57540 5246
rect 57036 5234 57540 5236
rect 57036 5182 57486 5234
rect 57538 5182 57540 5234
rect 57036 5180 57540 5182
rect 56588 4340 56644 4350
rect 56588 4246 56644 4284
rect 56700 3556 56756 3566
rect 56476 3554 56756 3556
rect 56476 3502 56702 3554
rect 56754 3502 56756 3554
rect 56476 3500 56756 3502
rect 55692 800 55748 3500
rect 56700 3490 56756 3500
rect 56364 3444 56420 3454
rect 56364 800 56420 3388
rect 57036 800 57092 5180
rect 57484 5170 57540 5180
rect 57596 4338 57652 6076
rect 57708 6066 57764 6076
rect 58156 6356 58212 6366
rect 58156 6132 58212 6300
rect 58156 6130 58436 6132
rect 58156 6078 58158 6130
rect 58210 6078 58436 6130
rect 58156 6076 58436 6078
rect 58156 6066 58212 6076
rect 58380 4900 58436 6076
rect 58716 6130 58772 43652
rect 59612 6244 59668 56812
rect 59724 56644 59780 56654
rect 59836 56644 59892 57148
rect 59724 56642 59892 56644
rect 59724 56590 59726 56642
rect 59778 56590 59892 56642
rect 59724 56588 59892 56590
rect 59724 56578 59780 56588
rect 59836 52164 59892 52174
rect 59836 52070 59892 52108
rect 60172 51380 60228 59276
rect 60284 59218 60340 59724
rect 60284 59166 60286 59218
rect 60338 59166 60340 59218
rect 60284 59154 60340 59166
rect 60396 59108 60452 60062
rect 60732 60674 60788 60686
rect 60732 60622 60734 60674
rect 60786 60622 60788 60674
rect 60620 60004 60676 60014
rect 60620 59910 60676 59948
rect 60396 59042 60452 59052
rect 60396 58548 60452 58558
rect 60396 58454 60452 58492
rect 60284 52388 60340 52398
rect 60284 52294 60340 52332
rect 60396 52276 60452 52286
rect 60396 52182 60452 52220
rect 59948 51324 60228 51380
rect 59948 31948 60004 51324
rect 59836 31892 60004 31948
rect 60172 51156 60228 51166
rect 59836 6356 59892 31892
rect 59836 6290 59892 6300
rect 59612 6178 59668 6188
rect 58716 6078 58718 6130
rect 58770 6078 58772 6130
rect 58492 5124 58548 5134
rect 58716 5124 58772 6078
rect 58492 5122 58772 5124
rect 58492 5070 58494 5122
rect 58546 5070 58772 5122
rect 58492 5068 58772 5070
rect 59164 6132 59220 6142
rect 58492 5058 58548 5068
rect 58380 4844 58548 4900
rect 57596 4286 57598 4338
rect 57650 4286 57652 4338
rect 57596 4274 57652 4286
rect 57708 4228 57764 4238
rect 57372 3668 57428 3678
rect 57372 3574 57428 3612
rect 57708 800 57764 4172
rect 58156 4226 58212 4238
rect 58156 4174 58158 4226
rect 58210 4174 58212 4226
rect 58156 3556 58212 4174
rect 58156 3490 58212 3500
rect 58380 3668 58436 3678
rect 58380 800 58436 3612
rect 58492 3554 58548 4844
rect 59164 4340 59220 6076
rect 60172 6132 60228 51100
rect 60732 50428 60788 60622
rect 60956 60116 61012 60844
rect 61740 60788 61796 60798
rect 61068 60676 61124 60686
rect 61068 60582 61124 60620
rect 61292 60564 61348 60574
rect 61292 60470 61348 60508
rect 60956 59444 61012 60060
rect 61516 60228 61572 60238
rect 61516 60114 61572 60172
rect 61516 60062 61518 60114
rect 61570 60062 61572 60114
rect 61516 60050 61572 60062
rect 61404 59780 61460 59790
rect 61404 59686 61460 59724
rect 61068 59444 61124 59454
rect 60956 59442 61124 59444
rect 60956 59390 61070 59442
rect 61122 59390 61124 59442
rect 60956 59388 61124 59390
rect 61068 59378 61124 59388
rect 61292 59218 61348 59230
rect 61292 59166 61294 59218
rect 61346 59166 61348 59218
rect 61292 59108 61348 59166
rect 61740 59108 61796 60732
rect 61852 60786 61908 61292
rect 62300 61012 62356 61022
rect 62300 60918 62356 60956
rect 62524 60900 62580 60910
rect 62524 60806 62580 60844
rect 61852 60734 61854 60786
rect 61906 60734 61908 60786
rect 61852 60722 61908 60734
rect 62076 60676 62132 60686
rect 62076 60582 62132 60620
rect 62412 60674 62468 60686
rect 62412 60622 62414 60674
rect 62466 60622 62468 60674
rect 62076 60228 62132 60238
rect 62076 60114 62132 60172
rect 62076 60062 62078 60114
rect 62130 60062 62132 60114
rect 62076 60050 62132 60062
rect 61852 59108 61908 59118
rect 61292 59106 61908 59108
rect 61292 59054 61854 59106
rect 61906 59054 61908 59106
rect 61292 59052 61908 59054
rect 61292 57316 61348 59052
rect 61852 59042 61908 59052
rect 61292 57250 61348 57260
rect 61404 52276 61460 52286
rect 61404 52182 61460 52220
rect 60732 50372 61236 50428
rect 59500 5234 59556 5246
rect 59500 5182 59502 5234
rect 59554 5182 59556 5234
rect 59276 4340 59332 4350
rect 59164 4338 59332 4340
rect 59164 4286 59278 4338
rect 59330 4286 59332 4338
rect 59164 4284 59332 4286
rect 59276 4274 59332 4284
rect 58492 3502 58494 3554
rect 58546 3502 58548 3554
rect 58492 3490 58548 3502
rect 59388 3444 59444 3454
rect 59388 3350 59444 3388
rect 59500 2660 59556 5182
rect 60172 5124 60228 6076
rect 60284 6692 60340 6702
rect 60284 6132 60340 6636
rect 61068 6244 61124 6254
rect 60732 6132 60788 6142
rect 60284 6130 60676 6132
rect 60284 6078 60286 6130
rect 60338 6078 60676 6130
rect 60284 6076 60676 6078
rect 60284 6066 60340 6076
rect 60284 5124 60340 5134
rect 60172 5122 60340 5124
rect 60172 5070 60286 5122
rect 60338 5070 60340 5122
rect 60172 5068 60340 5070
rect 60284 5058 60340 5068
rect 59948 4228 60004 4238
rect 59948 4134 60004 4172
rect 59052 2604 59556 2660
rect 59724 3556 59780 3566
rect 59052 800 59108 2604
rect 59724 800 59780 3500
rect 60620 3554 60676 6076
rect 60732 6038 60788 6076
rect 60620 3502 60622 3554
rect 60674 3502 60676 3554
rect 60620 3490 60676 3502
rect 60956 5236 61012 5246
rect 60396 3444 60452 3454
rect 60396 800 60452 3388
rect 60956 2548 61012 5180
rect 61068 4338 61124 6188
rect 61180 6130 61236 50372
rect 62076 6356 62132 6366
rect 61180 6078 61182 6130
rect 61234 6078 61236 6130
rect 61180 5124 61236 6078
rect 61628 6244 61684 6254
rect 61628 6130 61684 6188
rect 61628 6078 61630 6130
rect 61682 6078 61684 6130
rect 61628 6066 61684 6078
rect 62076 6132 62132 6300
rect 62076 6130 62244 6132
rect 62076 6078 62078 6130
rect 62130 6078 62244 6130
rect 62076 6076 62244 6078
rect 62076 6066 62132 6076
rect 62076 5236 62132 5246
rect 62076 5142 62132 5180
rect 61404 5124 61460 5134
rect 61180 5122 61460 5124
rect 61180 5070 61406 5122
rect 61458 5070 61460 5122
rect 61180 5068 61460 5070
rect 61404 5058 61460 5068
rect 61068 4286 61070 4338
rect 61122 4286 61124 4338
rect 61068 4274 61124 4286
rect 61740 4228 61796 4238
rect 61292 3668 61348 3678
rect 61292 3574 61348 3612
rect 60956 2492 61124 2548
rect 61068 800 61124 2492
rect 61740 800 61796 4172
rect 61852 4226 61908 4238
rect 61852 4174 61854 4226
rect 61906 4174 61908 4226
rect 61852 3556 61908 4174
rect 62188 3556 62244 6076
rect 62412 4340 62468 60622
rect 62748 57652 62804 57662
rect 62748 57558 62804 57596
rect 62636 57428 62692 57438
rect 62636 57334 62692 57372
rect 62860 6244 62916 62132
rect 62972 62132 63140 62188
rect 63196 62914 63252 62926
rect 63196 62862 63198 62914
rect 63250 62862 63252 62914
rect 62972 61460 63028 62132
rect 62972 61394 63028 61404
rect 63196 60900 63252 62862
rect 63308 62914 63364 62926
rect 63308 62862 63310 62914
rect 63362 62862 63364 62914
rect 63308 62804 63364 62862
rect 63308 62738 63364 62748
rect 63644 62578 63700 63084
rect 63644 62526 63646 62578
rect 63698 62526 63700 62578
rect 63644 62514 63700 62526
rect 63868 62356 63924 62366
rect 63868 62262 63924 62300
rect 63980 62354 64036 63756
rect 64876 63250 64932 64204
rect 64876 63198 64878 63250
rect 64930 63198 64932 63250
rect 64876 63186 64932 63198
rect 65100 64148 65156 64158
rect 65100 63924 65156 64092
rect 65100 62916 65156 63868
rect 65212 63140 65268 64430
rect 65324 64484 65380 64494
rect 65324 64390 65380 64428
rect 65548 64148 65604 64766
rect 65548 64082 65604 64092
rect 65660 64876 65828 64932
rect 66108 64876 66388 64932
rect 65548 63924 65604 63934
rect 65548 63830 65604 63868
rect 65212 63084 65492 63140
rect 65212 62916 65268 62926
rect 65100 62914 65268 62916
rect 65100 62862 65214 62914
rect 65266 62862 65268 62914
rect 65100 62860 65268 62862
rect 65212 62850 65268 62860
rect 63980 62302 63982 62354
rect 64034 62302 64036 62354
rect 63980 62290 64036 62302
rect 65324 62468 65380 62478
rect 63756 62242 63812 62254
rect 63756 62190 63758 62242
rect 63810 62190 63812 62242
rect 63644 62132 63700 62142
rect 63308 61460 63364 61470
rect 63308 61366 63364 61404
rect 63644 61458 63700 62076
rect 63644 61406 63646 61458
rect 63698 61406 63700 61458
rect 63196 60834 63252 60844
rect 63420 61124 63476 61134
rect 63084 60788 63140 60798
rect 63084 60694 63140 60732
rect 63196 57652 63252 57662
rect 63196 57558 63252 57596
rect 63420 6692 63476 61068
rect 63420 6626 63476 6636
rect 63532 60900 63588 60910
rect 63532 6356 63588 60844
rect 63644 60788 63700 61406
rect 63644 60722 63700 60732
rect 63532 6290 63588 6300
rect 62860 6178 62916 6188
rect 63756 6132 63812 62190
rect 64316 62244 64372 62254
rect 64316 62150 64372 62188
rect 64204 61572 64260 61582
rect 64204 61478 64260 61516
rect 65324 61012 65380 62412
rect 64652 61010 65380 61012
rect 64652 60958 65326 61010
rect 65378 60958 65380 61010
rect 64652 60956 65380 60958
rect 64652 60898 64708 60956
rect 65324 60946 65380 60956
rect 64652 60846 64654 60898
rect 64706 60846 64708 60898
rect 64652 60834 64708 60846
rect 64540 60564 64596 60574
rect 64540 60470 64596 60508
rect 63532 5236 63588 5246
rect 62412 4274 62468 4284
rect 63196 5234 63588 5236
rect 63196 5182 63534 5234
rect 63586 5182 63588 5234
rect 63196 5180 63588 5182
rect 63084 4228 63140 4238
rect 63084 4134 63140 4172
rect 62524 3668 62580 3678
rect 62412 3556 62468 3566
rect 62188 3554 62468 3556
rect 62188 3502 62414 3554
rect 62466 3502 62468 3554
rect 62188 3500 62468 3502
rect 61852 3490 61908 3500
rect 62412 3490 62468 3500
rect 62524 1764 62580 3612
rect 63196 2548 63252 5180
rect 63532 5170 63588 5180
rect 63756 5124 63812 6076
rect 63756 5058 63812 5068
rect 64204 6244 64260 6254
rect 64204 6130 64260 6188
rect 65436 6244 65492 63084
rect 65660 62188 65716 64876
rect 65772 64706 65828 64718
rect 65772 64654 65774 64706
rect 65826 64654 65828 64706
rect 65772 64596 65828 64654
rect 65772 64530 65828 64540
rect 65884 64148 65940 64158
rect 65884 64054 65940 64092
rect 66108 63700 66164 64876
rect 66444 64818 66500 65772
rect 66444 64766 66446 64818
rect 66498 64766 66500 64818
rect 66444 64754 66500 64766
rect 66556 65716 66612 65726
rect 66332 64596 66388 64606
rect 66332 64502 66388 64540
rect 66444 64372 66500 64382
rect 66444 64146 66500 64316
rect 66444 64094 66446 64146
rect 66498 64094 66500 64146
rect 66444 64082 66500 64094
rect 66108 63644 66388 63700
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 66108 62914 66164 62926
rect 66108 62862 66110 62914
rect 66162 62862 66164 62914
rect 65660 62132 65828 62188
rect 65772 6916 65828 62132
rect 66108 62132 66164 62862
rect 66108 62066 66164 62076
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 65772 6860 65940 6916
rect 65436 6178 65492 6188
rect 65772 6356 65828 6366
rect 64204 6078 64206 6130
rect 64258 6078 64260 6130
rect 63868 4340 63924 4350
rect 63868 4246 63924 4284
rect 63756 4228 63812 4238
rect 63308 3444 63364 3454
rect 63308 3350 63364 3388
rect 62412 1708 62580 1764
rect 63084 2492 63252 2548
rect 62412 800 62468 1708
rect 63084 800 63140 2492
rect 63756 800 63812 4172
rect 64204 3780 64260 6078
rect 65324 6132 65380 6142
rect 65324 6038 65380 6076
rect 65772 6130 65828 6300
rect 65772 6078 65774 6130
rect 65826 6078 65828 6130
rect 65548 5236 65604 5246
rect 65100 5234 65604 5236
rect 65100 5182 65550 5234
rect 65602 5182 65604 5234
rect 65100 5180 65604 5182
rect 64316 5124 64372 5134
rect 64316 5030 64372 5068
rect 64540 4340 64596 4350
rect 64540 4246 64596 4284
rect 64204 3724 64596 3780
rect 64428 3556 64484 3566
rect 64428 800 64484 3500
rect 64540 3554 64596 3724
rect 64540 3502 64542 3554
rect 64594 3502 64596 3554
rect 64540 3490 64596 3502
rect 65100 800 65156 5180
rect 65548 5170 65604 5180
rect 65660 4340 65716 4350
rect 65772 4340 65828 6078
rect 65884 5908 65940 6860
rect 66108 6692 66164 6702
rect 66108 6132 66164 6636
rect 66332 6692 66388 63644
rect 66556 62188 66612 65660
rect 66668 64372 66724 65884
rect 67004 65828 67060 65838
rect 67004 64818 67060 65772
rect 67676 65492 67732 65998
rect 67788 66052 67844 66062
rect 67788 65958 67844 65996
rect 68012 65828 68068 67172
rect 68348 67172 68404 68348
rect 68796 68402 68852 68414
rect 68796 68350 68798 68402
rect 68850 68350 68852 68402
rect 68572 68068 68628 68078
rect 68572 67954 68628 68012
rect 68572 67902 68574 67954
rect 68626 67902 68628 67954
rect 68572 67890 68628 67902
rect 68460 67618 68516 67630
rect 68460 67566 68462 67618
rect 68514 67566 68516 67618
rect 68460 67396 68516 67566
rect 68460 67340 68628 67396
rect 68460 67172 68516 67182
rect 68348 67170 68516 67172
rect 68348 67118 68462 67170
rect 68514 67118 68516 67170
rect 68348 67116 68516 67118
rect 68460 67106 68516 67116
rect 68236 67060 68292 67070
rect 68236 66966 68292 67004
rect 68348 66946 68404 66958
rect 68348 66894 68350 66946
rect 68402 66894 68404 66946
rect 68348 66724 68404 66894
rect 68348 66658 68404 66668
rect 68124 66500 68180 66510
rect 68124 66386 68180 66444
rect 68348 66500 68404 66510
rect 68572 66500 68628 67340
rect 68796 67060 68852 68350
rect 69132 67228 69188 72268
rect 69580 72322 69636 72334
rect 69580 72270 69582 72322
rect 69634 72270 69636 72322
rect 69580 71988 69636 72270
rect 69580 71922 69636 71932
rect 69468 70196 69524 70206
rect 69468 70102 69524 70140
rect 69356 70084 69412 70094
rect 69356 69298 69412 70028
rect 69356 69246 69358 69298
rect 69410 69246 69412 69298
rect 69356 69234 69412 69246
rect 69692 69300 69748 69310
rect 69692 69206 69748 69244
rect 69468 67956 69524 67966
rect 69468 67862 69524 67900
rect 69356 67618 69412 67630
rect 69356 67566 69358 67618
rect 69410 67566 69412 67618
rect 69356 67228 69412 67566
rect 69804 67228 69860 72604
rect 71820 72434 71876 73164
rect 72492 73218 72548 73230
rect 72492 73166 72494 73218
rect 72546 73166 72548 73218
rect 72156 72548 72212 72558
rect 72156 72454 72212 72492
rect 72492 72548 72548 73166
rect 72492 72482 72548 72492
rect 73052 72548 73108 72558
rect 73052 72454 73108 72492
rect 71820 72382 71822 72434
rect 71874 72382 71876 72434
rect 71820 72370 71876 72382
rect 73276 72434 73332 73276
rect 73388 73108 73444 73838
rect 73724 73554 73780 74844
rect 75068 74900 75124 74910
rect 75068 74806 75124 74844
rect 76860 74898 76916 74910
rect 76860 74846 76862 74898
rect 76914 74846 76916 74898
rect 76076 74786 76132 74798
rect 76076 74734 76078 74786
rect 76130 74734 76132 74786
rect 76076 74564 76132 74734
rect 76076 74498 76132 74508
rect 73724 73502 73726 73554
rect 73778 73502 73780 73554
rect 73724 73490 73780 73502
rect 74060 74004 74116 74014
rect 73836 73444 73892 73454
rect 73612 73108 73668 73118
rect 73388 73106 73668 73108
rect 73388 73054 73614 73106
rect 73666 73054 73668 73106
rect 73388 73052 73668 73054
rect 73612 72660 73668 73052
rect 73612 72594 73668 72604
rect 73276 72382 73278 72434
rect 73330 72382 73332 72434
rect 73276 72370 73332 72382
rect 73724 72548 73780 72558
rect 72492 72324 72548 72334
rect 72492 71986 72548 72268
rect 73724 72212 73780 72492
rect 73836 72436 73892 73388
rect 74060 72658 74116 73948
rect 76860 74004 76916 74846
rect 77868 74786 77924 74798
rect 77868 74734 77870 74786
rect 77922 74734 77924 74786
rect 76860 73938 76916 73948
rect 77308 74004 77364 74014
rect 77308 73910 77364 73948
rect 77756 73892 77812 73902
rect 77532 73890 77812 73892
rect 77532 73838 77758 73890
rect 77810 73838 77812 73890
rect 77532 73836 77812 73838
rect 75068 73332 75124 73342
rect 75068 73238 75124 73276
rect 76860 73330 76916 73342
rect 76860 73278 76862 73330
rect 76914 73278 76916 73330
rect 76076 73218 76132 73230
rect 76076 73166 76078 73218
rect 76130 73166 76132 73218
rect 74060 72606 74062 72658
rect 74114 72606 74116 72658
rect 74060 72594 74116 72606
rect 74172 72660 74228 72670
rect 74172 72566 74228 72604
rect 74620 72660 74676 72670
rect 74620 72566 74676 72604
rect 75068 72548 75124 72558
rect 75068 72454 75124 72492
rect 76076 72548 76132 73166
rect 76076 72482 76132 72492
rect 73836 72370 73892 72380
rect 74060 72436 74116 72446
rect 73948 72322 74004 72334
rect 73948 72270 73950 72322
rect 74002 72270 74004 72322
rect 73724 72156 73892 72212
rect 72492 71934 72494 71986
rect 72546 71934 72548 71986
rect 72492 71922 72548 71934
rect 73388 71988 73444 71998
rect 73388 71894 73444 71932
rect 71148 71876 71204 71886
rect 71148 71782 71204 71820
rect 70700 71764 70756 71774
rect 70700 71670 70756 71708
rect 71484 71764 71540 71774
rect 71484 71670 71540 71708
rect 72268 71764 72324 71774
rect 72268 71670 72324 71708
rect 72828 71764 72884 71774
rect 70588 71652 70644 71662
rect 70588 70866 70644 71596
rect 71708 70980 71764 70990
rect 71708 70978 71876 70980
rect 71708 70926 71710 70978
rect 71762 70926 71876 70978
rect 71708 70924 71876 70926
rect 71708 70914 71764 70924
rect 70588 70814 70590 70866
rect 70642 70814 70644 70866
rect 70588 70802 70644 70814
rect 70924 70866 70980 70878
rect 70924 70814 70926 70866
rect 70978 70814 70980 70866
rect 70140 70756 70196 70766
rect 70140 70662 70196 70700
rect 70924 70756 70980 70814
rect 70924 70690 70980 70700
rect 71820 70756 71876 70924
rect 71932 70868 71988 70878
rect 71932 70774 71988 70812
rect 71260 70644 71316 70654
rect 71260 70418 71316 70588
rect 71260 70366 71262 70418
rect 71314 70366 71316 70418
rect 71260 70354 71316 70366
rect 69916 70308 69972 70318
rect 69916 70214 69972 70252
rect 70252 70196 70308 70206
rect 70252 70102 70308 70140
rect 70924 70196 70980 70206
rect 70252 69300 70308 69310
rect 69020 67172 69188 67228
rect 69244 67172 69412 67228
rect 69692 67172 69860 67228
rect 69916 68516 69972 68526
rect 70252 68516 70308 69244
rect 70588 69300 70644 69310
rect 70588 69206 70644 69244
rect 69916 68514 70308 68516
rect 69916 68462 69918 68514
rect 69970 68462 70308 68514
rect 69916 68460 70308 68462
rect 69916 67228 69972 68460
rect 70028 68068 70084 68078
rect 70028 67954 70084 68012
rect 70028 67902 70030 67954
rect 70082 67902 70084 67954
rect 70028 67890 70084 67902
rect 69916 67172 70420 67228
rect 68908 67060 68964 67070
rect 68796 67058 68964 67060
rect 68796 67006 68910 67058
rect 68962 67006 68964 67058
rect 68796 67004 68964 67006
rect 68908 66994 68964 67004
rect 68684 66948 68740 66958
rect 68684 66946 68852 66948
rect 68684 66894 68686 66946
rect 68738 66894 68852 66946
rect 68684 66892 68852 66894
rect 68684 66882 68740 66892
rect 68348 66498 68628 66500
rect 68348 66446 68350 66498
rect 68402 66446 68628 66498
rect 68348 66444 68628 66446
rect 68796 66500 68852 66892
rect 68348 66434 68404 66444
rect 68124 66334 68126 66386
rect 68178 66334 68180 66386
rect 68124 66322 68180 66334
rect 68684 66388 68740 66398
rect 68572 66052 68628 66062
rect 68012 65772 68180 65828
rect 68124 65604 68180 65772
rect 68348 65716 68404 65726
rect 68124 65548 68292 65604
rect 68012 65492 68068 65502
rect 67676 65490 68068 65492
rect 67676 65438 68014 65490
rect 68066 65438 68068 65490
rect 67676 65436 68068 65438
rect 67228 65380 67284 65390
rect 67228 65378 67508 65380
rect 67228 65326 67230 65378
rect 67282 65326 67508 65378
rect 67228 65324 67508 65326
rect 67228 65314 67284 65324
rect 67004 64766 67006 64818
rect 67058 64766 67060 64818
rect 67004 64754 67060 64766
rect 66668 64306 66724 64316
rect 67452 64706 67508 65324
rect 67452 64654 67454 64706
rect 67506 64654 67508 64706
rect 66332 6626 66388 6636
rect 66444 62132 66612 62188
rect 66668 64036 66724 64046
rect 66668 63922 66724 63980
rect 67452 64036 67508 64654
rect 67788 64484 67844 64494
rect 67788 64390 67844 64428
rect 68012 64484 68068 65436
rect 68236 65490 68292 65548
rect 68236 65438 68238 65490
rect 68290 65438 68292 65490
rect 68236 65426 68292 65438
rect 68012 64418 68068 64428
rect 68124 65378 68180 65390
rect 68124 65326 68126 65378
rect 68178 65326 68180 65378
rect 67676 64148 67732 64158
rect 67676 64054 67732 64092
rect 67452 63970 67508 63980
rect 66668 63870 66670 63922
rect 66722 63870 66724 63922
rect 66668 62132 66724 63870
rect 67004 63924 67060 63934
rect 67004 63250 67060 63868
rect 67340 63924 67396 63934
rect 67340 63830 67396 63868
rect 67004 63198 67006 63250
rect 67058 63198 67060 63250
rect 67004 63186 67060 63198
rect 66332 6244 66388 6254
rect 66220 6132 66276 6142
rect 66108 6130 66276 6132
rect 66108 6078 66222 6130
rect 66274 6078 66276 6130
rect 66108 6076 66276 6078
rect 65884 5842 65940 5852
rect 66220 5682 66276 6076
rect 66220 5630 66222 5682
rect 66274 5630 66276 5682
rect 66220 5618 66276 5630
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 66332 5122 66388 6188
rect 66444 6132 66500 62132
rect 66668 62066 66724 62076
rect 66668 60116 66724 60126
rect 66668 60022 66724 60060
rect 67228 60116 67284 60126
rect 67228 60022 67284 60060
rect 66556 60004 66612 60014
rect 66556 59910 66612 59948
rect 68124 50428 68180 65326
rect 68236 62580 68292 62590
rect 68348 62580 68404 65660
rect 68460 65492 68516 65502
rect 68460 65378 68516 65436
rect 68460 65326 68462 65378
rect 68514 65326 68516 65378
rect 68460 64596 68516 65326
rect 68460 64148 68516 64540
rect 68460 64082 68516 64092
rect 68348 62524 68516 62580
rect 68236 62468 68292 62524
rect 68236 62412 68404 62468
rect 68236 62244 68292 62254
rect 68236 62150 68292 62188
rect 68348 62242 68404 62412
rect 68348 62190 68350 62242
rect 68402 62190 68404 62242
rect 68348 62178 68404 62190
rect 67900 50372 68180 50428
rect 67676 6692 67732 6702
rect 66444 6066 66500 6076
rect 66780 6244 66836 6254
rect 66780 6130 66836 6188
rect 66780 6078 66782 6130
rect 66834 6078 66836 6130
rect 66780 6066 66836 6078
rect 67228 6132 67284 6142
rect 67228 5796 67284 6076
rect 67676 6130 67732 6636
rect 67676 6078 67678 6130
rect 67730 6078 67732 6130
rect 67228 5794 67396 5796
rect 67228 5742 67230 5794
rect 67282 5742 67396 5794
rect 67228 5740 67396 5742
rect 67228 5730 67284 5740
rect 66332 5070 66334 5122
rect 66386 5070 66388 5122
rect 66332 5058 66388 5070
rect 66556 5682 66612 5694
rect 66556 5630 66558 5682
rect 66610 5630 66612 5682
rect 65660 4338 65828 4340
rect 65660 4286 65662 4338
rect 65714 4286 65828 4338
rect 65660 4284 65828 4286
rect 65660 4274 65716 4284
rect 66108 4228 66164 4238
rect 66108 4134 66164 4172
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 65212 3668 65268 3678
rect 65212 3574 65268 3612
rect 65772 3556 65828 3566
rect 65772 800 65828 3500
rect 66556 3554 66612 5630
rect 67116 5236 67172 5246
rect 67004 3668 67060 3678
rect 67004 3574 67060 3612
rect 66556 3502 66558 3554
rect 66610 3502 66612 3554
rect 66556 3490 66612 3502
rect 66444 3444 66500 3454
rect 66444 800 66500 3388
rect 67116 800 67172 5180
rect 67340 5122 67396 5740
rect 67340 5070 67342 5122
rect 67394 5070 67396 5122
rect 67340 5058 67396 5070
rect 67452 4340 67508 4350
rect 67676 4340 67732 6078
rect 67900 4452 67956 50372
rect 68012 49924 68068 49934
rect 68012 49140 68068 49868
rect 68012 49008 68068 49084
rect 68124 48804 68180 48814
rect 68124 48710 68180 48748
rect 68460 6132 68516 62524
rect 68572 50428 68628 65996
rect 68684 65490 68740 66332
rect 68684 65438 68686 65490
rect 68738 65438 68740 65490
rect 68684 65426 68740 65438
rect 68796 65492 68852 66444
rect 68796 65426 68852 65436
rect 68684 64484 68740 64494
rect 68684 64034 68740 64428
rect 68684 63982 68686 64034
rect 68738 63982 68740 64034
rect 68684 63970 68740 63982
rect 69020 64034 69076 67172
rect 69244 66388 69300 67172
rect 69356 66948 69412 66958
rect 69356 66854 69412 66892
rect 69244 66322 69300 66332
rect 69356 64596 69412 64606
rect 69356 64502 69412 64540
rect 69020 63982 69022 64034
rect 69074 63982 69076 64034
rect 68796 62580 68852 62590
rect 68796 62486 68852 62524
rect 69020 62188 69076 63982
rect 69692 64482 69748 67172
rect 69692 64430 69694 64482
rect 69746 64430 69748 64482
rect 69692 62188 69748 64430
rect 69020 62132 69300 62188
rect 69692 62132 70308 62188
rect 68684 50708 68740 50718
rect 68684 50614 68740 50652
rect 68572 50372 68740 50428
rect 68572 49140 68628 49150
rect 68572 49046 68628 49084
rect 68684 31948 68740 50372
rect 68908 49812 68964 49822
rect 68908 49718 68964 49756
rect 69244 49812 69300 62132
rect 70028 50820 70084 50830
rect 69356 50708 69412 50718
rect 69356 50614 69412 50652
rect 70028 50706 70084 50764
rect 70028 50654 70030 50706
rect 70082 50654 70084 50706
rect 70028 50642 70084 50654
rect 69468 50370 69524 50382
rect 69468 50318 69470 50370
rect 69522 50318 69524 50370
rect 69468 50036 69524 50318
rect 70140 50370 70196 50382
rect 70140 50318 70142 50370
rect 70194 50318 70196 50370
rect 69804 50036 69860 50046
rect 69468 50034 69860 50036
rect 69468 49982 69806 50034
rect 69858 49982 69860 50034
rect 69468 49980 69860 49982
rect 69804 49970 69860 49980
rect 69244 49746 69300 49756
rect 69580 49812 69636 49850
rect 69580 49746 69636 49756
rect 69916 49812 69972 49822
rect 70140 49812 70196 50318
rect 70252 50036 70308 62132
rect 70252 49970 70308 49980
rect 70252 49812 70308 49822
rect 70140 49810 70308 49812
rect 70140 49758 70254 49810
rect 70306 49758 70308 49810
rect 70140 49756 70308 49758
rect 69692 49698 69748 49710
rect 69692 49646 69694 49698
rect 69746 49646 69748 49698
rect 69580 49588 69636 49598
rect 69580 49138 69636 49532
rect 69580 49086 69582 49138
rect 69634 49086 69636 49138
rect 69580 49074 69636 49086
rect 69356 49028 69412 49038
rect 68908 49026 69412 49028
rect 68908 48974 69358 49026
rect 69410 48974 69412 49026
rect 68908 48972 69412 48974
rect 68796 48468 68852 48478
rect 68796 48354 68852 48412
rect 68908 48466 68964 48972
rect 69356 48962 69412 48972
rect 69692 48580 69748 49646
rect 69916 49476 69972 49756
rect 70252 49746 70308 49756
rect 70028 49700 70084 49710
rect 70028 49606 70084 49644
rect 69916 49420 70084 49476
rect 69804 48804 69860 48814
rect 69804 48710 69860 48748
rect 69916 48802 69972 48814
rect 69916 48750 69918 48802
rect 69970 48750 69972 48802
rect 69692 48524 69860 48580
rect 68908 48414 68910 48466
rect 68962 48414 68964 48466
rect 68908 48402 68964 48414
rect 69356 48468 69412 48478
rect 69356 48374 69412 48412
rect 68796 48302 68798 48354
rect 68850 48302 68852 48354
rect 68796 48290 68852 48302
rect 69468 48356 69524 48366
rect 68572 31892 68740 31948
rect 68572 6244 68628 31892
rect 69468 8428 69524 48300
rect 69804 38668 69860 48524
rect 69916 48356 69972 48750
rect 69916 48290 69972 48300
rect 70028 48802 70084 49420
rect 70028 48750 70030 48802
rect 70082 48750 70084 48802
rect 69916 48132 69972 48142
rect 70028 48132 70084 48750
rect 69916 48130 70084 48132
rect 69916 48078 69918 48130
rect 69970 48078 70084 48130
rect 69916 48076 70084 48078
rect 69916 48066 69972 48076
rect 69244 8372 69524 8428
rect 69692 38612 69860 38668
rect 68572 6178 68628 6188
rect 69132 6244 69188 6254
rect 68460 6066 68516 6076
rect 69020 6132 69076 6142
rect 69020 6038 69076 6076
rect 68124 5908 68180 5918
rect 68124 5794 68180 5852
rect 68124 5742 68126 5794
rect 68178 5742 68180 5794
rect 68012 5236 68068 5246
rect 68012 5142 68068 5180
rect 67900 4386 67956 4396
rect 67452 4338 67732 4340
rect 67452 4286 67454 4338
rect 67506 4286 67732 4338
rect 67452 4284 67732 4286
rect 67452 4274 67508 4284
rect 67788 4228 67844 4238
rect 67788 800 67844 4172
rect 67900 4226 67956 4238
rect 67900 4174 67902 4226
rect 67954 4174 67956 4226
rect 67900 3556 67956 4174
rect 68124 3556 68180 5742
rect 69132 4338 69188 6188
rect 69244 5796 69300 8372
rect 69468 6244 69524 6254
rect 69244 5730 69300 5740
rect 69356 6132 69412 6142
rect 69356 5122 69412 6076
rect 69468 6130 69524 6188
rect 69468 6078 69470 6130
rect 69522 6078 69524 6130
rect 69468 6066 69524 6078
rect 69692 5460 69748 38612
rect 69692 5394 69748 5404
rect 70028 5236 70084 5246
rect 69356 5070 69358 5122
rect 69410 5070 69412 5122
rect 69356 5058 69412 5070
rect 69468 5234 70084 5236
rect 69468 5182 70030 5234
rect 70082 5182 70084 5234
rect 69468 5180 70084 5182
rect 69132 4286 69134 4338
rect 69186 4286 69188 4338
rect 69132 4274 69188 4286
rect 68460 3556 68516 3566
rect 68124 3554 68516 3556
rect 68124 3502 68462 3554
rect 68514 3502 68516 3554
rect 68124 3500 68516 3502
rect 67900 3490 67956 3500
rect 68460 3490 68516 3500
rect 68572 3556 68628 3566
rect 68572 1764 68628 3500
rect 69356 3444 69412 3454
rect 69356 3350 69412 3388
rect 69468 2660 69524 5180
rect 70028 5170 70084 5180
rect 70364 4564 70420 67172
rect 70700 50820 70756 50830
rect 70700 50706 70756 50764
rect 70700 50654 70702 50706
rect 70754 50654 70756 50706
rect 70700 50642 70756 50654
rect 70700 49700 70756 49710
rect 70700 49138 70756 49644
rect 70700 49086 70702 49138
rect 70754 49086 70756 49138
rect 70700 49074 70756 49086
rect 70924 8428 70980 70140
rect 71708 70196 71764 70206
rect 71708 70102 71764 70140
rect 71148 69188 71204 69198
rect 71148 69094 71204 69132
rect 71820 50428 71876 70700
rect 72380 70756 72436 70766
rect 72380 70662 72436 70700
rect 72828 70754 72884 71708
rect 73500 71652 73556 71662
rect 73500 71650 73668 71652
rect 73500 71598 73502 71650
rect 73554 71598 73668 71650
rect 73500 71596 73668 71598
rect 73500 71586 73556 71596
rect 72828 70702 72830 70754
rect 72882 70702 72884 70754
rect 72828 50428 72884 70702
rect 73612 70756 73668 71596
rect 73724 70756 73780 70766
rect 73612 70754 73780 70756
rect 73612 70702 73726 70754
rect 73778 70702 73780 70754
rect 73612 70700 73780 70702
rect 73612 50428 73668 70700
rect 73724 70690 73780 70700
rect 73836 50428 73892 72156
rect 73948 71988 74004 72270
rect 73948 71922 74004 71932
rect 74060 71986 74116 72380
rect 76860 72324 76916 73278
rect 76860 72258 76916 72268
rect 74060 71934 74062 71986
rect 74114 71934 74116 71986
rect 74060 71922 74116 71934
rect 75068 71762 75124 71774
rect 75068 71710 75070 71762
rect 75122 71710 75124 71762
rect 74172 71650 74228 71662
rect 74172 71598 74174 71650
rect 74226 71598 74228 71650
rect 74172 70756 74228 71598
rect 75068 70868 75124 71710
rect 76860 71762 76916 71774
rect 76860 71710 76862 71762
rect 76914 71710 76916 71762
rect 76076 71650 76132 71662
rect 76076 71598 76078 71650
rect 76130 71598 76132 71650
rect 76076 71204 76132 71598
rect 76076 71138 76132 71148
rect 75068 70802 75124 70812
rect 74396 70756 74452 70766
rect 74172 70754 74452 70756
rect 74172 70702 74398 70754
rect 74450 70702 74452 70754
rect 74172 70700 74452 70702
rect 74396 67228 74452 70700
rect 76860 70644 76916 71710
rect 76860 70578 76916 70588
rect 76860 70194 76916 70206
rect 76860 70142 76862 70194
rect 76914 70142 76916 70194
rect 76524 69298 76580 69310
rect 76524 69246 76526 69298
rect 76578 69246 76580 69298
rect 76188 69186 76244 69198
rect 76188 69134 76190 69186
rect 76242 69134 76244 69186
rect 76188 68740 76244 69134
rect 76524 69188 76580 69246
rect 76860 69300 76916 70142
rect 76860 69234 76916 69244
rect 76524 69122 76580 69132
rect 77308 69188 77364 69198
rect 77308 69094 77364 69132
rect 76188 68674 76244 68684
rect 76860 68738 76916 68750
rect 76860 68686 76862 68738
rect 76914 68686 76916 68738
rect 75964 68628 76020 68638
rect 75964 68534 76020 68572
rect 76412 68516 76468 68526
rect 76412 68422 76468 68460
rect 76860 67956 76916 68686
rect 77196 68626 77252 68638
rect 77196 68574 77198 68626
rect 77250 68574 77252 68626
rect 77196 68516 77252 68574
rect 77196 68450 77252 68460
rect 76860 67890 76916 67900
rect 77308 67844 77364 67854
rect 77308 67750 77364 67788
rect 74396 67172 75236 67228
rect 70364 4498 70420 4508
rect 70700 8372 70980 8428
rect 71708 50372 71876 50428
rect 72380 50372 72884 50428
rect 73500 50372 73668 50428
rect 73724 50372 73892 50428
rect 69804 4340 69860 4350
rect 69692 4228 69748 4238
rect 69692 4134 69748 4172
rect 68460 1708 68628 1764
rect 69132 2604 69524 2660
rect 68460 800 68516 1708
rect 69132 800 69188 2604
rect 69804 800 69860 4284
rect 70588 3556 70644 3566
rect 70588 3462 70644 3500
rect 70476 3444 70532 3454
rect 70476 800 70532 3388
rect 70700 3332 70756 8372
rect 71036 4898 71092 4910
rect 71036 4846 71038 4898
rect 71090 4846 71092 4898
rect 70812 4340 70868 4350
rect 71036 4340 71092 4846
rect 71596 4898 71652 4910
rect 71596 4846 71598 4898
rect 71650 4846 71652 4898
rect 71148 4564 71204 4574
rect 71148 4470 71204 4508
rect 71260 4452 71316 4462
rect 70868 4284 71092 4340
rect 71148 4340 71204 4350
rect 70812 4246 70868 4284
rect 70700 3266 70756 3276
rect 71148 800 71204 4284
rect 71260 3668 71316 4396
rect 71260 3554 71316 3612
rect 71260 3502 71262 3554
rect 71314 3502 71316 3554
rect 71260 3490 71316 3502
rect 71596 4340 71652 4846
rect 71708 4562 71764 50372
rect 72044 5012 72100 5022
rect 71708 4510 71710 4562
rect 71762 4510 71764 4562
rect 71708 4498 71764 4510
rect 71932 5010 72100 5012
rect 71932 4958 72046 5010
rect 72098 4958 72100 5010
rect 71932 4956 72100 4958
rect 71932 4340 71988 4956
rect 72044 4946 72100 4956
rect 72380 5010 72436 50372
rect 72380 4958 72382 5010
rect 72434 4958 72436 5010
rect 72380 4946 72436 4958
rect 72828 4900 72884 4910
rect 72716 4898 72884 4900
rect 72716 4846 72830 4898
rect 72882 4846 72884 4898
rect 72716 4844 72884 4846
rect 71596 4284 71988 4340
rect 72044 4340 72100 4350
rect 71596 3332 71652 4284
rect 72044 4246 72100 4284
rect 72492 4340 72548 4350
rect 72492 4246 72548 4284
rect 72716 3444 72772 4844
rect 72828 4834 72884 4844
rect 73388 4898 73444 4910
rect 73388 4846 73390 4898
rect 73442 4846 73444 4898
rect 73388 4338 73444 4846
rect 73500 4564 73556 50372
rect 73500 4498 73556 4508
rect 73724 4562 73780 50372
rect 75068 48244 75124 48254
rect 74620 48242 75124 48244
rect 74620 48190 75070 48242
rect 75122 48190 75124 48242
rect 74620 48188 75124 48190
rect 74620 48130 74676 48188
rect 75068 48178 75124 48188
rect 74620 48078 74622 48130
rect 74674 48078 74676 48130
rect 74620 47236 74676 48078
rect 74620 47170 74676 47180
rect 75068 46676 75124 46686
rect 74620 46674 75124 46676
rect 74620 46622 75070 46674
rect 75122 46622 75124 46674
rect 74620 46620 75124 46622
rect 74620 46562 74676 46620
rect 75068 46610 75124 46620
rect 74620 46510 74622 46562
rect 74674 46510 74676 46562
rect 74620 45780 74676 46510
rect 74620 45714 74676 45724
rect 74732 45668 74788 45678
rect 74732 45574 74788 45612
rect 75068 45108 75124 45118
rect 74620 45106 75124 45108
rect 74620 45054 75070 45106
rect 75122 45054 75124 45106
rect 74620 45052 75124 45054
rect 74620 44994 74676 45052
rect 75068 45042 75124 45052
rect 74620 44942 74622 44994
rect 74674 44942 74676 44994
rect 74620 44212 74676 44942
rect 74620 44146 74676 44156
rect 75068 41972 75124 41982
rect 74620 41970 75124 41972
rect 74620 41918 75070 41970
rect 75122 41918 75124 41970
rect 74620 41916 75124 41918
rect 74620 41858 74676 41916
rect 75068 41906 75124 41916
rect 74620 41806 74622 41858
rect 74674 41806 74676 41858
rect 74620 41076 74676 41806
rect 74620 41010 74676 41020
rect 74620 40404 74676 40414
rect 75068 40404 75124 40414
rect 74620 40402 75124 40404
rect 74620 40350 74622 40402
rect 74674 40350 75070 40402
rect 75122 40350 75124 40402
rect 74620 40348 75124 40350
rect 74620 39508 74676 40348
rect 75068 40338 75124 40348
rect 74620 39442 74676 39452
rect 74732 39394 74788 39406
rect 74732 39342 74734 39394
rect 74786 39342 74788 39394
rect 74732 39060 74788 39342
rect 74732 38994 74788 39004
rect 75068 38836 75124 38846
rect 74620 38834 75124 38836
rect 74620 38782 75070 38834
rect 75122 38782 75124 38834
rect 74620 38780 75124 38782
rect 74620 38722 74676 38780
rect 75068 38770 75124 38780
rect 74620 38670 74622 38722
rect 74674 38670 74676 38722
rect 74620 37828 74676 38670
rect 74620 37762 74676 37772
rect 75068 37268 75124 37278
rect 74620 37266 75124 37268
rect 74620 37214 75070 37266
rect 75122 37214 75124 37266
rect 74620 37212 75124 37214
rect 74620 37154 74676 37212
rect 75068 37202 75124 37212
rect 74620 37102 74622 37154
rect 74674 37102 74676 37154
rect 74620 36260 74676 37102
rect 74620 36194 74676 36204
rect 75068 35700 75124 35710
rect 74620 35698 75124 35700
rect 74620 35646 75070 35698
rect 75122 35646 75124 35698
rect 74620 35644 75124 35646
rect 74620 35586 74676 35644
rect 75068 35634 75124 35644
rect 74620 35534 74622 35586
rect 74674 35534 74676 35586
rect 74620 34804 74676 35534
rect 74620 34738 74676 34748
rect 74732 34690 74788 34702
rect 74732 34638 74734 34690
rect 74786 34638 74788 34690
rect 74732 34356 74788 34638
rect 74732 34290 74788 34300
rect 75068 34132 75124 34142
rect 74620 34130 75124 34132
rect 74620 34078 75070 34130
rect 75122 34078 75124 34130
rect 74620 34076 75124 34078
rect 74620 34018 74676 34076
rect 75068 34066 75124 34076
rect 74620 33966 74622 34018
rect 74674 33966 74676 34018
rect 74620 33124 74676 33966
rect 74620 33058 74676 33068
rect 74620 32564 74676 32574
rect 75068 32564 75124 32574
rect 74620 32562 75124 32564
rect 74620 32510 74622 32562
rect 74674 32510 75070 32562
rect 75122 32510 75124 32562
rect 74620 32508 75124 32510
rect 74620 31556 74676 32508
rect 75068 32498 75124 32508
rect 74620 31490 74676 31500
rect 75068 30996 75124 31006
rect 74620 30994 75124 30996
rect 74620 30942 75070 30994
rect 75122 30942 75124 30994
rect 74620 30940 75124 30942
rect 74620 30882 74676 30940
rect 75068 30930 75124 30940
rect 74620 30830 74622 30882
rect 74674 30830 74676 30882
rect 74620 30100 74676 30830
rect 74620 30034 74676 30044
rect 74732 29986 74788 29998
rect 74732 29934 74734 29986
rect 74786 29934 74788 29986
rect 74732 29652 74788 29934
rect 74732 29586 74788 29596
rect 75068 29428 75124 29438
rect 74620 29426 75124 29428
rect 74620 29374 75070 29426
rect 75122 29374 75124 29426
rect 74620 29372 75124 29374
rect 74620 29314 74676 29372
rect 75068 29362 75124 29372
rect 74620 29262 74622 29314
rect 74674 29262 74676 29314
rect 74620 28420 74676 29262
rect 74620 28354 74676 28364
rect 75068 27860 75124 27870
rect 74620 27858 75124 27860
rect 74620 27806 75070 27858
rect 75122 27806 75124 27858
rect 74620 27804 75124 27806
rect 74620 27746 74676 27804
rect 75068 27794 75124 27804
rect 74620 27694 74622 27746
rect 74674 27694 74676 27746
rect 74620 26852 74676 27694
rect 74620 26786 74676 26796
rect 75068 26290 75124 26302
rect 75068 26238 75070 26290
rect 75122 26238 75124 26290
rect 74620 26180 74676 26190
rect 75068 26180 75124 26238
rect 74620 26178 75124 26180
rect 74620 26126 74622 26178
rect 74674 26126 75124 26178
rect 74620 26124 75124 26126
rect 74620 25284 74676 26124
rect 74620 25218 74676 25228
rect 74732 25282 74788 25294
rect 74732 25230 74734 25282
rect 74786 25230 74788 25282
rect 74732 25172 74788 25230
rect 74732 24836 74788 25116
rect 74508 24780 74788 24836
rect 74508 23716 74564 24780
rect 75068 24724 75124 24734
rect 74620 24722 75124 24724
rect 74620 24670 75070 24722
rect 75122 24670 75124 24722
rect 74620 24668 75124 24670
rect 74620 24610 74676 24668
rect 75068 24658 75124 24668
rect 74620 24558 74622 24610
rect 74674 24558 74676 24610
rect 74620 23828 74676 24558
rect 74620 23762 74676 23772
rect 74508 23650 74564 23660
rect 75068 23156 75124 23166
rect 74620 23154 75124 23156
rect 74620 23102 75070 23154
rect 75122 23102 75124 23154
rect 74620 23100 75124 23102
rect 74620 23042 74676 23100
rect 75068 23090 75124 23100
rect 74620 22990 74622 23042
rect 74674 22990 74676 23042
rect 74620 22148 74676 22990
rect 74620 22082 74676 22092
rect 75068 21588 75124 21598
rect 74620 21586 75124 21588
rect 74620 21534 75070 21586
rect 75122 21534 75124 21586
rect 74620 21532 75124 21534
rect 74620 21476 74676 21532
rect 75068 21522 75124 21532
rect 74508 21474 74676 21476
rect 74508 21422 74622 21474
rect 74674 21422 74676 21474
rect 74508 21420 74676 21422
rect 74508 20580 74564 21420
rect 74620 21410 74676 21420
rect 74732 20580 74788 20590
rect 74508 20514 74564 20524
rect 74620 20578 74788 20580
rect 74620 20526 74734 20578
rect 74786 20526 74788 20578
rect 74620 20524 74788 20526
rect 74620 20188 74676 20524
rect 74732 20514 74788 20524
rect 74508 20132 74676 20188
rect 74508 19012 74564 20076
rect 75068 20020 75124 20030
rect 74620 20018 75124 20020
rect 74620 19966 75070 20018
rect 75122 19966 75124 20018
rect 74620 19964 75124 19966
rect 74620 19906 74676 19964
rect 75068 19954 75124 19964
rect 74620 19854 74622 19906
rect 74674 19854 74676 19906
rect 74620 19124 74676 19854
rect 74620 19058 74676 19068
rect 74508 18946 74564 18956
rect 75068 18452 75124 18462
rect 74620 18450 75124 18452
rect 74620 18398 75070 18450
rect 75122 18398 75124 18450
rect 74620 18396 75124 18398
rect 74620 18338 74676 18396
rect 75068 18386 75124 18396
rect 74620 18286 74622 18338
rect 74674 18286 74676 18338
rect 74620 17892 74676 18286
rect 74620 17826 74676 17836
rect 74508 17780 74564 17790
rect 74508 17108 74564 17724
rect 74620 17108 74676 17118
rect 74508 17106 74676 17108
rect 74508 17054 74622 17106
rect 74674 17054 74676 17106
rect 74508 17052 74676 17054
rect 74620 16884 74676 17052
rect 75068 16884 75124 16894
rect 74620 16882 75124 16884
rect 74620 16830 75070 16882
rect 75122 16830 75124 16882
rect 74620 16828 75124 16830
rect 75068 16818 75124 16828
rect 74732 16100 74788 16110
rect 74732 15874 74788 16044
rect 74732 15822 74734 15874
rect 74786 15822 74788 15874
rect 74732 15428 74788 15822
rect 74732 15362 74788 15372
rect 75068 15314 75124 15326
rect 75068 15262 75070 15314
rect 75122 15262 75124 15314
rect 74620 15204 74676 15214
rect 74620 15110 74676 15148
rect 75068 15204 75124 15262
rect 75068 15138 75124 15148
rect 74620 13748 74676 13758
rect 74620 13654 74676 13692
rect 75068 13748 75124 13758
rect 75068 13654 75124 13692
rect 75068 12180 75124 12190
rect 74620 12178 75124 12180
rect 74620 12126 75070 12178
rect 75122 12126 75124 12178
rect 74620 12124 75124 12126
rect 74620 12066 74676 12124
rect 75068 12114 75124 12124
rect 74620 12014 74622 12066
rect 74674 12014 74676 12066
rect 74620 11284 74676 12014
rect 74620 11218 74676 11228
rect 74732 11170 74788 11182
rect 74732 11118 74734 11170
rect 74786 11118 74788 11170
rect 74732 10836 74788 11118
rect 74732 10770 74788 10780
rect 75068 10612 75124 10622
rect 74620 10610 75124 10612
rect 74620 10558 75070 10610
rect 75122 10558 75124 10610
rect 74620 10556 75124 10558
rect 74620 10498 74676 10556
rect 75068 10546 75124 10556
rect 74620 10446 74622 10498
rect 74674 10446 74676 10498
rect 74620 9604 74676 10446
rect 74620 9538 74676 9548
rect 74620 9044 74676 9054
rect 75068 9044 75124 9054
rect 74620 9042 75124 9044
rect 74620 8990 74622 9042
rect 74674 8990 75070 9042
rect 75122 8990 75124 9042
rect 74620 8988 75124 8990
rect 74620 8036 74676 8988
rect 75068 8978 75124 8988
rect 74620 7970 74676 7980
rect 75068 7476 75124 7486
rect 74620 7474 75124 7476
rect 74620 7422 75070 7474
rect 75122 7422 75124 7474
rect 74620 7420 75124 7422
rect 74620 7362 74676 7420
rect 75068 7410 75124 7420
rect 74620 7310 74622 7362
rect 74674 7310 74676 7362
rect 74620 6580 74676 7310
rect 74620 6514 74676 6524
rect 74732 6692 74788 6702
rect 74732 6466 74788 6636
rect 74732 6414 74734 6466
rect 74786 6414 74788 6466
rect 74732 6020 74788 6414
rect 74732 5954 74788 5964
rect 75068 5906 75124 5918
rect 75068 5854 75070 5906
rect 75122 5854 75124 5906
rect 74620 5796 74676 5806
rect 75068 5796 75124 5854
rect 74620 5794 75124 5796
rect 74620 5742 74622 5794
rect 74674 5742 75124 5794
rect 74620 5740 75124 5742
rect 74396 5460 74452 5470
rect 74396 5234 74452 5404
rect 74396 5182 74398 5234
rect 74450 5182 74452 5234
rect 73724 4510 73726 4562
rect 73778 4510 73780 4562
rect 73724 4498 73780 4510
rect 74060 4898 74116 4910
rect 74060 4846 74062 4898
rect 74114 4846 74116 4898
rect 73388 4286 73390 4338
rect 73442 4286 73444 4338
rect 73164 3668 73220 3678
rect 73164 3574 73220 3612
rect 72716 3350 72772 3388
rect 72380 3332 72436 3342
rect 71596 3276 71876 3332
rect 71820 800 71876 3276
rect 72380 3238 72436 3276
rect 73388 2996 73444 4286
rect 72492 2940 73444 2996
rect 73500 4340 73556 4350
rect 72492 800 72548 2940
rect 73500 2884 73556 4284
rect 74060 4340 74116 4846
rect 74284 4564 74340 4574
rect 74284 4470 74340 4508
rect 74060 4274 74116 4284
rect 74284 3556 74340 3566
rect 74396 3556 74452 5182
rect 74620 4900 74676 5740
rect 74620 4834 74676 4844
rect 74956 4898 75012 4910
rect 74956 4846 74958 4898
rect 75010 4846 75012 4898
rect 74508 4340 74564 4350
rect 74956 4340 75012 4846
rect 75180 4562 75236 67172
rect 77308 67060 77364 67070
rect 77308 66966 77364 67004
rect 77308 66052 77364 66062
rect 77308 65958 77364 65996
rect 77308 65380 77364 65390
rect 77308 65286 77364 65324
rect 76636 64596 76692 64606
rect 76636 64502 76692 64540
rect 77308 64482 77364 64494
rect 77308 64430 77310 64482
rect 77362 64430 77364 64482
rect 76860 64260 76916 64270
rect 76860 64146 76916 64204
rect 77308 64260 77364 64430
rect 77308 64194 77364 64204
rect 76860 64094 76862 64146
rect 76914 64094 76916 64146
rect 76860 64082 76916 64094
rect 77420 64036 77476 64046
rect 76412 63924 76468 63934
rect 76412 63830 76468 63868
rect 77196 63924 77252 63934
rect 77196 63830 77252 63868
rect 77308 63028 77364 63038
rect 77308 62934 77364 62972
rect 77308 62244 77364 62254
rect 77308 62150 77364 62188
rect 77420 61572 77476 63980
rect 77420 61506 77476 61516
rect 77308 61460 77364 61470
rect 77308 61366 77364 61404
rect 77308 60676 77364 60686
rect 77308 60582 77364 60620
rect 76636 59780 76692 59790
rect 76636 59686 76692 59724
rect 77308 59778 77364 59790
rect 77308 59726 77310 59778
rect 77362 59726 77364 59778
rect 76860 59330 76916 59342
rect 76860 59278 76862 59330
rect 76914 59278 76916 59330
rect 76412 59108 76468 59118
rect 76412 59014 76468 59052
rect 76860 58436 76916 59278
rect 77196 59218 77252 59230
rect 77196 59166 77198 59218
rect 77250 59166 77252 59218
rect 77196 59108 77252 59166
rect 77308 59220 77364 59726
rect 77308 59154 77364 59164
rect 77196 59042 77252 59052
rect 76860 58370 76916 58380
rect 77308 58324 77364 58334
rect 77308 58230 77364 58268
rect 77308 57540 77364 57550
rect 77308 57446 77364 57484
rect 77308 56644 77364 56654
rect 77308 56550 77364 56588
rect 77308 55972 77364 55982
rect 77308 55878 77364 55916
rect 77532 55468 77588 73836
rect 77756 73826 77812 73836
rect 77868 73444 77924 74734
rect 78092 74004 78148 74014
rect 78092 73910 78148 73948
rect 77868 73378 77924 73388
rect 77868 73218 77924 73230
rect 77868 73166 77870 73218
rect 77922 73166 77924 73218
rect 77868 71876 77924 73166
rect 77868 71810 77924 71820
rect 77868 71650 77924 71662
rect 77868 71598 77870 71650
rect 77922 71598 77924 71650
rect 77868 70644 77924 71598
rect 77868 70578 77924 70588
rect 78204 70754 78260 70766
rect 78204 70702 78206 70754
rect 78258 70702 78260 70754
rect 77868 70082 77924 70094
rect 77868 70030 77870 70082
rect 77922 70030 77924 70082
rect 77868 69860 77924 70030
rect 77868 69794 77924 69804
rect 78092 69300 78148 69310
rect 78204 69300 78260 70702
rect 78092 69298 78260 69300
rect 78092 69246 78094 69298
rect 78146 69246 78260 69298
rect 78092 69244 78260 69246
rect 78092 69234 78148 69244
rect 77756 69188 77812 69198
rect 77756 69186 77924 69188
rect 77756 69134 77758 69186
rect 77810 69134 77924 69186
rect 77756 69132 77924 69134
rect 77756 69122 77812 69132
rect 77756 68740 77812 68750
rect 77644 68738 77812 68740
rect 77644 68686 77758 68738
rect 77810 68686 77812 68738
rect 77644 68684 77812 68686
rect 77644 66948 77700 68684
rect 77756 68674 77812 68684
rect 77868 68068 77924 69132
rect 77980 68628 78036 68638
rect 78036 68572 78148 68628
rect 77980 68534 78036 68572
rect 77868 68002 77924 68012
rect 77980 67844 78036 67854
rect 77756 67620 77812 67630
rect 77756 67618 77924 67620
rect 77756 67566 77758 67618
rect 77810 67566 77924 67618
rect 77756 67564 77924 67566
rect 77756 67554 77812 67564
rect 77644 66882 77700 66892
rect 77756 67170 77812 67182
rect 77756 67118 77758 67170
rect 77810 67118 77812 67170
rect 77756 66276 77812 67118
rect 77868 67172 77924 67564
rect 77868 67106 77924 67116
rect 77980 66500 78036 67788
rect 78092 67396 78148 68572
rect 78204 67844 78260 69244
rect 78204 67778 78260 67788
rect 78092 67330 78148 67340
rect 78092 67060 78148 67070
rect 78148 67004 78260 67060
rect 78092 66928 78148 67004
rect 77980 66434 78036 66444
rect 77756 66210 77812 66220
rect 78092 66162 78148 66174
rect 78092 66110 78094 66162
rect 78146 66110 78148 66162
rect 77756 66050 77812 66062
rect 77756 65998 77758 66050
rect 77810 65998 77812 66050
rect 77756 65828 77812 65998
rect 77756 65762 77812 65772
rect 78092 66052 78148 66110
rect 77756 65602 77812 65614
rect 77756 65550 77758 65602
rect 77810 65550 77812 65602
rect 77756 64708 77812 65550
rect 77756 64642 77812 64652
rect 77980 65490 78036 65502
rect 77980 65438 77982 65490
rect 78034 65438 78036 65490
rect 77980 65380 78036 65438
rect 77756 64484 77812 64494
rect 77644 64482 77812 64484
rect 77644 64430 77758 64482
rect 77810 64430 77812 64482
rect 77644 64428 77812 64430
rect 77644 62580 77700 64428
rect 77756 64418 77812 64428
rect 77980 64484 78036 65324
rect 78092 65156 78148 65996
rect 78204 65828 78260 67004
rect 78204 65762 78260 65772
rect 78092 65090 78148 65100
rect 77980 64418 78036 64428
rect 78092 64596 78148 64606
rect 77980 64260 78036 64270
rect 77756 64036 77812 64046
rect 77756 63942 77812 63980
rect 77980 63922 78036 64204
rect 77980 63870 77982 63922
rect 78034 63870 78036 63922
rect 77756 62916 77812 62926
rect 77756 62914 77924 62916
rect 77756 62862 77758 62914
rect 77810 62862 77924 62914
rect 77756 62860 77924 62862
rect 77756 62850 77812 62860
rect 77644 62514 77700 62524
rect 77756 62468 77812 62478
rect 77756 62374 77812 62412
rect 77756 61348 77812 61358
rect 77644 61346 77812 61348
rect 77644 61294 77758 61346
rect 77810 61294 77812 61346
rect 77644 61292 77812 61294
rect 77644 60116 77700 61292
rect 77756 61282 77812 61292
rect 77868 61348 77924 62860
rect 77980 62580 78036 63870
rect 78092 63252 78148 64540
rect 78092 63186 78148 63196
rect 77980 62514 78036 62524
rect 78092 63028 78148 63038
rect 77868 61282 77924 61292
rect 77980 62354 78036 62366
rect 77980 62302 77982 62354
rect 78034 62302 78036 62354
rect 77980 62244 78036 62302
rect 77980 61124 78036 62188
rect 78092 61796 78148 62972
rect 78092 61730 78148 61740
rect 78092 61460 78148 61470
rect 78148 61404 78260 61460
rect 78092 61328 78148 61404
rect 77980 61058 78036 61068
rect 77756 60898 77812 60910
rect 77756 60846 77758 60898
rect 77810 60846 77812 60898
rect 77756 60228 77812 60846
rect 77756 60162 77812 60172
rect 78092 60786 78148 60798
rect 78092 60734 78094 60786
rect 78146 60734 78148 60786
rect 78092 60676 78148 60734
rect 77644 60050 77700 60060
rect 77980 60002 78036 60014
rect 77980 59950 77982 60002
rect 78034 59950 78036 60002
rect 77756 59780 77812 59790
rect 77644 59778 77812 59780
rect 77644 59726 77758 59778
rect 77810 59726 77812 59778
rect 77644 59724 77812 59726
rect 77644 58548 77700 59724
rect 77756 59714 77812 59724
rect 77980 59780 78036 59950
rect 78092 59892 78148 60620
rect 78204 60564 78260 61404
rect 78204 60498 78260 60508
rect 78092 59826 78148 59836
rect 77756 59332 77812 59342
rect 77756 59330 77924 59332
rect 77756 59278 77758 59330
rect 77810 59278 77924 59330
rect 77756 59276 77924 59278
rect 77756 59266 77812 59276
rect 77644 58482 77700 58492
rect 77756 58212 77812 58222
rect 77756 58118 77812 58156
rect 77756 57764 77812 57774
rect 77644 57762 77812 57764
rect 77644 57710 77758 57762
rect 77810 57710 77812 57762
rect 77644 57708 77812 57710
rect 77644 56084 77700 57708
rect 77756 57698 77812 57708
rect 77868 57652 77924 59276
rect 77980 58884 78036 59724
rect 77980 58818 78036 58828
rect 78092 59220 78148 59230
rect 77868 57586 77924 57596
rect 77980 58434 78036 58446
rect 77980 58382 77982 58434
rect 78034 58382 78036 58434
rect 77980 58324 78036 58382
rect 77980 57316 78036 58268
rect 78092 57876 78148 59164
rect 78092 57810 78148 57820
rect 77980 57250 78036 57260
rect 78092 57650 78148 57662
rect 78092 57598 78094 57650
rect 78146 57598 78148 57650
rect 78092 57540 78148 57598
rect 77980 56866 78036 56878
rect 77980 56814 77982 56866
rect 78034 56814 78036 56866
rect 77756 56644 77812 56654
rect 77980 56644 78036 56814
rect 77756 56642 77924 56644
rect 77756 56590 77758 56642
rect 77810 56590 77924 56642
rect 77756 56588 77924 56590
rect 77756 56578 77812 56588
rect 77756 56196 77812 56206
rect 77756 56102 77812 56140
rect 77644 56018 77700 56028
rect 77420 55412 77588 55468
rect 76636 55076 76692 55086
rect 76636 54982 76692 55020
rect 77308 55074 77364 55086
rect 77308 55022 77310 55074
rect 77362 55022 77364 55074
rect 76860 54740 76916 54750
rect 76860 54646 76916 54684
rect 77196 54514 77252 54526
rect 77196 54462 77198 54514
rect 77250 54462 77252 54514
rect 76412 54404 76468 54414
rect 76412 54310 76468 54348
rect 77196 54404 77252 54462
rect 77308 54516 77364 55022
rect 77308 54450 77364 54460
rect 77196 54338 77252 54348
rect 77308 53508 77364 53518
rect 77308 53414 77364 53452
rect 77308 52836 77364 52846
rect 77308 52742 77364 52780
rect 77308 51940 77364 51950
rect 77308 51846 77364 51884
rect 77308 51268 77364 51278
rect 77308 51174 77364 51212
rect 77420 50820 77476 55412
rect 77756 55076 77812 55086
rect 77644 55074 77812 55076
rect 77644 55022 77758 55074
rect 77810 55022 77812 55074
rect 77644 55020 77812 55022
rect 77644 53732 77700 55020
rect 77756 55010 77812 55020
rect 77868 54852 77924 56588
rect 77980 55748 78036 56588
rect 78092 56420 78148 57484
rect 78092 56354 78148 56364
rect 77980 55682 78036 55692
rect 78092 56082 78148 56094
rect 78092 56030 78094 56082
rect 78146 56030 78148 56082
rect 78092 55972 78148 56030
rect 78092 55524 78148 55916
rect 78092 55458 78148 55468
rect 77868 54786 77924 54796
rect 77980 55298 78036 55310
rect 77980 55246 77982 55298
rect 78034 55246 78036 55298
rect 77980 55076 78036 55246
rect 77756 54628 77812 54638
rect 77756 54534 77812 54572
rect 77980 53844 78036 55020
rect 78092 54516 78148 54526
rect 78148 54460 78260 54516
rect 78092 54384 78148 54460
rect 77980 53778 78036 53788
rect 77644 53666 77700 53676
rect 78092 53618 78148 53630
rect 78092 53566 78094 53618
rect 78146 53566 78148 53618
rect 77756 53508 77812 53518
rect 77644 53506 77812 53508
rect 77644 53454 77758 53506
rect 77810 53454 77812 53506
rect 77644 53452 77812 53454
rect 77644 52276 77700 53452
rect 77756 53442 77812 53452
rect 78092 53508 78148 53566
rect 77644 52210 77700 52220
rect 77756 53058 77812 53070
rect 77756 53006 77758 53058
rect 77810 53006 77812 53058
rect 77756 52164 77812 53006
rect 77756 52098 77812 52108
rect 77980 52946 78036 52958
rect 77980 52894 77982 52946
rect 78034 52894 78036 52946
rect 77980 52836 78036 52894
rect 77756 51940 77812 51950
rect 77420 50754 77476 50764
rect 77644 51938 77812 51940
rect 77644 51886 77758 51938
rect 77810 51886 77812 51938
rect 77644 51884 77812 51886
rect 77308 50708 77364 50718
rect 77308 50614 77364 50652
rect 77644 50596 77700 51884
rect 77756 51874 77812 51884
rect 77980 51716 78036 52780
rect 78092 52388 78148 53452
rect 78204 53060 78260 54460
rect 78204 52994 78260 53004
rect 78092 52322 78148 52332
rect 77980 51650 78036 51660
rect 78092 52050 78148 52062
rect 78092 51998 78094 52050
rect 78146 51998 78148 52050
rect 78092 51940 78148 51998
rect 77756 51492 77812 51502
rect 77756 51398 77812 51436
rect 77644 50530 77700 50540
rect 77980 51378 78036 51390
rect 77980 51326 77982 51378
rect 78034 51326 78036 51378
rect 77980 51268 78036 51326
rect 77980 50484 78036 51212
rect 78092 51044 78148 51884
rect 78092 50978 78148 50988
rect 77980 50418 78036 50428
rect 78092 50708 78148 50718
rect 78092 50482 78148 50652
rect 78092 50430 78094 50482
rect 78146 50430 78148 50482
rect 77756 50372 77812 50382
rect 77756 50278 77812 50316
rect 77756 49922 77812 49934
rect 77756 49870 77758 49922
rect 77810 49870 77812 49922
rect 77308 49700 77364 49710
rect 77308 49606 77364 49644
rect 77756 49028 77812 49870
rect 77756 48962 77812 48972
rect 77980 49810 78036 49822
rect 77980 49758 77982 49810
rect 78034 49758 78036 49810
rect 77980 49700 78036 49758
rect 78092 49812 78148 50430
rect 78092 49746 78148 49756
rect 77980 49028 78036 49644
rect 77980 48962 78036 48972
rect 78092 48914 78148 48926
rect 78092 48862 78094 48914
rect 78146 48862 78148 48914
rect 76636 48802 76692 48814
rect 76636 48750 76638 48802
rect 76690 48750 76692 48802
rect 76636 48244 76692 48750
rect 77308 48804 77364 48814
rect 77308 48710 77364 48748
rect 77756 48802 77812 48814
rect 77756 48750 77758 48802
rect 77810 48750 77812 48802
rect 77756 48468 77812 48750
rect 77756 48402 77812 48412
rect 78092 48804 78148 48862
rect 78092 48356 78148 48748
rect 78092 48290 78148 48300
rect 76972 48244 77028 48254
rect 76636 48242 77028 48244
rect 76636 48190 76974 48242
rect 77026 48190 77028 48242
rect 76636 48188 77028 48190
rect 76076 48130 76132 48142
rect 76076 48078 76078 48130
rect 76130 48078 76132 48130
rect 76076 47684 76132 48078
rect 76076 47618 76132 47628
rect 76636 47234 76692 47246
rect 76636 47182 76638 47234
rect 76690 47182 76692 47234
rect 76076 46562 76132 46574
rect 76076 46510 76078 46562
rect 76130 46510 76132 46562
rect 76076 46340 76132 46510
rect 76636 46564 76692 47182
rect 76972 46788 77028 48188
rect 77868 48130 77924 48142
rect 77868 48078 77870 48130
rect 77922 48078 77924 48130
rect 77868 47124 77924 48078
rect 77868 47058 77924 47068
rect 76972 46722 77028 46732
rect 77084 46674 77140 46686
rect 77084 46622 77086 46674
rect 77138 46622 77140 46674
rect 77084 46564 77140 46622
rect 76636 46508 77140 46564
rect 76076 46274 76132 46284
rect 75292 45890 75348 45902
rect 75292 45838 75294 45890
rect 75346 45838 75348 45890
rect 75292 45668 75348 45838
rect 75292 45602 75348 45612
rect 76188 45778 76244 45790
rect 76188 45726 76190 45778
rect 76242 45726 76244 45778
rect 76188 45668 76244 45726
rect 76188 45602 76244 45612
rect 76860 45108 76916 45118
rect 76524 45106 76916 45108
rect 76524 45054 76862 45106
rect 76914 45054 76916 45106
rect 76524 45052 76916 45054
rect 76076 44994 76132 45006
rect 76076 44942 76078 44994
rect 76130 44942 76132 44994
rect 76076 44324 76132 44942
rect 76076 44258 76132 44268
rect 76524 44098 76580 45052
rect 76860 45042 76916 45052
rect 76524 44046 76526 44098
rect 76578 44046 76580 44098
rect 76524 43764 76580 44046
rect 77084 44100 77140 46508
rect 77756 46562 77812 46574
rect 77756 46510 77758 46562
rect 77810 46510 77812 46562
rect 77756 44996 77812 46510
rect 77756 44930 77812 44940
rect 77868 44994 77924 45006
rect 77868 44942 77870 44994
rect 77922 44942 77924 44994
rect 77084 44034 77140 44044
rect 76524 43698 76580 43708
rect 77868 43764 77924 44942
rect 77868 43698 77924 43708
rect 76860 43540 76916 43550
rect 76412 43538 76916 43540
rect 76412 43486 76862 43538
rect 76914 43486 76916 43538
rect 76412 43484 76916 43486
rect 76412 43426 76468 43484
rect 76860 43474 76916 43484
rect 76412 43374 76414 43426
rect 76466 43374 76468 43426
rect 76412 42532 76468 43374
rect 77868 43426 77924 43438
rect 77868 43374 77870 43426
rect 77922 43374 77924 43426
rect 77868 42980 77924 43374
rect 77868 42914 77924 42924
rect 76412 42466 76468 42476
rect 76860 41972 76916 41982
rect 76636 41970 76916 41972
rect 76636 41918 76862 41970
rect 76914 41918 76916 41970
rect 76636 41916 76916 41918
rect 76076 41858 76132 41870
rect 76076 41806 76078 41858
rect 76130 41806 76132 41858
rect 76076 41636 76132 41806
rect 76076 41570 76132 41580
rect 76636 40964 76692 41916
rect 76860 41906 76916 41916
rect 77756 41972 77812 41982
rect 77756 41878 77812 41916
rect 76636 40870 76692 40908
rect 77756 40964 77812 40974
rect 76860 40516 76916 40526
rect 75964 40404 76020 40414
rect 75964 40310 76020 40348
rect 76860 40402 76916 40460
rect 76860 40350 76862 40402
rect 76914 40350 76916 40402
rect 76860 40338 76916 40350
rect 77196 40516 77252 40526
rect 77196 39730 77252 40460
rect 77756 40514 77812 40908
rect 77756 40462 77758 40514
rect 77810 40462 77812 40514
rect 77756 40450 77812 40462
rect 77196 39678 77198 39730
rect 77250 39678 77252 39730
rect 77196 39666 77252 39678
rect 75292 39618 75348 39630
rect 75292 39566 75294 39618
rect 75346 39566 75348 39618
rect 75292 39060 75348 39566
rect 77756 39620 77812 39630
rect 75292 38994 75348 39004
rect 76188 39506 76244 39518
rect 76188 39454 76190 39506
rect 76242 39454 76244 39506
rect 76188 38948 76244 39454
rect 76188 38882 76244 38892
rect 76860 39396 76916 39406
rect 76860 38836 76916 39340
rect 77756 38946 77812 39564
rect 77756 38894 77758 38946
rect 77810 38894 77812 38946
rect 77756 38882 77812 38894
rect 76636 38834 76916 38836
rect 76636 38782 76862 38834
rect 76914 38782 76916 38834
rect 76636 38780 76916 38782
rect 76076 38722 76132 38734
rect 76076 38670 76078 38722
rect 76130 38670 76132 38722
rect 76076 38276 76132 38670
rect 76076 38210 76132 38220
rect 76636 38162 76692 38780
rect 76860 38770 76916 38780
rect 76636 38110 76638 38162
rect 76690 38110 76692 38162
rect 76636 38098 76692 38110
rect 77756 37604 77812 37614
rect 76636 37380 76692 37390
rect 76076 37154 76132 37166
rect 76076 37102 76078 37154
rect 76130 37102 76132 37154
rect 76076 37044 76132 37102
rect 76076 36978 76132 36988
rect 76636 36594 76692 37324
rect 76860 37380 76916 37390
rect 76860 37266 76916 37324
rect 77756 37378 77812 37548
rect 77756 37326 77758 37378
rect 77810 37326 77812 37378
rect 77756 37314 77812 37326
rect 76860 37214 76862 37266
rect 76914 37214 76916 37266
rect 76860 37202 76916 37214
rect 76636 36542 76638 36594
rect 76690 36542 76692 36594
rect 76636 36530 76692 36542
rect 77756 36260 77812 36270
rect 76860 35812 76916 35822
rect 76860 35698 76916 35756
rect 76860 35646 76862 35698
rect 76914 35646 76916 35698
rect 76860 35634 76916 35646
rect 77196 35812 77252 35822
rect 76076 35588 76132 35598
rect 76076 35494 76132 35532
rect 77196 35026 77252 35756
rect 77756 35810 77812 36204
rect 77756 35758 77758 35810
rect 77810 35758 77812 35810
rect 77756 35746 77812 35758
rect 77196 34974 77198 35026
rect 77250 34974 77252 35026
rect 77196 34962 77252 34974
rect 75292 34914 75348 34926
rect 75292 34862 75294 34914
rect 75346 34862 75348 34914
rect 75292 34356 75348 34862
rect 77756 34916 77812 34926
rect 75292 34290 75348 34300
rect 76188 34802 76244 34814
rect 76188 34750 76190 34802
rect 76242 34750 76244 34802
rect 76188 34244 76244 34750
rect 76188 34178 76244 34188
rect 76860 34692 76916 34702
rect 76860 34132 76916 34636
rect 77756 34242 77812 34860
rect 77756 34190 77758 34242
rect 77810 34190 77812 34242
rect 77756 34178 77812 34190
rect 76636 34130 76916 34132
rect 76636 34078 76862 34130
rect 76914 34078 76916 34130
rect 76636 34076 76916 34078
rect 76076 34018 76132 34030
rect 76076 33966 76078 34018
rect 76130 33966 76132 34018
rect 76076 33684 76132 33966
rect 76076 33618 76132 33628
rect 76636 33458 76692 34076
rect 76860 34066 76916 34076
rect 76636 33406 76638 33458
rect 76690 33406 76692 33458
rect 76636 33394 76692 33406
rect 77756 32900 77812 32910
rect 76636 32676 76692 32686
rect 76636 32564 76692 32620
rect 77756 32674 77812 32844
rect 77756 32622 77758 32674
rect 77810 32622 77812 32674
rect 77756 32610 77812 32622
rect 76860 32564 76916 32574
rect 76636 32562 76916 32564
rect 76636 32510 76862 32562
rect 76914 32510 76916 32562
rect 76636 32508 76916 32510
rect 76076 32450 76132 32462
rect 76076 32398 76078 32450
rect 76130 32398 76132 32450
rect 76076 32228 76132 32398
rect 76076 32162 76132 32172
rect 76636 31890 76692 32508
rect 76860 32498 76916 32508
rect 76636 31838 76638 31890
rect 76690 31838 76692 31890
rect 76636 31826 76692 31838
rect 77756 31556 77812 31566
rect 76860 31108 76916 31118
rect 76860 30994 76916 31052
rect 76860 30942 76862 30994
rect 76914 30942 76916 30994
rect 76860 30930 76916 30942
rect 77196 31108 77252 31118
rect 76076 30884 76132 30894
rect 76076 30790 76132 30828
rect 77196 30322 77252 31052
rect 77756 31106 77812 31500
rect 77756 31054 77758 31106
rect 77810 31054 77812 31106
rect 77756 31042 77812 31054
rect 77196 30270 77198 30322
rect 77250 30270 77252 30322
rect 77196 30258 77252 30270
rect 75292 30210 75348 30222
rect 75292 30158 75294 30210
rect 75346 30158 75348 30210
rect 75292 29652 75348 30158
rect 77756 30212 77812 30222
rect 75292 29586 75348 29596
rect 76188 30098 76244 30110
rect 76188 30046 76190 30098
rect 76242 30046 76244 30098
rect 76188 29540 76244 30046
rect 76188 29474 76244 29484
rect 76860 29988 76916 29998
rect 76860 29428 76916 29932
rect 77756 29538 77812 30156
rect 77756 29486 77758 29538
rect 77810 29486 77812 29538
rect 77756 29474 77812 29486
rect 76636 29426 76916 29428
rect 76636 29374 76862 29426
rect 76914 29374 76916 29426
rect 76636 29372 76916 29374
rect 76076 29314 76132 29326
rect 76076 29262 76078 29314
rect 76130 29262 76132 29314
rect 76076 28868 76132 29262
rect 76076 28802 76132 28812
rect 76636 28754 76692 29372
rect 76860 29362 76916 29372
rect 76636 28702 76638 28754
rect 76690 28702 76692 28754
rect 76636 28690 76692 28702
rect 77756 28196 77812 28206
rect 76636 27972 76692 27982
rect 76076 27746 76132 27758
rect 76076 27694 76078 27746
rect 76130 27694 76132 27746
rect 76076 27524 76132 27694
rect 76076 27458 76132 27468
rect 76636 27186 76692 27916
rect 76860 27972 76916 27982
rect 76860 27858 76916 27916
rect 77756 27970 77812 28140
rect 77756 27918 77758 27970
rect 77810 27918 77812 27970
rect 77756 27906 77812 27918
rect 76860 27806 76862 27858
rect 76914 27806 76916 27858
rect 76860 27794 76916 27806
rect 76636 27134 76638 27186
rect 76690 27134 76692 27186
rect 76636 27122 76692 27134
rect 77756 26852 77812 26862
rect 76860 26404 76916 26414
rect 76860 26290 76916 26348
rect 76860 26238 76862 26290
rect 76914 26238 76916 26290
rect 76860 26226 76916 26238
rect 77196 26404 77252 26414
rect 76076 26180 76132 26190
rect 76076 26086 76132 26124
rect 77196 25618 77252 26348
rect 77756 26402 77812 26796
rect 77756 26350 77758 26402
rect 77810 26350 77812 26402
rect 77756 26338 77812 26350
rect 77196 25566 77198 25618
rect 77250 25566 77252 25618
rect 77196 25554 77252 25566
rect 75292 25506 75348 25518
rect 75292 25454 75294 25506
rect 75346 25454 75348 25506
rect 75292 25172 75348 25454
rect 77756 25508 77812 25518
rect 75292 25106 75348 25116
rect 76188 25394 76244 25406
rect 76188 25342 76190 25394
rect 76242 25342 76244 25394
rect 76188 24836 76244 25342
rect 76188 24770 76244 24780
rect 77756 24834 77812 25452
rect 77756 24782 77758 24834
rect 77810 24782 77812 24834
rect 77756 24770 77812 24782
rect 76636 24724 76692 24734
rect 76076 24610 76132 24622
rect 76076 24558 76078 24610
rect 76130 24558 76132 24610
rect 76076 24164 76132 24558
rect 76076 24098 76132 24108
rect 76636 24050 76692 24668
rect 76860 24724 76916 24734
rect 76860 24630 76916 24668
rect 76636 23998 76638 24050
rect 76690 23998 76692 24050
rect 76636 23986 76692 23998
rect 77756 23492 77812 23502
rect 76636 23268 76692 23278
rect 76076 23042 76132 23054
rect 76076 22990 76078 23042
rect 76130 22990 76132 23042
rect 76076 22820 76132 22990
rect 76076 22754 76132 22764
rect 76636 22482 76692 23212
rect 76860 23268 76916 23278
rect 76860 23154 76916 23212
rect 77756 23266 77812 23436
rect 77756 23214 77758 23266
rect 77810 23214 77812 23266
rect 77756 23202 77812 23214
rect 76860 23102 76862 23154
rect 76914 23102 76916 23154
rect 76860 23090 76916 23102
rect 76636 22430 76638 22482
rect 76690 22430 76692 22482
rect 76636 22418 76692 22430
rect 77756 22148 77812 22158
rect 76860 21700 76916 21710
rect 76860 21586 76916 21644
rect 76860 21534 76862 21586
rect 76914 21534 76916 21586
rect 76860 21522 76916 21534
rect 77196 21700 77252 21710
rect 76076 21476 76132 21486
rect 76076 21382 76132 21420
rect 77196 20914 77252 21644
rect 77756 21698 77812 22092
rect 77756 21646 77758 21698
rect 77810 21646 77812 21698
rect 77756 21634 77812 21646
rect 77196 20862 77198 20914
rect 77250 20862 77252 20914
rect 77196 20850 77252 20862
rect 75292 20802 75348 20814
rect 75292 20750 75294 20802
rect 75346 20750 75348 20802
rect 75292 20132 75348 20750
rect 76188 20690 76244 20702
rect 76188 20638 76190 20690
rect 76242 20638 76244 20690
rect 76188 20244 76244 20638
rect 76188 20178 76244 20188
rect 75292 20066 75348 20076
rect 77756 20132 77812 20142
rect 77756 20038 77812 20076
rect 76860 20018 76916 20030
rect 76860 19966 76862 20018
rect 76914 19966 76916 20018
rect 76076 19906 76132 19918
rect 76076 19854 76078 19906
rect 76130 19854 76132 19906
rect 76076 19460 76132 19854
rect 76076 19394 76132 19404
rect 76636 19908 76692 19918
rect 76636 19346 76692 19852
rect 76860 19908 76916 19966
rect 76860 19842 76916 19852
rect 76636 19294 76638 19346
rect 76690 19294 76692 19346
rect 76636 19282 76692 19294
rect 76860 18452 76916 18462
rect 76636 18450 76916 18452
rect 76636 18398 76862 18450
rect 76914 18398 76916 18450
rect 76636 18396 76916 18398
rect 76076 18338 76132 18350
rect 76076 18286 76078 18338
rect 76130 18286 76132 18338
rect 76076 18116 76132 18286
rect 76076 18050 76132 18060
rect 76636 17668 76692 18396
rect 76860 18386 76916 18396
rect 77756 18452 77812 18462
rect 77756 18358 77812 18396
rect 76636 17574 76692 17612
rect 77756 17444 77812 17454
rect 76860 16996 76916 17006
rect 75964 16884 76020 16894
rect 75964 16790 76020 16828
rect 76860 16882 76916 16940
rect 76860 16830 76862 16882
rect 76914 16830 76916 16882
rect 76860 16818 76916 16830
rect 77196 16996 77252 17006
rect 77196 16210 77252 16940
rect 77756 16994 77812 17388
rect 77756 16942 77758 16994
rect 77810 16942 77812 16994
rect 77756 16930 77812 16942
rect 77196 16158 77198 16210
rect 77250 16158 77252 16210
rect 77196 16146 77252 16158
rect 75292 16100 75348 16110
rect 75292 16006 75348 16044
rect 77756 16100 77812 16110
rect 76188 15986 76244 15998
rect 76188 15934 76190 15986
rect 76242 15934 76244 15986
rect 76188 15428 76244 15934
rect 76188 15362 76244 15372
rect 76860 15876 76916 15886
rect 76860 15316 76916 15820
rect 77756 15426 77812 16044
rect 77756 15374 77758 15426
rect 77810 15374 77812 15426
rect 77756 15362 77812 15374
rect 76636 15314 76916 15316
rect 76636 15262 76862 15314
rect 76914 15262 76916 15314
rect 76636 15260 76916 15262
rect 76076 15202 76132 15214
rect 76076 15150 76078 15202
rect 76130 15150 76132 15202
rect 76076 14756 76132 15150
rect 76076 14690 76132 14700
rect 76636 14642 76692 15260
rect 76860 15250 76916 15260
rect 76636 14590 76638 14642
rect 76690 14590 76692 14642
rect 76636 14578 76692 14590
rect 77756 14084 77812 14094
rect 76636 13860 76692 13870
rect 76076 13634 76132 13646
rect 76076 13582 76078 13634
rect 76130 13582 76132 13634
rect 76076 13524 76132 13582
rect 76076 13458 76132 13468
rect 76636 13074 76692 13804
rect 76860 13860 76916 13870
rect 76860 13746 76916 13804
rect 77756 13858 77812 14028
rect 77756 13806 77758 13858
rect 77810 13806 77812 13858
rect 77756 13794 77812 13806
rect 76860 13694 76862 13746
rect 76914 13694 76916 13746
rect 76860 13682 76916 13694
rect 76636 13022 76638 13074
rect 76690 13022 76692 13074
rect 76636 13010 76692 13022
rect 77756 12740 77812 12750
rect 76860 12292 76916 12302
rect 76860 12178 76916 12236
rect 76860 12126 76862 12178
rect 76914 12126 76916 12178
rect 76860 12114 76916 12126
rect 77196 12292 77252 12302
rect 76076 12068 76132 12078
rect 76076 11974 76132 12012
rect 77196 11506 77252 12236
rect 77756 12290 77812 12684
rect 77756 12238 77758 12290
rect 77810 12238 77812 12290
rect 77756 12226 77812 12238
rect 77196 11454 77198 11506
rect 77250 11454 77252 11506
rect 77196 11442 77252 11454
rect 75292 11394 75348 11406
rect 75292 11342 75294 11394
rect 75346 11342 75348 11394
rect 75292 10836 75348 11342
rect 77756 11396 77812 11406
rect 75292 10770 75348 10780
rect 76188 11282 76244 11294
rect 76188 11230 76190 11282
rect 76242 11230 76244 11282
rect 76188 10724 76244 11230
rect 76188 10658 76244 10668
rect 76860 11172 76916 11182
rect 76860 10612 76916 11116
rect 77756 10722 77812 11340
rect 77756 10670 77758 10722
rect 77810 10670 77812 10722
rect 77756 10658 77812 10670
rect 76636 10610 76916 10612
rect 76636 10558 76862 10610
rect 76914 10558 76916 10610
rect 76636 10556 76916 10558
rect 76076 10498 76132 10510
rect 76076 10446 76078 10498
rect 76130 10446 76132 10498
rect 76076 10164 76132 10446
rect 76076 10098 76132 10108
rect 76636 9938 76692 10556
rect 76860 10546 76916 10556
rect 76636 9886 76638 9938
rect 76690 9886 76692 9938
rect 76636 9874 76692 9886
rect 77756 9380 77812 9390
rect 76636 9156 76692 9166
rect 76636 9044 76692 9100
rect 77756 9154 77812 9324
rect 77756 9102 77758 9154
rect 77810 9102 77812 9154
rect 77756 9090 77812 9102
rect 76860 9044 76916 9054
rect 76636 9042 76916 9044
rect 76636 8990 76862 9042
rect 76914 8990 76916 9042
rect 76636 8988 76916 8990
rect 76076 8930 76132 8942
rect 76076 8878 76078 8930
rect 76130 8878 76132 8930
rect 76076 8708 76132 8878
rect 76076 8642 76132 8652
rect 76636 8370 76692 8988
rect 76860 8978 76916 8988
rect 76636 8318 76638 8370
rect 76690 8318 76692 8370
rect 76636 8306 76692 8318
rect 77756 8036 77812 8046
rect 76860 7588 76916 7598
rect 76860 7474 76916 7532
rect 76860 7422 76862 7474
rect 76914 7422 76916 7474
rect 76860 7410 76916 7422
rect 77196 7588 77252 7598
rect 76076 7364 76132 7374
rect 76076 7270 76132 7308
rect 77196 6802 77252 7532
rect 77756 7586 77812 7980
rect 77756 7534 77758 7586
rect 77810 7534 77812 7586
rect 77756 7522 77812 7534
rect 77196 6750 77198 6802
rect 77250 6750 77252 6802
rect 77196 6738 77252 6750
rect 75292 6692 75348 6702
rect 75292 6598 75348 6636
rect 77756 6692 77812 6702
rect 76188 6578 76244 6590
rect 76188 6526 76190 6578
rect 76242 6526 76244 6578
rect 76188 6020 76244 6526
rect 76188 5954 76244 5964
rect 76860 6468 76916 6478
rect 76860 5908 76916 6412
rect 77756 6018 77812 6636
rect 77756 5966 77758 6018
rect 77810 5966 77812 6018
rect 77756 5954 77812 5966
rect 76636 5906 76916 5908
rect 76636 5854 76862 5906
rect 76914 5854 76916 5906
rect 76636 5852 76916 5854
rect 76076 5794 76132 5806
rect 76076 5742 76078 5794
rect 76130 5742 76132 5794
rect 76076 5348 76132 5742
rect 76076 5282 76132 5292
rect 76636 5234 76692 5852
rect 76860 5842 76916 5852
rect 76636 5182 76638 5234
rect 76690 5182 76692 5234
rect 76636 5170 76692 5182
rect 75180 4510 75182 4562
rect 75234 4510 75236 4562
rect 75180 4498 75236 4510
rect 75404 4340 75460 4350
rect 74956 4338 75460 4340
rect 74956 4286 75406 4338
rect 75458 4286 75460 4338
rect 74956 4284 75460 4286
rect 74508 4246 74564 4284
rect 74284 3554 74452 3556
rect 74284 3502 74286 3554
rect 74338 3502 74452 3554
rect 74284 3500 74452 3502
rect 74284 3490 74340 3500
rect 73164 2828 73556 2884
rect 73836 3444 73892 3454
rect 73164 800 73220 2828
rect 73836 800 73892 3388
rect 74956 3444 75012 3454
rect 74956 3350 75012 3388
rect 74508 924 74788 980
rect 74508 800 74564 924
rect 5264 0 5376 800
rect 5936 0 6048 800
rect 6608 0 6720 800
rect 7280 0 7392 800
rect 7952 0 8064 800
rect 8624 0 8736 800
rect 9296 0 9408 800
rect 9968 0 10080 800
rect 10640 0 10752 800
rect 11312 0 11424 800
rect 11984 0 12096 800
rect 12656 0 12768 800
rect 13328 0 13440 800
rect 14000 0 14112 800
rect 14672 0 14784 800
rect 15344 0 15456 800
rect 16016 0 16128 800
rect 16688 0 16800 800
rect 17360 0 17472 800
rect 18032 0 18144 800
rect 18704 0 18816 800
rect 19376 0 19488 800
rect 20048 0 20160 800
rect 20720 0 20832 800
rect 21392 0 21504 800
rect 22064 0 22176 800
rect 22736 0 22848 800
rect 23408 0 23520 800
rect 24080 0 24192 800
rect 24752 0 24864 800
rect 25424 0 25536 800
rect 26096 0 26208 800
rect 26768 0 26880 800
rect 27440 0 27552 800
rect 28112 0 28224 800
rect 28784 0 28896 800
rect 29456 0 29568 800
rect 30128 0 30240 800
rect 30800 0 30912 800
rect 31472 0 31584 800
rect 32144 0 32256 800
rect 32816 0 32928 800
rect 33488 0 33600 800
rect 34160 0 34272 800
rect 34832 0 34944 800
rect 35504 0 35616 800
rect 36176 0 36288 800
rect 36848 0 36960 800
rect 37520 0 37632 800
rect 38192 0 38304 800
rect 38864 0 38976 800
rect 39536 0 39648 800
rect 40208 0 40320 800
rect 40880 0 40992 800
rect 41552 0 41664 800
rect 42224 0 42336 800
rect 42896 0 43008 800
rect 43568 0 43680 800
rect 44240 0 44352 800
rect 44912 0 45024 800
rect 45584 0 45696 800
rect 46256 0 46368 800
rect 46928 0 47040 800
rect 47600 0 47712 800
rect 48272 0 48384 800
rect 48944 0 49056 800
rect 49616 0 49728 800
rect 50288 0 50400 800
rect 50960 0 51072 800
rect 51632 0 51744 800
rect 52304 0 52416 800
rect 52976 0 53088 800
rect 53648 0 53760 800
rect 54320 0 54432 800
rect 54992 0 55104 800
rect 55664 0 55776 800
rect 56336 0 56448 800
rect 57008 0 57120 800
rect 57680 0 57792 800
rect 58352 0 58464 800
rect 59024 0 59136 800
rect 59696 0 59808 800
rect 60368 0 60480 800
rect 61040 0 61152 800
rect 61712 0 61824 800
rect 62384 0 62496 800
rect 63056 0 63168 800
rect 63728 0 63840 800
rect 64400 0 64512 800
rect 65072 0 65184 800
rect 65744 0 65856 800
rect 66416 0 66528 800
rect 67088 0 67200 800
rect 67760 0 67872 800
rect 68432 0 68544 800
rect 69104 0 69216 800
rect 69776 0 69888 800
rect 70448 0 70560 800
rect 71120 0 71232 800
rect 71792 0 71904 800
rect 72464 0 72576 800
rect 73136 0 73248 800
rect 73808 0 73920 800
rect 74480 0 74592 800
rect 74732 756 74788 924
rect 75404 756 75460 4284
rect 74732 700 75460 756
<< via2 >>
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 73724 74844 73780 74900
rect 3052 74732 3108 74788
rect 2044 74508 2100 74564
rect 3052 74114 3108 74116
rect 3052 74062 3054 74114
rect 3054 74062 3106 74114
rect 3106 74062 3108 74114
rect 3052 74060 3108 74062
rect 4060 74786 4116 74788
rect 4060 74734 4062 74786
rect 4062 74734 4114 74786
rect 4114 74734 4116 74786
rect 4060 74732 4116 74734
rect 4844 74732 4900 74788
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 4284 74060 4340 74116
rect 3612 73836 3668 73892
rect 2156 73164 2212 73220
rect 3052 73164 3108 73220
rect 3612 73218 3668 73220
rect 3612 73166 3614 73218
rect 3614 73166 3666 73218
rect 3666 73166 3668 73218
rect 3612 73164 3668 73166
rect 2044 72492 2100 72548
rect 2156 71820 2212 71876
rect 3500 71820 3556 71876
rect 3052 71596 3108 71652
rect 3612 71650 3668 71652
rect 3612 71598 3614 71650
rect 3614 71598 3666 71650
rect 3666 71598 3668 71650
rect 3612 71596 3668 71598
rect 2044 71148 2100 71204
rect 2156 70476 2212 70532
rect 3500 70252 3556 70308
rect 3052 70028 3108 70084
rect 3612 70082 3668 70084
rect 3612 70030 3614 70082
rect 3614 70030 3666 70082
rect 3666 70030 3668 70082
rect 3612 70028 3668 70030
rect 2044 69804 2100 69860
rect 1820 69298 1876 69300
rect 1820 69246 1822 69298
rect 1822 69246 1874 69298
rect 1874 69246 1876 69298
rect 1820 69244 1876 69246
rect 3948 69298 4004 69300
rect 3948 69246 3950 69298
rect 3950 69246 4002 69298
rect 4002 69246 4004 69298
rect 3948 69244 4004 69246
rect 1820 67900 1876 67956
rect 1932 68626 1988 68628
rect 1932 68574 1934 68626
rect 1934 68574 1986 68626
rect 1986 68574 1988 68626
rect 1932 68572 1988 68574
rect 2716 69132 2772 69188
rect 3052 68738 3108 68740
rect 3052 68686 3054 68738
rect 3054 68686 3106 68738
rect 3106 68686 3108 68738
rect 3052 68684 3108 68686
rect 2716 68460 2772 68516
rect 3500 69186 3556 69188
rect 3500 69134 3502 69186
rect 3502 69134 3554 69186
rect 3554 69134 3556 69186
rect 3500 69132 3556 69134
rect 3500 68626 3556 68628
rect 3500 68574 3502 68626
rect 3502 68574 3554 68626
rect 3554 68574 3556 68626
rect 3500 68572 3556 68574
rect 3164 68460 3220 68516
rect 2268 67788 2324 67844
rect 1932 67228 1988 67284
rect 1820 67116 1876 67172
rect 1820 66444 1876 66500
rect 1932 66892 1988 66948
rect 1932 65772 1988 65828
rect 1820 65100 1876 65156
rect 2268 66220 2324 66276
rect 3052 67116 3108 67172
rect 2604 66946 2660 66948
rect 2604 66894 2606 66946
rect 2606 66894 2658 66946
rect 2658 66894 2660 66946
rect 2604 66892 2660 66894
rect 2044 65436 2100 65492
rect 1932 65324 1988 65380
rect 1932 64428 1988 64484
rect 2380 65996 2436 66052
rect 2604 65378 2660 65380
rect 2604 65326 2606 65378
rect 2606 65326 2658 65378
rect 2658 65326 2660 65378
rect 2604 65324 2660 65326
rect 2492 65100 2548 65156
rect 2268 64652 2324 64708
rect 1708 63644 1764 63700
rect 1708 63084 1764 63140
rect 1932 63980 1988 64036
rect 2044 63868 2100 63924
rect 2156 63084 2212 63140
rect 1932 62524 1988 62580
rect 1820 61740 1876 61796
rect 1932 62076 1988 62132
rect 1820 61458 1876 61460
rect 1820 61406 1822 61458
rect 1822 61406 1874 61458
rect 1874 61406 1876 61458
rect 1820 61404 1876 61406
rect 1932 61068 1988 61124
rect 1708 60396 1764 60452
rect 2604 63644 2660 63700
rect 2716 63756 2772 63812
rect 2380 62188 2436 62244
rect 2604 62076 2660 62132
rect 3500 64034 3556 64036
rect 3500 63982 3502 64034
rect 3502 63982 3554 64034
rect 3554 63982 3556 64034
rect 3500 63980 3556 63982
rect 3164 62860 3220 62916
rect 3052 61740 3108 61796
rect 2268 61516 2324 61572
rect 2604 61458 2660 61460
rect 2604 61406 2606 61458
rect 2606 61406 2658 61458
rect 2658 61406 2660 61458
rect 2604 61404 2660 61406
rect 2044 60620 2100 60676
rect 1932 60396 1988 60452
rect 2604 60396 2660 60452
rect 2268 60060 2324 60116
rect 2156 59948 2212 60004
rect 1932 59724 1988 59780
rect 1708 58380 1764 58436
rect 1932 59218 1988 59220
rect 1932 59166 1934 59218
rect 1934 59166 1986 59218
rect 1986 59166 1988 59218
rect 1932 59164 1988 59166
rect 2156 58604 2212 58660
rect 2268 58492 2324 58548
rect 2716 59052 2772 59108
rect 2604 58380 2660 58436
rect 3500 59218 3556 59220
rect 3500 59166 3502 59218
rect 3502 59166 3554 59218
rect 3554 59166 3556 59218
rect 3500 59164 3556 59166
rect 3052 58380 3108 58436
rect 3276 58604 3332 58660
rect 1932 57820 1988 57876
rect 1820 57036 1876 57092
rect 1932 56924 1988 56980
rect 1820 56588 1876 56644
rect 1932 56364 1988 56420
rect 1820 55692 1876 55748
rect 2604 56924 2660 56980
rect 3276 57484 3332 57540
rect 3052 57036 3108 57092
rect 2716 56700 2772 56756
rect 2044 55916 2100 55972
rect 1932 55020 1988 55076
rect 2604 56642 2660 56644
rect 2604 56590 2606 56642
rect 2606 56590 2658 56642
rect 2658 56590 2660 56642
rect 2604 56588 2660 56590
rect 2268 55356 2324 55412
rect 2044 54684 2100 54740
rect 1708 53676 1764 53732
rect 1932 54514 1988 54516
rect 1932 54462 1934 54514
rect 1934 54462 1986 54514
rect 1986 54462 1988 54514
rect 1932 54460 1988 54462
rect 1820 53452 1876 53508
rect 2156 53618 2212 53620
rect 2156 53566 2158 53618
rect 2158 53566 2210 53618
rect 2210 53566 2212 53618
rect 2156 53564 2212 53566
rect 2268 53340 2324 53396
rect 1932 53116 1988 53172
rect 2156 53058 2212 53060
rect 2156 53006 2158 53058
rect 2158 53006 2210 53058
rect 2210 53006 2212 53058
rect 2156 53004 2212 53006
rect 2492 55020 2548 55076
rect 3052 54626 3108 54628
rect 3052 54574 3054 54626
rect 3054 54574 3106 54626
rect 3106 54574 3108 54626
rect 3052 54572 3108 54574
rect 3500 54514 3556 54516
rect 3500 54462 3502 54514
rect 3502 54462 3554 54514
rect 3554 54462 3556 54514
rect 3500 54460 3556 54462
rect 2716 54348 2772 54404
rect 2604 53676 2660 53732
rect 3052 53506 3108 53508
rect 3052 53454 3054 53506
rect 3054 53454 3106 53506
rect 3106 53454 3108 53506
rect 3052 53452 3108 53454
rect 1820 52332 1876 52388
rect 1820 52050 1876 52052
rect 1820 51998 1822 52050
rect 1822 51998 1874 52050
rect 1874 51998 1876 52050
rect 1820 51996 1876 51998
rect 2716 52780 2772 52836
rect 2604 52050 2660 52052
rect 2604 51998 2606 52050
rect 2606 51998 2658 52050
rect 2658 51998 2660 52050
rect 2604 51996 2660 51998
rect 2156 51938 2212 51940
rect 2156 51886 2158 51938
rect 2158 51886 2210 51938
rect 2210 51886 2212 51938
rect 2156 51884 2212 51886
rect 1932 51660 1988 51716
rect 1820 50988 1876 51044
rect 1932 50316 1988 50372
rect 1708 50204 1764 50260
rect 2156 49922 2212 49924
rect 2156 49870 2158 49922
rect 2158 49870 2210 49922
rect 2210 49870 2212 49922
rect 2156 49868 2212 49870
rect 1708 48972 1764 49028
rect 1820 49532 1876 49588
rect 1820 48300 1876 48356
rect 2716 49644 2772 49700
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 69356 73442 69412 73444
rect 69356 73390 69358 73442
rect 69358 73390 69410 73442
rect 69410 73390 69412 73442
rect 69356 73388 69412 73390
rect 4844 73052 4900 73108
rect 69132 73276 69188 73332
rect 70028 73330 70084 73332
rect 70028 73278 70030 73330
rect 70030 73278 70082 73330
rect 70082 73278 70084 73330
rect 70028 73276 70084 73278
rect 73276 73276 73332 73332
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 4284 72380 4340 72436
rect 69244 73052 69300 73108
rect 71820 73164 71876 73220
rect 69804 72604 69860 72660
rect 69468 72434 69524 72436
rect 69468 72382 69470 72434
rect 69470 72382 69522 72434
rect 69522 72382 69524 72434
rect 69468 72380 69524 72382
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 67340 68738 67396 68740
rect 67340 68686 67342 68738
rect 67342 68686 67394 68738
rect 67394 68686 67396 68738
rect 67340 68684 67396 68686
rect 67676 68684 67732 68740
rect 66780 68514 66836 68516
rect 66780 68462 66782 68514
rect 66782 68462 66834 68514
rect 66834 68462 66836 68514
rect 66780 68460 66836 68462
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 68684 68738 68740 68740
rect 68684 68686 68686 68738
rect 68686 68686 68738 68738
rect 68738 68686 68740 68738
rect 68684 68684 68740 68686
rect 67788 68514 67844 68516
rect 67788 68462 67790 68514
rect 67790 68462 67842 68514
rect 67842 68462 67844 68514
rect 67788 68460 67844 68462
rect 66668 67842 66724 67844
rect 66668 67790 66670 67842
rect 66670 67790 66722 67842
rect 66722 67790 66724 67842
rect 66668 67788 66724 67790
rect 67116 67842 67172 67844
rect 67116 67790 67118 67842
rect 67118 67790 67170 67842
rect 67170 67790 67172 67842
rect 67116 67788 67172 67790
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 63420 67004 63476 67060
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 63308 66274 63364 66276
rect 63308 66222 63310 66274
rect 63310 66222 63362 66274
rect 63362 66222 63364 66274
rect 63308 66220 63364 66222
rect 63868 66274 63924 66276
rect 63868 66222 63870 66274
rect 63870 66222 63922 66274
rect 63922 66222 63924 66274
rect 63868 66220 63924 66222
rect 64540 66220 64596 66276
rect 61964 66050 62020 66052
rect 61964 65998 61966 66050
rect 61966 65998 62018 66050
rect 62018 65998 62020 66050
rect 61964 65996 62020 65998
rect 62524 66162 62580 66164
rect 62524 66110 62526 66162
rect 62526 66110 62578 66162
rect 62578 66110 62580 66162
rect 62524 66108 62580 66110
rect 62412 65996 62468 66052
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 61852 65548 61908 65604
rect 64876 66274 64932 66276
rect 64876 66222 64878 66274
rect 64878 66222 64930 66274
rect 64930 66222 64932 66274
rect 64876 66220 64932 66222
rect 65996 67058 66052 67060
rect 65996 67006 65998 67058
rect 65998 67006 66050 67058
rect 66050 67006 66052 67058
rect 65996 67004 66052 67006
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 67116 66946 67172 66948
rect 67116 66894 67118 66946
rect 67118 66894 67170 66946
rect 67170 66894 67172 66946
rect 67116 66892 67172 66894
rect 67564 67170 67620 67172
rect 67564 67118 67566 67170
rect 67566 67118 67618 67170
rect 67618 67118 67620 67170
rect 67564 67116 67620 67118
rect 65884 66162 65940 66164
rect 65884 66110 65886 66162
rect 65886 66110 65938 66162
rect 65938 66110 65940 66162
rect 65884 66108 65940 66110
rect 65660 66050 65716 66052
rect 65660 65998 65662 66050
rect 65662 65998 65714 66050
rect 65714 65998 65716 66050
rect 65660 65996 65716 65998
rect 65660 65772 65716 65828
rect 61740 65378 61796 65380
rect 61740 65326 61742 65378
rect 61742 65326 61794 65378
rect 61794 65326 61796 65378
rect 61740 65324 61796 65326
rect 62300 65378 62356 65380
rect 62300 65326 62302 65378
rect 62302 65326 62354 65378
rect 62354 65326 62356 65378
rect 62300 65324 62356 65326
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 65996 65660 66052 65716
rect 66108 65884 66164 65940
rect 67004 66386 67060 66388
rect 67004 66334 67006 66386
rect 67006 66334 67058 66386
rect 67058 66334 67060 66386
rect 67004 66332 67060 66334
rect 67564 66332 67620 66388
rect 67676 67004 67732 67060
rect 66668 65884 66724 65940
rect 66220 65772 66276 65828
rect 66444 65772 66500 65828
rect 65884 65602 65940 65604
rect 65884 65550 65886 65602
rect 65886 65550 65938 65602
rect 65938 65550 65940 65602
rect 65884 65548 65940 65550
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 60732 64706 60788 64708
rect 60732 64654 60734 64706
rect 60734 64654 60786 64706
rect 60786 64654 60788 64706
rect 60732 64652 60788 64654
rect 61404 64706 61460 64708
rect 61404 64654 61406 64706
rect 61406 64654 61458 64706
rect 61458 64654 61460 64706
rect 61404 64652 61460 64654
rect 63532 64706 63588 64708
rect 63532 64654 63534 64706
rect 63534 64654 63586 64706
rect 63586 64654 63588 64706
rect 63532 64652 63588 64654
rect 64204 64706 64260 64708
rect 64204 64654 64206 64706
rect 64206 64654 64258 64706
rect 64258 64654 64260 64706
rect 64204 64652 64260 64654
rect 61516 64482 61572 64484
rect 61516 64430 61518 64482
rect 61518 64430 61570 64482
rect 61570 64430 61572 64482
rect 61516 64428 61572 64430
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 59500 64092 59556 64148
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 59276 62860 59332 62916
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 59388 62748 59444 62804
rect 50764 62692 50820 62694
rect 62188 64092 62244 64148
rect 61180 64034 61236 64036
rect 61180 63982 61182 64034
rect 61182 63982 61234 64034
rect 61234 63982 61236 64034
rect 61180 63980 61236 63982
rect 61068 63922 61124 63924
rect 61068 63870 61070 63922
rect 61070 63870 61122 63922
rect 61122 63870 61124 63922
rect 61068 63868 61124 63870
rect 61628 63922 61684 63924
rect 61628 63870 61630 63922
rect 61630 63870 61682 63922
rect 61682 63870 61684 63922
rect 61628 63868 61684 63870
rect 63420 64034 63476 64036
rect 63420 63982 63422 64034
rect 63422 63982 63474 64034
rect 63474 63982 63476 64034
rect 63420 63980 63476 63982
rect 62524 63756 62580 63812
rect 61404 63138 61460 63140
rect 61404 63086 61406 63138
rect 61406 63086 61458 63138
rect 61458 63086 61460 63138
rect 61404 63084 61460 63086
rect 61964 63138 62020 63140
rect 61964 63086 61966 63138
rect 61966 63086 62018 63138
rect 62018 63086 62020 63138
rect 61964 63084 62020 63086
rect 59836 62914 59892 62916
rect 59836 62862 59838 62914
rect 59838 62862 59890 62914
rect 59890 62862 59892 62914
rect 59836 62860 59892 62862
rect 61516 62524 61572 62580
rect 59836 62354 59892 62356
rect 59836 62302 59838 62354
rect 59838 62302 59890 62354
rect 59890 62302 59892 62354
rect 59836 62300 59892 62302
rect 63532 63868 63588 63924
rect 63308 63196 63364 63252
rect 63420 63756 63476 63812
rect 63644 63810 63700 63812
rect 63644 63758 63646 63810
rect 63646 63758 63698 63810
rect 63698 63758 63700 63810
rect 63644 63756 63700 63758
rect 65100 64316 65156 64372
rect 64540 64204 64596 64260
rect 64876 64204 64932 64260
rect 64428 63922 64484 63924
rect 64428 63870 64430 63922
rect 64430 63870 64482 63922
rect 64482 63870 64484 63922
rect 64428 63868 64484 63870
rect 63980 63756 64036 63812
rect 63196 63084 63252 63140
rect 62636 62578 62692 62580
rect 62636 62526 62638 62578
rect 62638 62526 62690 62578
rect 62690 62526 62692 62578
rect 62636 62524 62692 62526
rect 59724 62242 59780 62244
rect 59724 62190 59726 62242
rect 59726 62190 59778 62242
rect 59778 62190 59780 62242
rect 59724 62188 59780 62190
rect 60284 62242 60340 62244
rect 60284 62190 60286 62242
rect 60286 62190 60338 62242
rect 60338 62190 60340 62242
rect 60284 62188 60340 62190
rect 63644 63084 63700 63140
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 57596 60786 57652 60788
rect 57596 60734 57598 60786
rect 57598 60734 57650 60786
rect 57650 60734 57652 60786
rect 57596 60732 57652 60734
rect 62748 61570 62804 61572
rect 62748 61518 62750 61570
rect 62750 61518 62802 61570
rect 62802 61518 62804 61570
rect 62748 61516 62804 61518
rect 59724 61458 59780 61460
rect 59724 61406 59726 61458
rect 59726 61406 59778 61458
rect 59778 61406 59780 61458
rect 59724 61404 59780 61406
rect 60172 61458 60228 61460
rect 60172 61406 60174 61458
rect 60174 61406 60226 61458
rect 60226 61406 60228 61458
rect 60172 61404 60228 61406
rect 61404 61458 61460 61460
rect 61404 61406 61406 61458
rect 61406 61406 61458 61458
rect 61458 61406 61460 61458
rect 61404 61404 61460 61406
rect 62076 61458 62132 61460
rect 62076 61406 62078 61458
rect 62078 61406 62130 61458
rect 62130 61406 62132 61458
rect 62076 61404 62132 61406
rect 60284 60956 60340 61012
rect 57484 60674 57540 60676
rect 57484 60622 57486 60674
rect 57486 60622 57538 60674
rect 57538 60622 57540 60674
rect 57484 60620 57540 60622
rect 58044 60674 58100 60676
rect 58044 60622 58046 60674
rect 58046 60622 58098 60674
rect 58098 60622 58100 60674
rect 58044 60620 58100 60622
rect 58380 60620 58436 60676
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 57372 60002 57428 60004
rect 57372 59950 57374 60002
rect 57374 59950 57426 60002
rect 57426 59950 57428 60002
rect 57372 59948 57428 59950
rect 57932 60002 57988 60004
rect 57932 59950 57934 60002
rect 57934 59950 57986 60002
rect 57986 59950 57988 60002
rect 57932 59948 57988 59950
rect 57484 59890 57540 59892
rect 57484 59838 57486 59890
rect 57486 59838 57538 59890
rect 57538 59838 57540 59890
rect 57484 59836 57540 59838
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 56140 58434 56196 58436
rect 56140 58382 56142 58434
rect 56142 58382 56194 58434
rect 56194 58382 56196 58434
rect 56140 58380 56196 58382
rect 56700 58434 56756 58436
rect 56700 58382 56702 58434
rect 56702 58382 56754 58434
rect 56754 58382 56756 58434
rect 56700 58380 56756 58382
rect 57260 58322 57316 58324
rect 57260 58270 57262 58322
rect 57262 58270 57314 58322
rect 57314 58270 57316 58322
rect 57260 58268 57316 58270
rect 57820 58322 57876 58324
rect 57820 58270 57822 58322
rect 57822 58270 57874 58322
rect 57874 58270 57876 58322
rect 57820 58268 57876 58270
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 55132 57650 55188 57652
rect 55132 57598 55134 57650
rect 55134 57598 55186 57650
rect 55186 57598 55188 57650
rect 55132 57596 55188 57598
rect 55020 57538 55076 57540
rect 55020 57486 55022 57538
rect 55022 57486 55074 57538
rect 55074 57486 55076 57538
rect 55020 57484 55076 57486
rect 55580 57538 55636 57540
rect 55580 57486 55582 57538
rect 55582 57486 55634 57538
rect 55634 57486 55636 57538
rect 55580 57484 55636 57486
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 57596 57932 57652 57988
rect 57932 57932 57988 57988
rect 57372 57708 57428 57764
rect 57820 57650 57876 57652
rect 57820 57598 57822 57650
rect 57822 57598 57874 57650
rect 57874 57598 57876 57650
rect 57820 57596 57876 57598
rect 56252 56924 56308 56980
rect 56252 56754 56308 56756
rect 56252 56702 56254 56754
rect 56254 56702 56306 56754
rect 56306 56702 56308 56754
rect 56252 56700 56308 56702
rect 56700 56754 56756 56756
rect 56700 56702 56702 56754
rect 56702 56702 56754 56754
rect 56754 56702 56756 56754
rect 56700 56700 56756 56702
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 52220 56082 52276 56084
rect 52220 56030 52222 56082
rect 52222 56030 52274 56082
rect 52274 56030 52276 56082
rect 52220 56028 52276 56030
rect 52108 55970 52164 55972
rect 52108 55918 52110 55970
rect 52110 55918 52162 55970
rect 52162 55918 52164 55970
rect 52108 55916 52164 55918
rect 52668 55970 52724 55972
rect 52668 55918 52670 55970
rect 52670 55918 52722 55970
rect 52722 55918 52724 55970
rect 52668 55916 52724 55918
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 50316 55410 50372 55412
rect 50316 55358 50318 55410
rect 50318 55358 50370 55410
rect 50370 55358 50372 55410
rect 50316 55356 50372 55358
rect 50876 55410 50932 55412
rect 50876 55358 50878 55410
rect 50878 55358 50930 55410
rect 50930 55358 50932 55410
rect 50876 55356 50932 55358
rect 52332 55244 52388 55300
rect 50428 55074 50484 55076
rect 50428 55022 50430 55074
rect 50430 55022 50482 55074
rect 50482 55022 50484 55074
rect 50428 55020 50484 55022
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 51660 54626 51716 54628
rect 51660 54574 51662 54626
rect 51662 54574 51714 54626
rect 51714 54574 51716 54626
rect 51660 54572 51716 54574
rect 52108 54626 52164 54628
rect 52108 54574 52110 54626
rect 52110 54574 52162 54626
rect 52162 54574 52164 54626
rect 52108 54572 52164 54574
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 52220 53676 52276 53732
rect 46956 53564 47012 53620
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 47740 53452 47796 53508
rect 54124 55298 54180 55300
rect 54124 55246 54126 55298
rect 54126 55246 54178 55298
rect 54178 55246 54180 55298
rect 54124 55244 54180 55246
rect 54684 55244 54740 55300
rect 55580 56082 55636 56084
rect 55580 56030 55582 56082
rect 55582 56030 55634 56082
rect 55634 56030 55636 56082
rect 55580 56028 55636 56030
rect 54348 55186 54404 55188
rect 54348 55134 54350 55186
rect 54350 55134 54402 55186
rect 54402 55134 54404 55186
rect 54348 55132 54404 55134
rect 52444 54684 52500 54740
rect 52780 54684 52836 54740
rect 53564 54684 53620 54740
rect 53788 54684 53844 54740
rect 52892 54514 52948 54516
rect 52892 54462 52894 54514
rect 52894 54462 52946 54514
rect 52946 54462 52948 54514
rect 52892 54460 52948 54462
rect 54796 54514 54852 54516
rect 54796 54462 54798 54514
rect 54798 54462 54850 54514
rect 54850 54462 54852 54514
rect 54796 54460 54852 54462
rect 54684 54402 54740 54404
rect 54684 54350 54686 54402
rect 54686 54350 54738 54402
rect 54738 54350 54740 54402
rect 54684 54348 54740 54350
rect 54572 54124 54628 54180
rect 52780 53618 52836 53620
rect 52780 53566 52782 53618
rect 52782 53566 52834 53618
rect 52834 53566 52836 53618
rect 52780 53564 52836 53566
rect 53452 53618 53508 53620
rect 53452 53566 53454 53618
rect 53454 53566 53506 53618
rect 53506 53566 53508 53618
rect 53452 53564 53508 53566
rect 48300 53452 48356 53508
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 48748 53004 48804 53060
rect 48412 52946 48468 52948
rect 48412 52894 48414 52946
rect 48414 52894 48466 52946
rect 48466 52894 48468 52946
rect 48412 52892 48468 52894
rect 46956 52274 47012 52276
rect 46956 52222 46958 52274
rect 46958 52222 47010 52274
rect 47010 52222 47012 52274
rect 46956 52220 47012 52222
rect 47516 52274 47572 52276
rect 47516 52222 47518 52274
rect 47518 52222 47570 52274
rect 47570 52222 47572 52274
rect 47516 52220 47572 52222
rect 50316 53058 50372 53060
rect 50316 53006 50318 53058
rect 50318 53006 50370 53058
rect 50370 53006 50372 53058
rect 50316 53004 50372 53006
rect 52668 53170 52724 53172
rect 52668 53118 52670 53170
rect 52670 53118 52722 53170
rect 52722 53118 52724 53170
rect 52668 53116 52724 53118
rect 53228 53116 53284 53172
rect 50204 52834 50260 52836
rect 50204 52782 50206 52834
rect 50206 52782 50258 52834
rect 50258 52782 50260 52834
rect 50204 52780 50260 52782
rect 50764 52834 50820 52836
rect 50764 52782 50766 52834
rect 50766 52782 50818 52834
rect 50818 52782 50820 52834
rect 50764 52780 50820 52782
rect 48748 52274 48804 52276
rect 48748 52222 48750 52274
rect 48750 52222 48802 52274
rect 48802 52222 48804 52274
rect 48748 52220 48804 52222
rect 52892 52946 52948 52948
rect 52892 52894 52894 52946
rect 52894 52894 52946 52946
rect 52946 52894 52948 52946
rect 52892 52892 52948 52894
rect 51884 52780 51940 52836
rect 52444 52780 52500 52836
rect 52668 52386 52724 52388
rect 52668 52334 52670 52386
rect 52670 52334 52722 52386
rect 52722 52334 52724 52386
rect 52668 52332 52724 52334
rect 49308 52274 49364 52276
rect 49308 52222 49310 52274
rect 49310 52222 49362 52274
rect 49362 52222 49364 52274
rect 49308 52220 49364 52222
rect 47068 52050 47124 52052
rect 47068 51998 47070 52050
rect 47070 51998 47122 52050
rect 47122 51998 47124 52050
rect 47068 51996 47124 51998
rect 52220 52050 52276 52052
rect 52220 51998 52222 52050
rect 52222 51998 52274 52050
rect 52274 51998 52276 52050
rect 52220 51996 52276 51998
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 48860 51548 48916 51604
rect 49196 51884 49252 51940
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 4172 50652 4228 50708
rect 51996 51938 52052 51940
rect 51996 51886 51998 51938
rect 51998 51886 52050 51938
rect 52050 51886 52052 51938
rect 51996 51884 52052 51886
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 52108 51490 52164 51492
rect 52108 51438 52110 51490
rect 52110 51438 52162 51490
rect 52162 51438 52164 51490
rect 52108 51436 52164 51438
rect 49756 50482 49812 50484
rect 49756 50430 49758 50482
rect 49758 50430 49810 50482
rect 49810 50430 49812 50482
rect 49756 50428 49812 50430
rect 50652 50482 50708 50484
rect 50652 50430 50654 50482
rect 50654 50430 50706 50482
rect 50706 50430 50708 50482
rect 50652 50428 50708 50430
rect 51772 50594 51828 50596
rect 51772 50542 51774 50594
rect 51774 50542 51826 50594
rect 51826 50542 51828 50594
rect 51772 50540 51828 50542
rect 3052 50204 3108 50260
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 46620 50034 46676 50036
rect 46620 49982 46622 50034
rect 46622 49982 46674 50034
rect 46674 49982 46676 50034
rect 46620 49980 46676 49982
rect 50540 50370 50596 50372
rect 50540 50318 50542 50370
rect 50542 50318 50594 50370
rect 50594 50318 50596 50370
rect 50540 50316 50596 50318
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 3052 49756 3108 49812
rect 47964 49756 48020 49812
rect 2940 49644 2996 49700
rect 46508 49698 46564 49700
rect 46508 49646 46510 49698
rect 46510 49646 46562 49698
rect 46562 49646 46564 49698
rect 46508 49644 46564 49646
rect 47068 49698 47124 49700
rect 47068 49646 47070 49698
rect 47070 49646 47122 49698
rect 47122 49646 47124 49698
rect 47068 49644 47124 49646
rect 3500 49532 3556 49588
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 49756 49698 49812 49700
rect 49756 49646 49758 49698
rect 49758 49646 49810 49698
rect 49810 49646 49812 49698
rect 49756 49644 49812 49646
rect 49196 49532 49252 49588
rect 48076 49250 48132 49252
rect 48076 49198 48078 49250
rect 48078 49198 48130 49250
rect 48130 49198 48132 49250
rect 48076 49196 48132 49198
rect 47964 49138 48020 49140
rect 47964 49086 47966 49138
rect 47966 49086 48018 49138
rect 48018 49086 48020 49138
rect 47964 49084 48020 49086
rect 48524 49138 48580 49140
rect 48524 49086 48526 49138
rect 48526 49086 48578 49138
rect 48578 49086 48580 49138
rect 48524 49084 48580 49086
rect 3052 48242 3108 48244
rect 3052 48190 3054 48242
rect 3054 48190 3106 48242
rect 3106 48190 3108 48242
rect 3052 48188 3108 48190
rect 2268 48076 2324 48132
rect 48636 48748 48692 48804
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 3612 48188 3668 48244
rect 2156 47628 2212 47684
rect 2044 46956 2100 47012
rect 3052 46674 3108 46676
rect 3052 46622 3054 46674
rect 3054 46622 3106 46674
rect 3106 46622 3108 46674
rect 3052 46620 3108 46622
rect 2156 46284 2212 46340
rect 2044 45612 2100 45668
rect 3612 47180 3668 47236
rect 47292 48130 47348 48132
rect 47292 48078 47294 48130
rect 47294 48078 47346 48130
rect 47346 48078 47348 48130
rect 47292 48076 47348 48078
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 47516 47346 47572 47348
rect 47516 47294 47518 47346
rect 47518 47294 47570 47346
rect 47570 47294 47572 47346
rect 47516 47292 47572 47294
rect 48412 48130 48468 48132
rect 48412 48078 48414 48130
rect 48414 48078 48466 48130
rect 48466 48078 48468 48130
rect 48412 48076 48468 48078
rect 47852 47292 47908 47348
rect 48188 47346 48244 47348
rect 48188 47294 48190 47346
rect 48190 47294 48242 47346
rect 48242 47294 48244 47346
rect 48188 47292 48244 47294
rect 47180 47234 47236 47236
rect 47180 47182 47182 47234
rect 47182 47182 47234 47234
rect 47234 47182 47236 47234
rect 47180 47180 47236 47182
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 3724 46732 3780 46788
rect 46508 46786 46564 46788
rect 46508 46734 46510 46786
rect 46510 46734 46562 46786
rect 46562 46734 46564 46786
rect 46508 46732 46564 46734
rect 47852 46786 47908 46788
rect 47852 46734 47854 46786
rect 47854 46734 47906 46786
rect 47906 46734 47908 46786
rect 47852 46732 47908 46734
rect 3500 45836 3556 45892
rect 3612 46620 3668 46676
rect 3500 45276 3556 45332
rect 46060 46562 46116 46564
rect 46060 46510 46062 46562
rect 46062 46510 46114 46562
rect 46114 46510 46116 46562
rect 46060 46508 46116 46510
rect 46844 46508 46900 46564
rect 47628 46508 47684 46564
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 46172 45778 46228 45780
rect 46172 45726 46174 45778
rect 46174 45726 46226 45778
rect 46226 45726 46228 45778
rect 46172 45724 46228 45726
rect 46844 45778 46900 45780
rect 46844 45726 46846 45778
rect 46846 45726 46898 45778
rect 46898 45726 46900 45778
rect 46844 45724 46900 45726
rect 45836 45666 45892 45668
rect 45836 45614 45838 45666
rect 45838 45614 45890 45666
rect 45890 45614 45892 45666
rect 45836 45612 45892 45614
rect 46508 45612 46564 45668
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 44380 45330 44436 45332
rect 44380 45278 44382 45330
rect 44382 45278 44434 45330
rect 44434 45278 44436 45330
rect 44380 45276 44436 45278
rect 3612 45164 3668 45220
rect 45276 45218 45332 45220
rect 45276 45166 45278 45218
rect 45278 45166 45330 45218
rect 45330 45166 45332 45218
rect 45276 45164 45332 45166
rect 2156 44940 2212 44996
rect 43932 45106 43988 45108
rect 43932 45054 43934 45106
rect 43934 45054 43986 45106
rect 43986 45054 43988 45106
rect 43932 45052 43988 45054
rect 44604 45106 44660 45108
rect 44604 45054 44606 45106
rect 44606 45054 44658 45106
rect 44658 45054 44660 45106
rect 44604 45052 44660 45054
rect 45612 45106 45668 45108
rect 45612 45054 45614 45106
rect 45614 45054 45666 45106
rect 45666 45054 45668 45106
rect 45612 45052 45668 45054
rect 46284 45106 46340 45108
rect 46284 45054 46286 45106
rect 46286 45054 46338 45106
rect 46338 45054 46340 45106
rect 46284 45052 46340 45054
rect 3052 44940 3108 44996
rect 3612 44994 3668 44996
rect 3612 44942 3614 44994
rect 3614 44942 3666 44994
rect 3666 44942 3668 44994
rect 3612 44940 3668 44942
rect 43708 44940 43764 44996
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 2044 44268 2100 44324
rect 46396 44940 46452 44996
rect 44044 44210 44100 44212
rect 44044 44158 44046 44210
rect 44046 44158 44098 44210
rect 44098 44158 44100 44210
rect 44044 44156 44100 44158
rect 44604 44210 44660 44212
rect 44604 44158 44606 44210
rect 44606 44158 44658 44210
rect 44658 44158 44660 44210
rect 44604 44156 44660 44158
rect 45276 44156 45332 44212
rect 3052 44044 3108 44100
rect 3500 44098 3556 44100
rect 3500 44046 3502 44098
rect 3502 44046 3554 44098
rect 3554 44046 3556 44098
rect 3500 44044 3556 44046
rect 42924 44044 42980 44100
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 44380 43762 44436 43764
rect 44380 43710 44382 43762
rect 44382 43710 44434 43762
rect 44434 43710 44436 43762
rect 44380 43708 44436 43710
rect 2156 43596 2212 43652
rect 3052 43372 3108 43428
rect 3612 43426 3668 43428
rect 3612 43374 3614 43426
rect 3614 43374 3666 43426
rect 3666 43374 3668 43426
rect 3612 43372 3668 43374
rect 42252 43372 42308 43428
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 2044 42924 2100 42980
rect 41916 42754 41972 42756
rect 41916 42702 41918 42754
rect 41918 42702 41970 42754
rect 41970 42702 41972 42754
rect 41916 42700 41972 42702
rect 42476 43426 42532 43428
rect 42476 43374 42478 43426
rect 42478 43374 42530 43426
rect 42530 43374 42532 43426
rect 42476 43372 42532 43374
rect 43260 43372 43316 43428
rect 44268 43372 44324 43428
rect 42588 42754 42644 42756
rect 42588 42702 42590 42754
rect 42590 42702 42642 42754
rect 42642 42702 42644 42754
rect 42588 42700 42644 42702
rect 43372 42754 43428 42756
rect 43372 42702 43374 42754
rect 43374 42702 43426 42754
rect 43426 42702 43428 42754
rect 43372 42700 43428 42702
rect 44044 42588 44100 42644
rect 3052 42476 3108 42532
rect 3500 42530 3556 42532
rect 3500 42478 3502 42530
rect 3502 42478 3554 42530
rect 3554 42478 3556 42530
rect 3500 42476 3556 42478
rect 41692 42476 41748 42532
rect 2156 42252 2212 42308
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 43708 42530 43764 42532
rect 43708 42478 43710 42530
rect 43710 42478 43762 42530
rect 43762 42478 43764 42530
rect 43708 42476 43764 42478
rect 3052 41804 3108 41860
rect 3612 41858 3668 41860
rect 3612 41806 3614 41858
rect 3614 41806 3666 41858
rect 3666 41806 3668 41858
rect 3612 41804 3668 41806
rect 41020 41804 41076 41860
rect 2044 41580 2100 41636
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 2156 40908 2212 40964
rect 42028 41804 42084 41860
rect 42924 41804 42980 41860
rect 3052 40908 3108 40964
rect 3500 40962 3556 40964
rect 3500 40910 3502 40962
rect 3502 40910 3554 40962
rect 3554 40910 3556 40962
rect 3500 40908 3556 40910
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 3052 40402 3108 40404
rect 3052 40350 3054 40402
rect 3054 40350 3106 40402
rect 3106 40350 3108 40402
rect 3052 40348 3108 40350
rect 3612 40402 3668 40404
rect 3612 40350 3614 40402
rect 3614 40350 3666 40402
rect 3666 40350 3668 40402
rect 3612 40348 3668 40350
rect 39340 40348 39396 40404
rect 40236 40908 40292 40964
rect 40572 40962 40628 40964
rect 40572 40910 40574 40962
rect 40574 40910 40626 40962
rect 40626 40910 40628 40962
rect 40572 40908 40628 40910
rect 41356 40908 41412 40964
rect 42364 41074 42420 41076
rect 42364 41022 42366 41074
rect 42366 41022 42418 41074
rect 42418 41022 42420 41074
rect 42364 41020 42420 41022
rect 42140 40908 42196 40964
rect 41916 40514 41972 40516
rect 41916 40462 41918 40514
rect 41918 40462 41970 40514
rect 41970 40462 41972 40514
rect 41916 40460 41972 40462
rect 2044 40290 2100 40292
rect 2044 40238 2046 40290
rect 2046 40238 2098 40290
rect 2098 40238 2100 40290
rect 2044 40236 2100 40238
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 2156 39618 2212 39620
rect 2156 39566 2158 39618
rect 2158 39566 2210 39618
rect 2210 39566 2212 39618
rect 2156 39564 2212 39566
rect 3052 39452 3108 39508
rect 3612 39506 3668 39508
rect 3612 39454 3614 39506
rect 3614 39454 3666 39506
rect 3666 39454 3668 39506
rect 3612 39452 3668 39454
rect 38780 39506 38836 39508
rect 38780 39454 38782 39506
rect 38782 39454 38834 39506
rect 38834 39454 38836 39506
rect 38780 39452 38836 39454
rect 38332 39394 38388 39396
rect 38332 39342 38334 39394
rect 38334 39342 38386 39394
rect 38386 39342 38388 39394
rect 38332 39340 38388 39342
rect 38892 39340 38948 39396
rect 39116 39506 39172 39508
rect 39116 39454 39118 39506
rect 39118 39454 39170 39506
rect 39170 39454 39172 39506
rect 39116 39452 39172 39454
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 2156 38946 2212 38948
rect 2156 38894 2158 38946
rect 2158 38894 2210 38946
rect 2210 38894 2212 38946
rect 2156 38892 2212 38894
rect 3052 38834 3108 38836
rect 3052 38782 3054 38834
rect 3054 38782 3106 38834
rect 3106 38782 3108 38834
rect 3052 38780 3108 38782
rect 3612 38834 3668 38836
rect 3612 38782 3614 38834
rect 3614 38782 3666 38834
rect 3666 38782 3668 38834
rect 3612 38780 3668 38782
rect 38332 38780 38388 38836
rect 38668 38834 38724 38836
rect 38668 38782 38670 38834
rect 38670 38782 38722 38834
rect 38722 38782 38724 38834
rect 38668 38780 38724 38782
rect 37884 38722 37940 38724
rect 37884 38670 37886 38722
rect 37886 38670 37938 38722
rect 37938 38670 37940 38722
rect 37884 38668 37940 38670
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 2044 38220 2100 38276
rect 37996 37938 38052 37940
rect 37996 37886 37998 37938
rect 37998 37886 38050 37938
rect 38050 37886 38052 37938
rect 37996 37884 38052 37886
rect 38668 37938 38724 37940
rect 38668 37886 38670 37938
rect 38670 37886 38722 37938
rect 38722 37886 38724 37938
rect 38668 37884 38724 37886
rect 3052 37772 3108 37828
rect 3612 37826 3668 37828
rect 3612 37774 3614 37826
rect 3614 37774 3666 37826
rect 3666 37774 3668 37826
rect 3612 37772 3668 37774
rect 37660 37826 37716 37828
rect 37660 37774 37662 37826
rect 37662 37774 37714 37826
rect 37714 37774 37716 37826
rect 37660 37772 37716 37774
rect 19836 37658 19892 37660
rect 2156 37548 2212 37604
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 3052 36988 3108 37044
rect 36540 37154 36596 37156
rect 36540 37102 36542 37154
rect 36542 37102 36594 37154
rect 36594 37102 36596 37154
rect 36540 37100 36596 37102
rect 3612 36988 3668 37044
rect 38332 37378 38388 37380
rect 38332 37326 38334 37378
rect 38334 37326 38386 37378
rect 38386 37326 38388 37378
rect 38332 37324 38388 37326
rect 36988 36988 37044 37044
rect 37212 37100 37268 37156
rect 2044 36876 2100 36932
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 2156 36204 2212 36260
rect 35868 36370 35924 36372
rect 35868 36318 35870 36370
rect 35870 36318 35922 36370
rect 35922 36318 35924 36370
rect 35868 36316 35924 36318
rect 36652 36370 36708 36372
rect 36652 36318 36654 36370
rect 36654 36318 36706 36370
rect 36706 36318 36708 36370
rect 36652 36316 36708 36318
rect 3052 36204 3108 36260
rect 3612 36258 3668 36260
rect 3612 36206 3614 36258
rect 3614 36206 3666 36258
rect 3666 36206 3668 36258
rect 3612 36204 3668 36206
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 3052 35756 3108 35812
rect 3612 35756 3668 35812
rect 2044 35532 2100 35588
rect 4844 35532 4900 35588
rect 5404 35586 5460 35588
rect 5404 35534 5406 35586
rect 5406 35534 5458 35586
rect 5458 35534 5460 35586
rect 5404 35532 5460 35534
rect 34188 35532 34244 35588
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 3836 34860 3892 34916
rect 33740 34914 33796 34916
rect 33740 34862 33742 34914
rect 33742 34862 33794 34914
rect 33794 34862 33796 34914
rect 33740 34860 33796 34862
rect 34524 34914 34580 34916
rect 34524 34862 34526 34914
rect 34526 34862 34578 34914
rect 34578 34862 34580 34914
rect 34524 34860 34580 34862
rect 3052 34636 3108 34692
rect 4060 34690 4116 34692
rect 4060 34638 4062 34690
rect 4062 34638 4114 34690
rect 4114 34638 4116 34690
rect 4060 34636 4116 34638
rect 34972 35698 35028 35700
rect 34972 35646 34974 35698
rect 34974 35646 35026 35698
rect 35026 35646 35028 35698
rect 34972 35644 35028 35646
rect 36316 36258 36372 36260
rect 36316 36206 36318 36258
rect 36318 36206 36370 36258
rect 36370 36206 36372 36258
rect 36316 36204 36372 36206
rect 35532 35810 35588 35812
rect 35532 35758 35534 35810
rect 35534 35758 35586 35810
rect 35586 35758 35588 35810
rect 35532 35756 35588 35758
rect 35868 35810 35924 35812
rect 35868 35758 35870 35810
rect 35870 35758 35922 35810
rect 35922 35758 35924 35810
rect 35868 35756 35924 35758
rect 36764 35756 36820 35812
rect 35308 35644 35364 35700
rect 36092 35644 36148 35700
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 34914 35252 34916
rect 35196 34862 35198 34914
rect 35198 34862 35250 34914
rect 35250 34862 35252 34914
rect 35196 34860 35252 34862
rect 34636 34636 34692 34692
rect 35420 34690 35476 34692
rect 35420 34638 35422 34690
rect 35422 34638 35474 34690
rect 35474 34638 35476 34690
rect 35420 34636 35476 34638
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 2156 34242 2212 34244
rect 2156 34190 2158 34242
rect 2158 34190 2210 34242
rect 2210 34190 2212 34242
rect 2156 34188 2212 34190
rect 32956 34130 33012 34132
rect 32956 34078 32958 34130
rect 32958 34078 33010 34130
rect 33010 34078 33012 34130
rect 32956 34076 33012 34078
rect 3052 33852 3108 33908
rect 3612 33852 3668 33908
rect 35084 34242 35140 34244
rect 35084 34190 35086 34242
rect 35086 34190 35138 34242
rect 35138 34190 35140 34242
rect 35084 34188 35140 34190
rect 33964 34130 34020 34132
rect 33964 34078 33966 34130
rect 33966 34078 34018 34130
rect 34018 34078 34020 34130
rect 33964 34076 34020 34078
rect 34860 34130 34916 34132
rect 34860 34078 34862 34130
rect 34862 34078 34914 34130
rect 34914 34078 34916 34130
rect 34860 34076 34916 34078
rect 33628 33852 33684 33908
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 2044 33516 2100 33572
rect 32508 33346 32564 33348
rect 32508 33294 32510 33346
rect 32510 33294 32562 33346
rect 32562 33294 32564 33346
rect 32508 33292 32564 33294
rect 33180 33346 33236 33348
rect 33180 33294 33182 33346
rect 33182 33294 33234 33346
rect 33234 33294 33236 33346
rect 33180 33292 33236 33294
rect 3052 33068 3108 33124
rect 3612 33122 3668 33124
rect 3612 33070 3614 33122
rect 3614 33070 3666 33122
rect 3666 33070 3668 33122
rect 3612 33068 3668 33070
rect 32956 33122 33012 33124
rect 32956 33070 32958 33122
rect 32958 33070 33010 33122
rect 33010 33070 33012 33122
rect 32956 33068 33012 33070
rect 19836 32954 19892 32956
rect 2156 32844 2212 32900
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 3052 32284 3108 32340
rect 31724 32450 31780 32452
rect 31724 32398 31726 32450
rect 31726 32398 31778 32450
rect 31778 32398 31780 32450
rect 31724 32396 31780 32398
rect 3612 32284 3668 32340
rect 32172 32284 32228 32340
rect 32508 32562 32564 32564
rect 32508 32510 32510 32562
rect 32510 32510 32562 32562
rect 32562 32510 32564 32562
rect 32508 32508 32564 32510
rect 2044 32172 2100 32228
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 34076 33346 34132 33348
rect 34076 33294 34078 33346
rect 34078 33294 34130 33346
rect 34130 33294 34132 33346
rect 34076 33292 34132 33294
rect 34412 33122 34468 33124
rect 34412 33070 34414 33122
rect 34414 33070 34466 33122
rect 34466 33070 34468 33122
rect 34412 33068 34468 33070
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 33964 32674 34020 32676
rect 33964 32622 33966 32674
rect 33966 32622 34018 32674
rect 34018 32622 34020 32674
rect 33964 32620 34020 32622
rect 33404 32508 33460 32564
rect 2156 31500 2212 31556
rect 31164 31666 31220 31668
rect 31164 31614 31166 31666
rect 31166 31614 31218 31666
rect 31218 31614 31220 31666
rect 31164 31612 31220 31614
rect 31948 31666 32004 31668
rect 31948 31614 31950 31666
rect 31950 31614 32002 31666
rect 32002 31614 32004 31666
rect 31948 31612 32004 31614
rect 3052 31500 3108 31556
rect 3612 31554 3668 31556
rect 3612 31502 3614 31554
rect 3614 31502 3666 31554
rect 3666 31502 3668 31554
rect 3612 31500 3668 31502
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 3052 31052 3108 31108
rect 3612 31052 3668 31108
rect 2156 30828 2212 30884
rect 4844 30828 4900 30884
rect 5404 30882 5460 30884
rect 5404 30830 5406 30882
rect 5406 30830 5458 30882
rect 5458 30830 5460 30882
rect 5404 30828 5460 30830
rect 29596 30828 29652 30884
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 3836 30156 3892 30212
rect 3052 29932 3108 29988
rect 4060 29986 4116 29988
rect 4060 29934 4062 29986
rect 4062 29934 4114 29986
rect 4114 29934 4116 29986
rect 4060 29932 4116 29934
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 2156 29538 2212 29540
rect 2156 29486 2158 29538
rect 2158 29486 2210 29538
rect 2210 29486 2212 29538
rect 2156 29484 2212 29486
rect 3052 29148 3108 29204
rect 28252 29314 28308 29316
rect 28252 29262 28254 29314
rect 28254 29262 28306 29314
rect 28306 29262 28308 29314
rect 28252 29260 28308 29262
rect 3612 29148 3668 29204
rect 28700 29148 28756 29204
rect 30044 29932 30100 29988
rect 31612 31554 31668 31556
rect 31612 31502 31614 31554
rect 31614 31502 31666 31554
rect 31666 31502 31668 31554
rect 31612 31500 31668 31502
rect 30940 31106 30996 31108
rect 30940 31054 30942 31106
rect 30942 31054 30994 31106
rect 30994 31054 30996 31106
rect 30940 31052 30996 31054
rect 31276 30994 31332 30996
rect 31276 30942 31278 30994
rect 31278 30942 31330 30994
rect 31330 30942 31332 30994
rect 31276 30940 31332 30942
rect 29932 29426 29988 29428
rect 29932 29374 29934 29426
rect 29934 29374 29986 29426
rect 29986 29374 29988 29426
rect 29932 29372 29988 29374
rect 29036 29260 29092 29316
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 2044 28812 2100 28868
rect 3052 28642 3108 28644
rect 3052 28590 3054 28642
rect 3054 28590 3106 28642
rect 3106 28590 3108 28642
rect 3052 28588 3108 28590
rect 3612 28642 3668 28644
rect 3612 28590 3614 28642
rect 3614 28590 3666 28642
rect 3666 28590 3668 28642
rect 3612 28588 3668 28590
rect 27804 28476 27860 28532
rect 28252 28588 28308 28644
rect 32060 30994 32116 30996
rect 32060 30942 32062 30994
rect 32062 30942 32114 30994
rect 32114 30942 32116 30994
rect 32060 30940 32116 30942
rect 30716 29986 30772 29988
rect 30716 29934 30718 29986
rect 30718 29934 30770 29986
rect 30770 29934 30772 29986
rect 30716 29932 30772 29934
rect 30828 29538 30884 29540
rect 30828 29486 30830 29538
rect 30830 29486 30882 29538
rect 30882 29486 30884 29538
rect 30828 29484 30884 29486
rect 30380 29372 30436 29428
rect 29036 28588 29092 28644
rect 29708 28588 29764 28644
rect 28588 28530 28644 28532
rect 28588 28478 28590 28530
rect 28590 28478 28642 28530
rect 28642 28478 28644 28530
rect 28588 28476 28644 28478
rect 29372 28476 29428 28532
rect 19836 28250 19892 28252
rect 2156 28140 2212 28196
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 27132 27858 27188 27860
rect 27132 27806 27134 27858
rect 27134 27806 27186 27858
rect 27186 27806 27188 27858
rect 27132 27804 27188 27806
rect 3052 27692 3108 27748
rect 3612 27746 3668 27748
rect 3612 27694 3614 27746
rect 3614 27694 3666 27746
rect 3666 27694 3668 27746
rect 3612 27692 3668 27694
rect 28924 27970 28980 27972
rect 28924 27918 28926 27970
rect 28926 27918 28978 27970
rect 28978 27918 28980 27970
rect 28924 27916 28980 27918
rect 27916 27858 27972 27860
rect 27916 27806 27918 27858
rect 27918 27806 27970 27858
rect 27970 27806 27972 27858
rect 27916 27804 27972 27806
rect 28476 27804 28532 27860
rect 27580 27692 27636 27748
rect 2044 27468 2100 27524
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 3052 27074 3108 27076
rect 3052 27022 3054 27074
rect 3054 27022 3106 27074
rect 3106 27022 3108 27074
rect 3052 27020 3108 27022
rect 3612 27074 3668 27076
rect 3612 27022 3614 27074
rect 3614 27022 3666 27074
rect 3666 27022 3668 27074
rect 3612 27020 3668 27022
rect 26908 27020 26964 27076
rect 26460 26962 26516 26964
rect 26460 26910 26462 26962
rect 26462 26910 26514 26962
rect 26514 26910 26516 26962
rect 26460 26908 26516 26910
rect 2156 26796 2212 26852
rect 27244 26962 27300 26964
rect 27244 26910 27246 26962
rect 27246 26910 27298 26962
rect 27298 26910 27300 26962
rect 27244 26908 27300 26910
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 2044 26124 2100 26180
rect 4844 26124 4900 26180
rect 5404 26178 5460 26180
rect 5404 26126 5406 26178
rect 5406 26126 5458 26178
rect 5458 26126 5460 26178
rect 5404 26124 5460 26126
rect 24332 26124 24388 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 3836 25452 3892 25508
rect 3052 25340 3108 25396
rect 4060 25394 4116 25396
rect 4060 25342 4062 25394
rect 4062 25342 4114 25394
rect 4114 25342 4116 25394
rect 4060 25340 4116 25342
rect 25788 26178 25844 26180
rect 25788 26126 25790 26178
rect 25790 26126 25842 26178
rect 25842 26126 25844 26178
rect 25788 26124 25844 26126
rect 25564 25506 25620 25508
rect 25564 25454 25566 25506
rect 25566 25454 25618 25506
rect 25618 25454 25620 25506
rect 25564 25452 25620 25454
rect 2940 25228 2996 25284
rect 3612 25282 3668 25284
rect 3612 25230 3614 25282
rect 3614 25230 3666 25282
rect 3666 25230 3668 25282
rect 3612 25228 3668 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 2156 24834 2212 24836
rect 2156 24782 2158 24834
rect 2158 24782 2210 24834
rect 2210 24782 2212 24834
rect 2156 24780 2212 24782
rect 3052 24556 3108 24612
rect 3612 24610 3668 24612
rect 3612 24558 3614 24610
rect 3614 24558 3666 24610
rect 3666 24558 3668 24610
rect 3612 24556 3668 24558
rect 24108 24556 24164 24612
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 2044 24108 2100 24164
rect 3052 23660 3108 23716
rect 3612 23714 3668 23716
rect 3612 23662 3614 23714
rect 3614 23662 3666 23714
rect 3666 23662 3668 23714
rect 3612 23660 3668 23662
rect 19836 23546 19892 23548
rect 2156 23436 2212 23492
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 3052 22988 3108 23044
rect 3612 23042 3668 23044
rect 3612 22990 3614 23042
rect 3614 22990 3666 23042
rect 3666 22990 3668 23042
rect 3612 22988 3668 22990
rect 22764 23154 22820 23156
rect 22764 23102 22766 23154
rect 22766 23102 22818 23154
rect 22818 23102 22820 23154
rect 22764 23100 22820 23102
rect 23660 23714 23716 23716
rect 23660 23662 23662 23714
rect 23662 23662 23714 23714
rect 23714 23662 23716 23714
rect 23660 23660 23716 23662
rect 25228 25394 25284 25396
rect 25228 25342 25230 25394
rect 25230 25342 25282 25394
rect 25282 25342 25284 25394
rect 25228 25340 25284 25342
rect 26460 26124 26516 26180
rect 26236 25228 26292 25284
rect 26348 25452 26404 25508
rect 26124 24834 26180 24836
rect 26124 24782 26126 24834
rect 26126 24782 26178 24834
rect 26178 24782 26180 24834
rect 26124 24780 26180 24782
rect 24892 24610 24948 24612
rect 24892 24558 24894 24610
rect 24894 24558 24946 24610
rect 24946 24558 24948 24610
rect 24892 24556 24948 24558
rect 25900 24556 25956 24612
rect 24668 23714 24724 23716
rect 24668 23662 24670 23714
rect 24670 23662 24722 23714
rect 24722 23662 24724 23714
rect 24668 23660 24724 23662
rect 25564 23660 25620 23716
rect 23996 23548 24052 23604
rect 23884 23266 23940 23268
rect 23884 23214 23886 23266
rect 23886 23214 23938 23266
rect 23938 23214 23940 23266
rect 23884 23212 23940 23214
rect 23100 23100 23156 23156
rect 23660 23154 23716 23156
rect 23660 23102 23662 23154
rect 23662 23102 23714 23154
rect 23714 23102 23716 23154
rect 23660 23100 23716 23102
rect 22428 22988 22484 23044
rect 2044 22764 2100 22820
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 3052 22204 3108 22260
rect 3612 22258 3668 22260
rect 3612 22206 3614 22258
rect 3614 22206 3666 22258
rect 3666 22206 3668 22258
rect 3612 22204 3668 22206
rect 22092 22258 22148 22260
rect 22092 22206 22094 22258
rect 22094 22206 22146 22258
rect 22146 22206 22148 22258
rect 22092 22204 22148 22206
rect 22428 22258 22484 22260
rect 22428 22206 22430 22258
rect 22430 22206 22482 22258
rect 22482 22206 22484 22258
rect 22428 22204 22484 22206
rect 2156 22092 2212 22148
rect 21644 22146 21700 22148
rect 21644 22094 21646 22146
rect 21646 22094 21698 22146
rect 21698 22094 21700 22146
rect 21644 22092 21700 22094
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 2044 21420 2100 21476
rect 4844 21420 4900 21476
rect 5404 21474 5460 21476
rect 5404 21422 5406 21474
rect 5406 21422 5458 21474
rect 5458 21422 5460 21474
rect 5404 21420 5460 21422
rect 19628 21420 19684 21476
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 3836 20748 3892 20804
rect 3052 20636 3108 20692
rect 4060 20690 4116 20692
rect 4060 20638 4062 20690
rect 4062 20638 4114 20690
rect 4114 20638 4116 20690
rect 4060 20636 4116 20638
rect 2940 20524 2996 20580
rect 3612 20578 3668 20580
rect 3612 20526 3614 20578
rect 3614 20526 3666 20578
rect 3666 20526 3668 20578
rect 3612 20524 3668 20526
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 2156 20130 2212 20132
rect 2156 20078 2158 20130
rect 2158 20078 2210 20130
rect 2210 20078 2212 20130
rect 2156 20076 2212 20078
rect 19516 20018 19572 20020
rect 19516 19966 19518 20018
rect 19518 19966 19570 20018
rect 19570 19966 19572 20018
rect 19516 19964 19572 19966
rect 20300 20018 20356 20020
rect 20300 19966 20302 20018
rect 20302 19966 20354 20018
rect 20354 19966 20356 20018
rect 20300 19964 20356 19966
rect 3052 19852 3108 19908
rect 3612 19906 3668 19908
rect 3612 19854 3614 19906
rect 3614 19854 3666 19906
rect 3666 19854 3668 19906
rect 3612 19852 3668 19854
rect 19404 19852 19460 19908
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 2044 19404 2100 19460
rect 3052 18844 3108 18900
rect 3612 18844 3668 18900
rect 2156 18732 2212 18788
rect 18620 18844 18676 18900
rect 18172 18620 18228 18676
rect 19852 19122 19908 19124
rect 19852 19070 19854 19122
rect 19854 19070 19906 19122
rect 19906 19070 19908 19122
rect 19852 19068 19908 19070
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 18956 18620 19012 18676
rect 3052 18284 3108 18340
rect 3612 18338 3668 18340
rect 3612 18286 3614 18338
rect 3614 18286 3666 18338
rect 3666 18286 3668 18338
rect 3612 18284 3668 18286
rect 2044 18060 2100 18116
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 2156 17388 2212 17444
rect 20076 18508 20132 18564
rect 18620 18284 18676 18340
rect 18956 17836 19012 17892
rect 3052 17388 3108 17444
rect 3612 17442 3668 17444
rect 3612 17390 3614 17442
rect 3614 17390 3666 17442
rect 3666 17390 3668 17442
rect 3612 17388 3668 17390
rect 3052 16940 3108 16996
rect 3612 16940 3668 16996
rect 2044 16716 2100 16772
rect 4844 16882 4900 16884
rect 4844 16830 4846 16882
rect 4846 16830 4898 16882
rect 4898 16830 4900 16882
rect 4844 16828 4900 16830
rect 5404 16882 5460 16884
rect 5404 16830 5406 16882
rect 5406 16830 5458 16882
rect 5458 16830 5460 16882
rect 5404 16828 5460 16830
rect 15596 16828 15652 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 3836 16044 3892 16100
rect 3052 15820 3108 15876
rect 4060 15874 4116 15876
rect 4060 15822 4062 15874
rect 4062 15822 4114 15874
rect 4114 15822 4116 15874
rect 4060 15820 4116 15822
rect 15820 15820 15876 15876
rect 16604 16994 16660 16996
rect 16604 16942 16606 16994
rect 16606 16942 16658 16994
rect 16658 16942 16660 16994
rect 16604 16940 16660 16942
rect 2156 15426 2212 15428
rect 2156 15374 2158 15426
rect 2158 15374 2210 15426
rect 2210 15374 2212 15426
rect 2156 15372 2212 15374
rect 3052 15148 3108 15204
rect 3612 15202 3668 15204
rect 3612 15150 3614 15202
rect 3614 15150 3666 15202
rect 3666 15150 3668 15202
rect 3612 15148 3668 15150
rect 14700 15148 14756 15204
rect 15484 15260 15540 15316
rect 17724 17442 17780 17444
rect 17724 17390 17726 17442
rect 17726 17390 17778 17442
rect 17778 17390 17780 17442
rect 17724 17388 17780 17390
rect 17052 16828 17108 16884
rect 15932 15148 15988 15204
rect 16044 15820 16100 15876
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 2044 14700 2100 14756
rect 14364 14418 14420 14420
rect 14364 14366 14366 14418
rect 14366 14366 14418 14418
rect 14418 14366 14420 14418
rect 14364 14364 14420 14366
rect 14812 14418 14868 14420
rect 14812 14366 14814 14418
rect 14814 14366 14866 14418
rect 14866 14366 14868 14418
rect 14812 14364 14868 14366
rect 3052 14252 3108 14308
rect 3612 14306 3668 14308
rect 3612 14254 3614 14306
rect 3614 14254 3666 14306
rect 3666 14254 3668 14306
rect 3612 14252 3668 14254
rect 14028 14306 14084 14308
rect 14028 14254 14030 14306
rect 14030 14254 14082 14306
rect 14082 14254 14084 14306
rect 14028 14252 14084 14254
rect 2156 14028 2212 14084
rect 12012 13746 12068 13748
rect 12012 13694 12014 13746
rect 12014 13694 12066 13746
rect 12066 13694 12068 13746
rect 12012 13692 12068 13694
rect 3052 13580 3108 13636
rect 3612 13634 3668 13636
rect 3612 13582 3614 13634
rect 3614 13582 3666 13634
rect 3666 13582 3668 13634
rect 3612 13580 3668 13582
rect 2044 13356 2100 13412
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 2156 12684 2212 12740
rect 3052 12684 3108 12740
rect 3612 12738 3668 12740
rect 3612 12686 3614 12738
rect 3614 12686 3666 12738
rect 3666 12686 3668 12738
rect 3612 12684 3668 12686
rect 3052 12236 3108 12292
rect 3612 12236 3668 12292
rect 2044 12012 2100 12068
rect 3052 11452 3108 11508
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4060 11506 4116 11508
rect 4060 11454 4062 11506
rect 4062 11454 4114 11506
rect 4114 11454 4116 11506
rect 4060 11452 4116 11454
rect 3836 11340 3892 11396
rect 12796 13746 12852 13748
rect 12796 13694 12798 13746
rect 12798 13694 12850 13746
rect 12850 13694 12852 13746
rect 12796 13692 12852 13694
rect 13356 13580 13412 13636
rect 13692 13468 13748 13524
rect 12460 12684 12516 12740
rect 12236 12290 12292 12292
rect 12236 12238 12238 12290
rect 12238 12238 12290 12290
rect 12290 12238 12292 12290
rect 12236 12236 12292 12238
rect 12684 12124 12740 12180
rect 11340 11452 11396 11508
rect 4844 11228 4900 11284
rect 10780 11282 10836 11284
rect 10780 11230 10782 11282
rect 10782 11230 10834 11282
rect 10834 11230 10836 11282
rect 10780 11228 10836 11230
rect 2156 10722 2212 10724
rect 2156 10670 2158 10722
rect 2158 10670 2210 10722
rect 2210 10670 2212 10722
rect 2156 10668 2212 10670
rect 3052 10668 3108 10724
rect 10108 10722 10164 10724
rect 10108 10670 10110 10722
rect 10110 10670 10162 10722
rect 10162 10670 10164 10722
rect 10108 10668 10164 10670
rect 11452 10722 11508 10724
rect 11452 10670 11454 10722
rect 11454 10670 11506 10722
rect 11506 10670 11508 10722
rect 11452 10668 11508 10670
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 2044 9996 2100 10052
rect 3052 9660 3108 9716
rect 9436 9714 9492 9716
rect 9436 9662 9438 9714
rect 9438 9662 9490 9714
rect 9490 9662 9492 9714
rect 9436 9660 9492 9662
rect 9660 9660 9716 9716
rect 2156 9324 2212 9380
rect 3052 9100 3108 9156
rect 8652 9154 8708 9156
rect 8652 9102 8654 9154
rect 8654 9102 8706 9154
rect 8706 9102 8708 9154
rect 8652 9100 8708 9102
rect 8988 9042 9044 9044
rect 8988 8990 8990 9042
rect 8990 8990 9042 9042
rect 9042 8990 9044 9042
rect 8988 8988 9044 8990
rect 2044 8652 2100 8708
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 3052 8092 3108 8148
rect 7980 8146 8036 8148
rect 7980 8094 7982 8146
rect 7982 8094 8034 8146
rect 8034 8094 8036 8146
rect 7980 8092 8036 8094
rect 8316 8146 8372 8148
rect 8316 8094 8318 8146
rect 8318 8094 8370 8146
rect 8370 8094 8372 8146
rect 8316 8092 8372 8094
rect 2156 7980 2212 8036
rect 3052 7532 3108 7588
rect 2156 7308 2212 7364
rect 3052 6748 3108 6804
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 3836 6636 3892 6692
rect 7420 7586 7476 7588
rect 7420 7534 7422 7586
rect 7422 7534 7474 7586
rect 7474 7534 7476 7586
rect 7420 7532 7476 7534
rect 8764 7586 8820 7588
rect 8764 7534 8766 7586
rect 8766 7534 8818 7586
rect 8818 7534 8820 7586
rect 8764 7532 8820 7534
rect 6524 6748 6580 6804
rect 6972 6636 7028 6692
rect 4844 6524 4900 6580
rect 5964 6578 6020 6580
rect 5964 6526 5966 6578
rect 5966 6526 6018 6578
rect 6018 6526 6020 6578
rect 5964 6524 6020 6526
rect 6300 6578 6356 6580
rect 6300 6526 6302 6578
rect 6302 6526 6354 6578
rect 6354 6526 6356 6578
rect 6300 6524 6356 6526
rect 6860 6578 6916 6580
rect 6860 6526 6862 6578
rect 6862 6526 6914 6578
rect 6914 6526 6916 6578
rect 6860 6524 6916 6526
rect 2156 6018 2212 6020
rect 2156 5966 2158 6018
rect 2158 5966 2210 6018
rect 2210 5966 2212 6018
rect 2156 5964 2212 5966
rect 3052 5964 3108 6020
rect 5292 6018 5348 6020
rect 5292 5966 5294 6018
rect 5294 5966 5346 6018
rect 5346 5966 5348 6018
rect 5292 5964 5348 5966
rect 6748 6018 6804 6020
rect 6748 5966 6750 6018
rect 6750 5966 6802 6018
rect 6802 5966 6804 6018
rect 6748 5964 6804 5966
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 2044 5292 2100 5348
rect 3052 4956 3108 5012
rect 4620 5010 4676 5012
rect 4620 4958 4622 5010
rect 4622 4958 4674 5010
rect 4674 4958 4676 5010
rect 4620 4956 4676 4958
rect 4956 5010 5012 5012
rect 4956 4958 4958 5010
rect 4958 4958 5010 5010
rect 5010 4958 5012 5010
rect 4956 4956 5012 4958
rect 5740 5010 5796 5012
rect 5740 4958 5742 5010
rect 5742 4958 5794 5010
rect 5794 4958 5796 5010
rect 5740 4956 5796 4958
rect 6076 4898 6132 4900
rect 6076 4846 6078 4898
rect 6078 4846 6130 4898
rect 6130 4846 6132 4898
rect 6076 4844 6132 4846
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 5068 3442 5124 3444
rect 5068 3390 5070 3442
rect 5070 3390 5122 3442
rect 5122 3390 5124 3442
rect 5068 3388 5124 3390
rect 5964 3388 6020 3444
rect 7644 7474 7700 7476
rect 7644 7422 7646 7474
rect 7646 7422 7698 7474
rect 7698 7422 7700 7474
rect 7644 7420 7700 7422
rect 7196 6466 7252 6468
rect 7196 6414 7198 6466
rect 7198 6414 7250 6466
rect 7250 6414 7252 6466
rect 7196 6412 7252 6414
rect 8428 7474 8484 7476
rect 8428 7422 8430 7474
rect 8430 7422 8482 7474
rect 8482 7422 8484 7474
rect 8428 7420 8484 7422
rect 7756 6690 7812 6692
rect 7756 6638 7758 6690
rect 7758 6638 7810 6690
rect 7810 6638 7812 6690
rect 7756 6636 7812 6638
rect 8092 6578 8148 6580
rect 8092 6526 8094 6578
rect 8094 6526 8146 6578
rect 8146 6526 8148 6578
rect 8092 6524 8148 6526
rect 6412 4284 6468 4340
rect 7084 4338 7140 4340
rect 7084 4286 7086 4338
rect 7086 4286 7138 4338
rect 7138 4286 7140 4338
rect 7084 4284 7140 4286
rect 8540 3442 8596 3444
rect 8540 3390 8542 3442
rect 8542 3390 8594 3442
rect 8594 3390 8596 3442
rect 8540 3388 8596 3390
rect 9100 8146 9156 8148
rect 9100 8094 9102 8146
rect 9102 8094 9154 8146
rect 9154 8094 9156 8146
rect 9100 8092 9156 8094
rect 9436 8034 9492 8036
rect 9436 7982 9438 8034
rect 9438 7982 9490 8034
rect 9490 7982 9492 8034
rect 9436 7980 9492 7982
rect 8988 4284 9044 4340
rect 9324 3388 9380 3444
rect 10556 9714 10612 9716
rect 10556 9662 10558 9714
rect 10558 9662 10610 9714
rect 10610 9662 10612 9714
rect 10556 9660 10612 9662
rect 10892 9602 10948 9604
rect 10892 9550 10894 9602
rect 10894 9550 10946 9602
rect 10946 9550 10948 9602
rect 10892 9548 10948 9550
rect 10220 9154 10276 9156
rect 10220 9102 10222 9154
rect 10222 9102 10274 9154
rect 10274 9102 10276 9154
rect 10220 9100 10276 9102
rect 9884 9042 9940 9044
rect 9884 8990 9886 9042
rect 9886 8990 9938 9042
rect 9938 8990 9940 9042
rect 9884 8988 9940 8990
rect 9772 8092 9828 8148
rect 9996 4338 10052 4340
rect 9996 4286 9998 4338
rect 9998 4286 10050 4338
rect 10050 4286 10052 4338
rect 9996 4284 10052 4286
rect 12012 11170 12068 11172
rect 12012 11118 12014 11170
rect 12014 11118 12066 11170
rect 12066 11118 12068 11170
rect 12012 11116 12068 11118
rect 11564 9660 11620 9716
rect 11900 9660 11956 9716
rect 13580 12290 13636 12292
rect 13580 12238 13582 12290
rect 13582 12238 13634 12290
rect 13634 12238 13636 12290
rect 13580 12236 13636 12238
rect 13020 12124 13076 12180
rect 13244 12178 13300 12180
rect 13244 12126 13246 12178
rect 13246 12126 13298 12178
rect 13298 12126 13300 12178
rect 13244 12124 13300 12126
rect 12908 11282 12964 11284
rect 12908 11230 12910 11282
rect 12910 11230 12962 11282
rect 12962 11230 12964 11282
rect 12908 11228 12964 11230
rect 13916 13692 13972 13748
rect 14140 13468 14196 13524
rect 14028 12178 14084 12180
rect 14028 12126 14030 12178
rect 14030 12126 14082 12178
rect 14082 12126 14084 12178
rect 14028 12124 14084 12126
rect 15708 9212 15764 9268
rect 15148 4338 15204 4340
rect 15148 4286 15150 4338
rect 15150 4286 15202 4338
rect 15202 4286 15204 4338
rect 15148 4284 15204 4286
rect 15372 4284 15428 4340
rect 15596 4338 15652 4340
rect 15596 4286 15598 4338
rect 15598 4286 15650 4338
rect 15650 4286 15652 4338
rect 15596 4284 15652 4286
rect 16268 9212 16324 9268
rect 16380 15148 16436 15204
rect 18060 16828 18116 16884
rect 17612 16156 17668 16212
rect 17276 15874 17332 15876
rect 17276 15822 17278 15874
rect 17278 15822 17330 15874
rect 17330 15822 17332 15874
rect 17276 15820 17332 15822
rect 18620 16994 18676 16996
rect 18620 16942 18622 16994
rect 18622 16942 18674 16994
rect 18674 16942 18676 16994
rect 18620 16940 18676 16942
rect 19628 17724 19684 17780
rect 19404 17052 19460 17108
rect 21644 20690 21700 20692
rect 21644 20638 21646 20690
rect 21646 20638 21698 20690
rect 21698 20638 21700 20690
rect 21644 20636 21700 20638
rect 21532 20524 21588 20580
rect 22988 22258 23044 22260
rect 22988 22206 22990 22258
rect 22990 22206 23042 22258
rect 23042 22206 23044 22258
rect 22988 22204 23044 22206
rect 23324 22146 23380 22148
rect 23324 22094 23326 22146
rect 23326 22094 23378 22146
rect 23378 22094 23380 22146
rect 23324 22092 23380 22094
rect 21868 20524 21924 20580
rect 20636 19964 20692 20020
rect 20860 20018 20916 20020
rect 20860 19966 20862 20018
rect 20862 19966 20914 20018
rect 20914 19966 20916 20018
rect 20860 19964 20916 19966
rect 21196 19964 21252 20020
rect 20524 19068 20580 19124
rect 20748 19010 20804 19012
rect 20748 18958 20750 19010
rect 20750 18958 20802 19010
rect 20802 18958 20804 19010
rect 20748 18956 20804 18958
rect 20524 18844 20580 18900
rect 20412 18508 20468 18564
rect 20860 18620 20916 18676
rect 20076 17388 20132 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 18508 16828 18564 16884
rect 18956 16210 19012 16212
rect 18956 16158 18958 16210
rect 18958 16158 19010 16210
rect 19010 16158 19012 16210
rect 18956 16156 19012 16158
rect 17724 15202 17780 15204
rect 17724 15150 17726 15202
rect 17726 15150 17778 15202
rect 17778 15150 17780 15202
rect 17724 15148 17780 15150
rect 19068 16098 19124 16100
rect 19068 16046 19070 16098
rect 19070 16046 19122 16098
rect 19122 16046 19124 16098
rect 19068 16044 19124 16046
rect 18732 15820 18788 15876
rect 17052 4338 17108 4340
rect 17052 4286 17054 4338
rect 17054 4286 17106 4338
rect 17106 4286 17108 4338
rect 17052 4284 17108 4286
rect 17388 4284 17444 4340
rect 17724 4338 17780 4340
rect 17724 4286 17726 4338
rect 17726 4286 17778 4338
rect 17778 4286 17780 4338
rect 17724 4284 17780 4286
rect 19628 16716 19684 16772
rect 19404 16156 19460 16212
rect 19292 15820 19348 15876
rect 19628 15820 19684 15876
rect 19964 15874 20020 15876
rect 19964 15822 19966 15874
rect 19966 15822 20018 15874
rect 20018 15822 20020 15874
rect 19964 15820 20020 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20300 17500 20356 17556
rect 21756 18844 21812 18900
rect 21532 18674 21588 18676
rect 21532 18622 21534 18674
rect 21534 18622 21586 18674
rect 21586 18622 21588 18674
rect 21532 18620 21588 18622
rect 20300 17106 20356 17108
rect 20300 17054 20302 17106
rect 20302 17054 20354 17106
rect 20354 17054 20356 17106
rect 20300 17052 20356 17054
rect 20636 17388 20692 17444
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19852 4338 19908 4340
rect 19852 4286 19854 4338
rect 19854 4286 19906 4338
rect 19906 4286 19908 4338
rect 19852 4284 19908 4286
rect 20300 4338 20356 4340
rect 20300 4286 20302 4338
rect 20302 4286 20354 4338
rect 20354 4286 20356 4338
rect 20300 4284 20356 4286
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21084 17612 21140 17668
rect 21532 17554 21588 17556
rect 21532 17502 21534 17554
rect 21534 17502 21586 17554
rect 21586 17502 21588 17554
rect 21532 17500 21588 17502
rect 20860 17164 20916 17220
rect 21532 16882 21588 16884
rect 21532 16830 21534 16882
rect 21534 16830 21586 16882
rect 21586 16830 21588 16882
rect 21532 16828 21588 16830
rect 22428 20578 22484 20580
rect 22428 20526 22430 20578
rect 22430 20526 22482 20578
rect 22482 20526 22484 20578
rect 22428 20524 22484 20526
rect 22204 19906 22260 19908
rect 22204 19854 22206 19906
rect 22206 19854 22258 19906
rect 22258 19854 22260 19906
rect 22204 19852 22260 19854
rect 21980 19122 22036 19124
rect 21980 19070 21982 19122
rect 21982 19070 22034 19122
rect 22034 19070 22036 19122
rect 21980 19068 22036 19070
rect 21980 18844 22036 18900
rect 20748 16716 20804 16772
rect 21196 4338 21252 4340
rect 21196 4286 21198 4338
rect 21198 4286 21250 4338
rect 21250 4286 21252 4338
rect 21196 4284 21252 4286
rect 21420 4284 21476 4340
rect 21644 4338 21700 4340
rect 21644 4286 21646 4338
rect 21646 4286 21698 4338
rect 21698 4286 21700 4338
rect 21644 4284 21700 4286
rect 21644 3554 21700 3556
rect 21644 3502 21646 3554
rect 21646 3502 21698 3554
rect 21698 3502 21700 3554
rect 21644 3500 21700 3502
rect 22428 16828 22484 16884
rect 22316 16770 22372 16772
rect 22316 16718 22318 16770
rect 22318 16718 22370 16770
rect 22370 16718 22372 16770
rect 22316 16716 22372 16718
rect 23100 20524 23156 20580
rect 23548 20578 23604 20580
rect 23548 20526 23550 20578
rect 23550 20526 23602 20578
rect 23602 20526 23604 20578
rect 23548 20524 23604 20526
rect 23660 20412 23716 20468
rect 22876 19906 22932 19908
rect 22876 19854 22878 19906
rect 22878 19854 22930 19906
rect 22930 19854 22932 19906
rect 22876 19852 22932 19854
rect 24780 23154 24836 23156
rect 24780 23102 24782 23154
rect 24782 23102 24834 23154
rect 24834 23102 24836 23154
rect 24780 23100 24836 23102
rect 23996 21698 24052 21700
rect 23996 21646 23998 21698
rect 23998 21646 24050 21698
rect 24050 21646 24052 21698
rect 23996 21644 24052 21646
rect 23212 17276 23268 17332
rect 22652 16828 22708 16884
rect 22988 16882 23044 16884
rect 22988 16830 22990 16882
rect 22990 16830 23042 16882
rect 23042 16830 23044 16882
rect 22988 16828 23044 16830
rect 23100 16658 23156 16660
rect 23100 16606 23102 16658
rect 23102 16606 23154 16658
rect 23154 16606 23156 16658
rect 23100 16604 23156 16606
rect 23324 16770 23380 16772
rect 23324 16718 23326 16770
rect 23326 16718 23378 16770
rect 23378 16718 23380 16770
rect 23324 16716 23380 16718
rect 25788 23714 25844 23716
rect 25788 23662 25790 23714
rect 25790 23662 25842 23714
rect 25842 23662 25844 23714
rect 25788 23660 25844 23662
rect 26012 23548 26068 23604
rect 25452 17500 25508 17556
rect 24332 17052 24388 17108
rect 24892 17052 24948 17108
rect 23884 16604 23940 16660
rect 22652 16098 22708 16100
rect 22652 16046 22654 16098
rect 22654 16046 22706 16098
rect 22706 16046 22708 16098
rect 22652 16044 22708 16046
rect 24444 16882 24500 16884
rect 24444 16830 24446 16882
rect 24446 16830 24498 16882
rect 24498 16830 24500 16882
rect 24444 16828 24500 16830
rect 22092 3500 22148 3556
rect 22428 3500 22484 3556
rect 23884 4338 23940 4340
rect 23884 4286 23886 4338
rect 23886 4286 23938 4338
rect 23938 4286 23940 4338
rect 23884 4284 23940 4286
rect 24108 4284 24164 4340
rect 24332 4338 24388 4340
rect 24332 4286 24334 4338
rect 24334 4286 24386 4338
rect 24386 4286 24388 4338
rect 24332 4284 24388 4286
rect 25788 17554 25844 17556
rect 25788 17502 25790 17554
rect 25790 17502 25842 17554
rect 25842 17502 25844 17554
rect 25788 17500 25844 17502
rect 26012 17442 26068 17444
rect 26012 17390 26014 17442
rect 26014 17390 26066 17442
rect 26066 17390 26068 17442
rect 26012 17388 26068 17390
rect 26012 17164 26068 17220
rect 25788 17052 25844 17108
rect 25676 16882 25732 16884
rect 25676 16830 25678 16882
rect 25678 16830 25730 16882
rect 25730 16830 25732 16882
rect 25676 16828 25732 16830
rect 26460 25340 26516 25396
rect 26348 23548 26404 23604
rect 26236 17388 26292 17444
rect 25900 4338 25956 4340
rect 25900 4286 25902 4338
rect 25902 4286 25954 4338
rect 25954 4286 25956 4338
rect 25900 4284 25956 4286
rect 26124 4284 26180 4340
rect 26348 4338 26404 4340
rect 26348 4286 26350 4338
rect 26350 4286 26402 4338
rect 26402 4286 26404 4338
rect 26348 4284 26404 4286
rect 27132 25394 27188 25396
rect 27132 25342 27134 25394
rect 27134 25342 27186 25394
rect 27186 25342 27188 25394
rect 27132 25340 27188 25342
rect 26684 25282 26740 25284
rect 26684 25230 26686 25282
rect 26686 25230 26738 25282
rect 26738 25230 26740 25282
rect 26684 25228 26740 25230
rect 27020 24610 27076 24612
rect 27020 24558 27022 24610
rect 27022 24558 27074 24610
rect 27074 24558 27076 24610
rect 27020 24556 27076 24558
rect 26684 23826 26740 23828
rect 26684 23774 26686 23826
rect 26686 23774 26738 23826
rect 26738 23774 26740 23826
rect 26684 23772 26740 23774
rect 27020 17554 27076 17556
rect 27020 17502 27022 17554
rect 27022 17502 27074 17554
rect 27074 17502 27076 17554
rect 27020 17500 27076 17502
rect 26572 17442 26628 17444
rect 26572 17390 26574 17442
rect 26574 17390 26626 17442
rect 26626 17390 26628 17442
rect 26572 17388 26628 17390
rect 26684 16882 26740 16884
rect 26684 16830 26686 16882
rect 26686 16830 26738 16882
rect 26738 16830 26740 16882
rect 26684 16828 26740 16830
rect 28028 26962 28084 26964
rect 28028 26910 28030 26962
rect 28030 26910 28082 26962
rect 28082 26910 28084 26962
rect 28028 26908 28084 26910
rect 28364 26850 28420 26852
rect 28364 26798 28366 26850
rect 28366 26798 28418 26850
rect 28418 26798 28420 26850
rect 28364 26796 28420 26798
rect 27692 26402 27748 26404
rect 27692 26350 27694 26402
rect 27694 26350 27746 26402
rect 27746 26350 27748 26402
rect 27692 26348 27748 26350
rect 27580 25506 27636 25508
rect 27580 25454 27582 25506
rect 27582 25454 27634 25506
rect 27634 25454 27636 25506
rect 27580 25452 27636 25454
rect 27356 25340 27412 25396
rect 28812 26962 28868 26964
rect 28812 26910 28814 26962
rect 28814 26910 28866 26962
rect 28866 26910 28868 26962
rect 28812 26908 28868 26910
rect 29932 28418 29988 28420
rect 29932 28366 29934 28418
rect 29934 28366 29986 28418
rect 29986 28366 29988 28418
rect 29932 28364 29988 28366
rect 29820 27858 29876 27860
rect 29820 27806 29822 27858
rect 29822 27806 29874 27858
rect 29874 27806 29876 27858
rect 29820 27804 29876 27806
rect 30156 4284 30212 4340
rect 30380 28642 30436 28644
rect 30380 28590 30382 28642
rect 30382 28590 30434 28642
rect 30434 28590 30436 28642
rect 30380 28588 30436 28590
rect 30604 29372 30660 29428
rect 31612 30098 31668 30100
rect 31612 30046 31614 30098
rect 31614 30046 31666 30098
rect 31666 30046 31668 30098
rect 31612 30044 31668 30046
rect 32620 31666 32676 31668
rect 32620 31614 32622 31666
rect 32622 31614 32674 31666
rect 32674 31614 32676 31666
rect 32620 31612 32676 31614
rect 32284 31106 32340 31108
rect 32284 31054 32286 31106
rect 32286 31054 32338 31106
rect 32338 31054 32340 31106
rect 32284 31052 32340 31054
rect 32956 31554 33012 31556
rect 32956 31502 32958 31554
rect 32958 31502 33010 31554
rect 33010 31502 33012 31554
rect 32956 31500 33012 31502
rect 32732 30994 32788 30996
rect 32732 30942 32734 30994
rect 32734 30942 32786 30994
rect 32786 30942 32788 30994
rect 32732 30940 32788 30942
rect 30380 4338 30436 4340
rect 30380 4286 30382 4338
rect 30382 4286 30434 4338
rect 30434 4286 30436 4338
rect 30380 4284 30436 4286
rect 31948 4284 32004 4340
rect 32396 4338 32452 4340
rect 32396 4286 32398 4338
rect 32398 4286 32450 4338
rect 32450 4286 32452 4338
rect 32396 4284 32452 4286
rect 33628 32562 33684 32564
rect 33628 32510 33630 32562
rect 33630 32510 33682 32562
rect 33682 32510 33684 32562
rect 33628 32508 33684 32510
rect 33852 31666 33908 31668
rect 33852 31614 33854 31666
rect 33854 31614 33906 31666
rect 33906 31614 33908 31666
rect 33852 31612 33908 31614
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 36988 35810 37044 35812
rect 36988 35758 36990 35810
rect 36990 35758 37042 35810
rect 37042 35758 37044 35810
rect 36988 35756 37044 35758
rect 36316 34802 36372 34804
rect 36316 34750 36318 34802
rect 36318 34750 36370 34802
rect 36370 34750 36372 34802
rect 36316 34748 36372 34750
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35084 3330 35140 3332
rect 35084 3278 35086 3330
rect 35086 3278 35138 3330
rect 35138 3278 35140 3330
rect 35084 3276 35140 3278
rect 36092 3276 36148 3332
rect 37996 37100 38052 37156
rect 39004 37826 39060 37828
rect 39004 37774 39006 37826
rect 39006 37774 39058 37826
rect 39058 37774 39060 37826
rect 39004 37772 39060 37774
rect 38332 37100 38388 37156
rect 37548 36370 37604 36372
rect 37548 36318 37550 36370
rect 37550 36318 37602 36370
rect 37602 36318 37604 36370
rect 37548 36316 37604 36318
rect 37436 35698 37492 35700
rect 37436 35646 37438 35698
rect 37438 35646 37490 35698
rect 37490 35646 37492 35698
rect 37436 35644 37492 35646
rect 37884 36258 37940 36260
rect 37884 36206 37886 36258
rect 37886 36206 37938 36258
rect 37938 36206 37940 36258
rect 37884 36204 37940 36206
rect 38780 36370 38836 36372
rect 38780 36318 38782 36370
rect 38782 36318 38834 36370
rect 38834 36318 38836 36370
rect 38780 36316 38836 36318
rect 39676 39506 39732 39508
rect 39676 39454 39678 39506
rect 39678 39454 39730 39506
rect 39730 39454 39732 39506
rect 39676 39452 39732 39454
rect 39788 38946 39844 38948
rect 39788 38894 39790 38946
rect 39790 38894 39842 38946
rect 39842 38894 39844 38946
rect 39788 38892 39844 38894
rect 39564 38834 39620 38836
rect 39564 38782 39566 38834
rect 39566 38782 39618 38834
rect 39618 38782 39620 38834
rect 39564 38780 39620 38782
rect 39452 37938 39508 37940
rect 39452 37886 39454 37938
rect 39454 37886 39506 37938
rect 39506 37886 39508 37938
rect 39452 37884 39508 37886
rect 40572 40402 40628 40404
rect 40572 40350 40574 40402
rect 40574 40350 40626 40402
rect 40626 40350 40628 40402
rect 40572 40348 40628 40350
rect 41580 40402 41636 40404
rect 41580 40350 41582 40402
rect 41582 40350 41634 40402
rect 41634 40350 41636 40402
rect 41580 40348 41636 40350
rect 40012 39394 40068 39396
rect 40012 39342 40014 39394
rect 40014 39342 40066 39394
rect 40066 39342 40068 39394
rect 40012 39340 40068 39342
rect 40908 39506 40964 39508
rect 40908 39454 40910 39506
rect 40910 39454 40962 39506
rect 40962 39454 40964 39506
rect 40908 39452 40964 39454
rect 40684 38834 40740 38836
rect 40684 38782 40686 38834
rect 40686 38782 40738 38834
rect 40738 38782 40740 38834
rect 40684 38780 40740 38782
rect 38668 4338 38724 4340
rect 38668 4286 38670 4338
rect 38670 4286 38722 4338
rect 38722 4286 38724 4338
rect 38668 4284 38724 4286
rect 38892 4284 38948 4340
rect 39116 4338 39172 4340
rect 39116 4286 39118 4338
rect 39118 4286 39170 4338
rect 39170 4286 39172 4338
rect 39116 4284 39172 4286
rect 40908 4284 40964 4340
rect 41580 4338 41636 4340
rect 41580 4286 41582 4338
rect 41582 4286 41634 4338
rect 41634 4286 41636 4338
rect 41580 4284 41636 4286
rect 42812 40962 42868 40964
rect 42812 40910 42814 40962
rect 42814 40910 42866 40962
rect 42866 40910 42868 40962
rect 42812 40908 42868 40910
rect 42364 40402 42420 40404
rect 42364 40350 42366 40402
rect 42366 40350 42418 40402
rect 42418 40350 42420 40402
rect 42364 40348 42420 40350
rect 43484 41858 43540 41860
rect 43484 41806 43486 41858
rect 43486 41806 43538 41858
rect 43538 41806 43540 41858
rect 43484 41804 43540 41806
rect 43932 41858 43988 41860
rect 43932 41806 43934 41858
rect 43934 41806 43986 41858
rect 43986 41806 43988 41858
rect 43932 41804 43988 41806
rect 43036 40908 43092 40964
rect 42924 3500 42980 3556
rect 43596 3554 43652 3556
rect 43596 3502 43598 3554
rect 43598 3502 43650 3554
rect 43650 3502 43652 3554
rect 43596 3500 43652 3502
rect 44828 43426 44884 43428
rect 44828 43374 44830 43426
rect 44830 43374 44882 43426
rect 44882 43374 44884 43426
rect 44828 43372 44884 43374
rect 45500 44210 45556 44212
rect 45500 44158 45502 44210
rect 45502 44158 45554 44210
rect 45554 44158 45556 44210
rect 45500 44156 45556 44158
rect 45836 44210 45892 44212
rect 45836 44158 45838 44210
rect 45838 44158 45890 44210
rect 45890 44158 45892 44210
rect 45836 44156 45892 44158
rect 46732 44098 46788 44100
rect 46732 44046 46734 44098
rect 46734 44046 46786 44098
rect 46786 44046 46788 44098
rect 46732 44044 46788 44046
rect 44268 3500 44324 3556
rect 44940 3554 44996 3556
rect 44940 3502 44942 3554
rect 44942 3502 44994 3554
rect 44994 3502 44996 3554
rect 44940 3500 44996 3502
rect 45052 3388 45108 3444
rect 46060 4284 46116 4340
rect 45612 3388 45668 3444
rect 45948 3388 46004 3444
rect 47180 45778 47236 45780
rect 47180 45726 47182 45778
rect 47182 45726 47234 45778
rect 47234 45726 47236 45778
rect 47180 45724 47236 45726
rect 46956 45052 47012 45108
rect 47740 45890 47796 45892
rect 47740 45838 47742 45890
rect 47742 45838 47794 45890
rect 47794 45838 47796 45890
rect 47740 45836 47796 45838
rect 48076 45890 48132 45892
rect 48076 45838 48078 45890
rect 48078 45838 48130 45890
rect 48130 45838 48132 45890
rect 48076 45836 48132 45838
rect 46508 4338 46564 4340
rect 46508 4286 46510 4338
rect 46510 4286 46562 4338
rect 46562 4286 46564 4338
rect 46508 4284 46564 4286
rect 46956 3500 47012 3556
rect 47068 3388 47124 3444
rect 48972 47346 49028 47348
rect 48972 47294 48974 47346
rect 48974 47294 49026 47346
rect 49026 47294 49028 47346
rect 48972 47292 49028 47294
rect 48524 47234 48580 47236
rect 48524 47182 48526 47234
rect 48526 47182 48578 47234
rect 48578 47182 48580 47234
rect 48524 47180 48580 47182
rect 48300 46562 48356 46564
rect 48300 46510 48302 46562
rect 48302 46510 48354 46562
rect 48354 46510 48356 46562
rect 48300 46508 48356 46510
rect 49420 48802 49476 48804
rect 49420 48750 49422 48802
rect 49422 48750 49474 48802
rect 49474 48750 49476 48802
rect 49420 48748 49476 48750
rect 49980 49196 50036 49252
rect 49868 49026 49924 49028
rect 49868 48974 49870 49026
rect 49870 48974 49922 49026
rect 49922 48974 49924 49026
rect 49868 48972 49924 48974
rect 49868 48748 49924 48804
rect 51772 50316 51828 50372
rect 50876 49644 50932 49700
rect 50988 50092 51044 50148
rect 50428 49532 50484 49588
rect 51212 50034 51268 50036
rect 51212 49982 51214 50034
rect 51214 49982 51266 50034
rect 51266 49982 51268 50034
rect 51212 49980 51268 49982
rect 50988 49532 51044 49588
rect 50316 49420 50372 49476
rect 50428 49026 50484 49028
rect 50428 48974 50430 49026
rect 50430 48974 50482 49026
rect 50482 48974 50484 49026
rect 50428 48972 50484 48974
rect 51436 49698 51492 49700
rect 51436 49646 51438 49698
rect 51438 49646 51490 49698
rect 51490 49646 51492 49698
rect 51436 49644 51492 49646
rect 51660 49586 51716 49588
rect 51660 49534 51662 49586
rect 51662 49534 51714 49586
rect 51714 49534 51716 49586
rect 51660 49532 51716 49534
rect 50316 48748 50372 48804
rect 50540 48748 50596 48804
rect 51100 48802 51156 48804
rect 51100 48750 51102 48802
rect 51102 48750 51154 48802
rect 51154 48750 51156 48802
rect 51100 48748 51156 48750
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 50316 5852 50372 5908
rect 49980 5234 50036 5236
rect 49980 5182 49982 5234
rect 49982 5182 50034 5234
rect 50034 5182 50036 5234
rect 49980 5180 50036 5182
rect 47964 4172 48020 4228
rect 48636 4226 48692 4228
rect 48636 4174 48638 4226
rect 48638 4174 48690 4226
rect 48690 4174 48692 4226
rect 48636 4172 48692 4174
rect 48972 4172 49028 4228
rect 47964 3554 48020 3556
rect 47964 3502 47966 3554
rect 47966 3502 48018 3554
rect 48018 3502 48020 3554
rect 47964 3500 48020 3502
rect 48300 3388 48356 3444
rect 50876 5180 50932 5236
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 50204 4226 50260 4228
rect 50204 4174 50206 4226
rect 50206 4174 50258 4226
rect 50258 4174 50260 4226
rect 50204 4172 50260 4174
rect 50316 3500 50372 3556
rect 49196 3442 49252 3444
rect 49196 3390 49198 3442
rect 49198 3390 49250 3442
rect 49250 3390 49252 3442
rect 49196 3388 49252 3390
rect 49644 3388 49700 3444
rect 51772 5234 51828 5236
rect 51772 5182 51774 5234
rect 51774 5182 51826 5234
rect 51826 5182 51828 5234
rect 51772 5180 51828 5182
rect 52556 52220 52612 52276
rect 52668 51436 52724 51492
rect 52332 50594 52388 50596
rect 52332 50542 52334 50594
rect 52334 50542 52386 50594
rect 52386 50542 52388 50594
rect 52332 50540 52388 50542
rect 53116 52834 53172 52836
rect 53116 52782 53118 52834
rect 53118 52782 53170 52834
rect 53170 52782 53172 52834
rect 53116 52780 53172 52782
rect 54460 53116 54516 53172
rect 54684 53730 54740 53732
rect 54684 53678 54686 53730
rect 54686 53678 54738 53730
rect 54738 53678 54740 53730
rect 54684 53676 54740 53678
rect 55356 55074 55412 55076
rect 55356 55022 55358 55074
rect 55358 55022 55410 55074
rect 55410 55022 55412 55074
rect 55356 55020 55412 55022
rect 55020 54514 55076 54516
rect 55020 54462 55022 54514
rect 55022 54462 55074 54514
rect 55074 54462 55076 54514
rect 55020 54460 55076 54462
rect 55356 54348 55412 54404
rect 55244 54290 55300 54292
rect 55244 54238 55246 54290
rect 55246 54238 55298 54290
rect 55298 54238 55300 54290
rect 55244 54236 55300 54238
rect 55132 54124 55188 54180
rect 54908 53730 54964 53732
rect 54908 53678 54910 53730
rect 54910 53678 54962 53730
rect 54962 53678 54964 53730
rect 54908 53676 54964 53678
rect 54348 53058 54404 53060
rect 54348 53006 54350 53058
rect 54350 53006 54402 53058
rect 54402 53006 54404 53058
rect 54348 53004 54404 53006
rect 54124 52834 54180 52836
rect 54124 52782 54126 52834
rect 54126 52782 54178 52834
rect 54178 52782 54180 52834
rect 54124 52780 54180 52782
rect 53340 52722 53396 52724
rect 53340 52670 53342 52722
rect 53342 52670 53394 52722
rect 53394 52670 53396 52722
rect 53340 52668 53396 52670
rect 53228 51884 53284 51940
rect 53676 51548 53732 51604
rect 53452 50092 53508 50148
rect 52220 49586 52276 49588
rect 52220 49534 52222 49586
rect 52222 49534 52274 49586
rect 52274 49534 52276 49586
rect 52220 49532 52276 49534
rect 52668 6076 52724 6132
rect 54012 17442 54068 17444
rect 54012 17390 54014 17442
rect 54014 17390 54066 17442
rect 54066 17390 54068 17442
rect 54012 17388 54068 17390
rect 53564 17052 53620 17108
rect 53900 15260 53956 15316
rect 53452 14418 53508 14420
rect 53452 14366 53454 14418
rect 53454 14366 53506 14418
rect 53506 14366 53508 14418
rect 53452 14364 53508 14366
rect 54572 18396 54628 18452
rect 54460 16882 54516 16884
rect 54460 16830 54462 16882
rect 54462 16830 54514 16882
rect 54514 16830 54516 16882
rect 54460 16828 54516 16830
rect 54572 17164 54628 17220
rect 54796 18508 54852 18564
rect 55020 18338 55076 18340
rect 55020 18286 55022 18338
rect 55022 18286 55074 18338
rect 55074 18286 55076 18338
rect 55020 18284 55076 18286
rect 55132 17164 55188 17220
rect 55020 17052 55076 17108
rect 55244 16828 55300 16884
rect 54796 15260 54852 15316
rect 55020 15314 55076 15316
rect 55020 15262 55022 15314
rect 55022 15262 55074 15314
rect 55074 15262 55076 15314
rect 55020 15260 55076 15262
rect 54348 13468 54404 13524
rect 54236 6130 54292 6132
rect 54236 6078 54238 6130
rect 54238 6078 54290 6130
rect 54290 6078 54292 6130
rect 54236 6076 54292 6078
rect 52332 5292 52388 5348
rect 52668 5180 52724 5236
rect 51660 3724 51716 3780
rect 50988 3612 51044 3668
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 51548 3442 51604 3444
rect 51548 3390 51550 3442
rect 51550 3390 51602 3442
rect 51602 3390 51604 3442
rect 51548 3388 51604 3390
rect 52108 3500 52164 3556
rect 53116 5292 53172 5348
rect 53564 5180 53620 5236
rect 53452 3666 53508 3668
rect 53452 3614 53454 3666
rect 53454 3614 53506 3666
rect 53506 3614 53508 3666
rect 53452 3612 53508 3614
rect 52332 3388 52388 3444
rect 54124 5234 54180 5236
rect 54124 5182 54126 5234
rect 54126 5182 54178 5234
rect 54178 5182 54180 5234
rect 54124 5180 54180 5182
rect 54572 14140 54628 14196
rect 55020 14364 55076 14420
rect 54796 14252 54852 14308
rect 54908 13468 54964 13524
rect 55244 13468 55300 13524
rect 56812 56252 56868 56308
rect 56252 56140 56308 56196
rect 55580 55132 55636 55188
rect 56700 55970 56756 55972
rect 56700 55918 56702 55970
rect 56702 55918 56754 55970
rect 56754 55918 56756 55970
rect 56700 55916 56756 55918
rect 56924 55244 56980 55300
rect 57260 55186 57316 55188
rect 57260 55134 57262 55186
rect 57262 55134 57314 55186
rect 57314 55134 57316 55186
rect 57260 55132 57316 55134
rect 55804 54908 55860 54964
rect 56924 55020 56980 55076
rect 56476 54908 56532 54964
rect 56588 54796 56644 54852
rect 55580 54460 55636 54516
rect 55804 54290 55860 54292
rect 55804 54238 55806 54290
rect 55806 54238 55858 54290
rect 55858 54238 55860 54290
rect 55804 54236 55860 54238
rect 55580 53676 55636 53732
rect 55916 53730 55972 53732
rect 55916 53678 55918 53730
rect 55918 53678 55970 53730
rect 55970 53678 55972 53730
rect 55916 53676 55972 53678
rect 56140 53676 56196 53732
rect 56028 52892 56084 52948
rect 56140 51602 56196 51604
rect 56140 51550 56142 51602
rect 56142 51550 56194 51602
rect 56194 51550 56196 51602
rect 56140 51548 56196 51550
rect 56252 52162 56308 52164
rect 56252 52110 56254 52162
rect 56254 52110 56306 52162
rect 56306 52110 56308 52162
rect 56252 52108 56308 52110
rect 55692 51324 55748 51380
rect 55580 18562 55636 18564
rect 55580 18510 55582 18562
rect 55582 18510 55634 18562
rect 55634 18510 55636 18562
rect 55580 18508 55636 18510
rect 56364 51378 56420 51380
rect 56364 51326 56366 51378
rect 56366 51326 56418 51378
rect 56418 51326 56420 51378
rect 56364 51324 56420 51326
rect 56028 18450 56084 18452
rect 56028 18398 56030 18450
rect 56030 18398 56082 18450
rect 56082 18398 56084 18450
rect 56028 18396 56084 18398
rect 55804 18284 55860 18340
rect 55468 17388 55524 17444
rect 56028 17388 56084 17444
rect 55916 15426 55972 15428
rect 55916 15374 55918 15426
rect 55918 15374 55970 15426
rect 55970 15374 55972 15426
rect 55916 15372 55972 15374
rect 55580 15314 55636 15316
rect 55580 15262 55582 15314
rect 55582 15262 55634 15314
rect 55634 15262 55636 15314
rect 55580 15260 55636 15262
rect 56140 15148 56196 15204
rect 55916 14530 55972 14532
rect 55916 14478 55918 14530
rect 55918 14478 55970 14530
rect 55970 14478 55972 14530
rect 55916 14476 55972 14478
rect 55580 13858 55636 13860
rect 55580 13806 55582 13858
rect 55582 13806 55634 13858
rect 55634 13806 55636 13858
rect 55580 13804 55636 13806
rect 55468 13692 55524 13748
rect 54572 6188 54628 6244
rect 54460 4284 54516 4340
rect 54684 6076 54740 6132
rect 53676 4172 53732 4228
rect 53788 3724 53844 3780
rect 54348 3612 54404 3668
rect 54908 6076 54964 6132
rect 56924 54572 56980 54628
rect 57148 53676 57204 53732
rect 56588 52892 56644 52948
rect 56588 52722 56644 52724
rect 56588 52670 56590 52722
rect 56590 52670 56642 52722
rect 56642 52670 56644 52722
rect 56588 52668 56644 52670
rect 56812 52162 56868 52164
rect 56812 52110 56814 52162
rect 56814 52110 56866 52162
rect 56866 52110 56868 52162
rect 56812 52108 56868 52110
rect 57260 52162 57316 52164
rect 57260 52110 57262 52162
rect 57262 52110 57314 52162
rect 57314 52110 57316 52162
rect 57260 52108 57316 52110
rect 57148 51324 57204 51380
rect 58156 57484 58212 57540
rect 58044 56924 58100 56980
rect 58268 57426 58324 57428
rect 58268 57374 58270 57426
rect 58270 57374 58322 57426
rect 58322 57374 58324 57426
rect 58268 57372 58324 57374
rect 57820 56306 57876 56308
rect 57820 56254 57822 56306
rect 57822 56254 57874 56306
rect 57874 56254 57876 56306
rect 57820 56252 57876 56254
rect 57708 55244 57764 55300
rect 57708 55074 57764 55076
rect 57708 55022 57710 55074
rect 57710 55022 57762 55074
rect 57762 55022 57764 55074
rect 57708 55020 57764 55022
rect 57596 54796 57652 54852
rect 57820 53170 57876 53172
rect 57820 53118 57822 53170
rect 57822 53118 57874 53170
rect 57874 53118 57876 53170
rect 57820 53116 57876 53118
rect 57484 52108 57540 52164
rect 57820 51602 57876 51604
rect 57820 51550 57822 51602
rect 57822 51550 57874 51602
rect 57874 51550 57876 51602
rect 57820 51548 57876 51550
rect 57484 51378 57540 51380
rect 57484 51326 57486 51378
rect 57486 51326 57538 51378
rect 57538 51326 57540 51378
rect 57484 51324 57540 51326
rect 56588 17442 56644 17444
rect 56588 17390 56590 17442
rect 56590 17390 56642 17442
rect 56642 17390 56644 17442
rect 56588 17388 56644 17390
rect 56588 14530 56644 14532
rect 56588 14478 56590 14530
rect 56590 14478 56642 14530
rect 56642 14478 56644 14530
rect 56588 14476 56644 14478
rect 56700 13746 56756 13748
rect 56700 13694 56702 13746
rect 56702 13694 56754 13746
rect 56754 13694 56756 13746
rect 56700 13692 56756 13694
rect 57484 13746 57540 13748
rect 57484 13694 57486 13746
rect 57486 13694 57538 13746
rect 57538 13694 57540 13746
rect 57484 13692 57540 13694
rect 56476 6300 56532 6356
rect 57372 6188 57428 6244
rect 55020 5180 55076 5236
rect 56364 6076 56420 6132
rect 57820 13692 57876 13748
rect 58268 56082 58324 56084
rect 58268 56030 58270 56082
rect 58270 56030 58322 56082
rect 58322 56030 58324 56082
rect 58268 56028 58324 56030
rect 58044 55132 58100 55188
rect 58828 60674 58884 60676
rect 58828 60622 58830 60674
rect 58830 60622 58882 60674
rect 58882 60622 58884 60674
rect 58828 60620 58884 60622
rect 59388 60620 59444 60676
rect 60620 60898 60676 60900
rect 60620 60846 60622 60898
rect 60622 60846 60674 60898
rect 60674 60846 60676 60898
rect 60620 60844 60676 60846
rect 60956 60844 61012 60900
rect 60844 60786 60900 60788
rect 60844 60734 60846 60786
rect 60846 60734 60898 60786
rect 60898 60734 60900 60786
rect 60844 60732 60900 60734
rect 59724 60620 59780 60676
rect 60396 60620 60452 60676
rect 59948 60060 60004 60116
rect 58716 59724 58772 59780
rect 59276 59778 59332 59780
rect 59276 59726 59278 59778
rect 59278 59726 59330 59778
rect 59330 59726 59332 59778
rect 59276 59724 59332 59726
rect 59612 59330 59668 59332
rect 59612 59278 59614 59330
rect 59614 59278 59666 59330
rect 59666 59278 59668 59330
rect 59612 59276 59668 59278
rect 60172 59890 60228 59892
rect 60172 59838 60174 59890
rect 60174 59838 60226 59890
rect 60226 59838 60228 59890
rect 60172 59836 60228 59838
rect 59948 59276 60004 59332
rect 60284 59724 60340 59780
rect 59388 58546 59444 58548
rect 59388 58494 59390 58546
rect 59390 58494 59442 58546
rect 59442 58494 59444 58546
rect 59388 58492 59444 58494
rect 58492 58434 58548 58436
rect 58492 58382 58494 58434
rect 58494 58382 58546 58434
rect 58546 58382 58548 58434
rect 58492 58380 58548 58382
rect 58492 57820 58548 57876
rect 59276 57820 59332 57876
rect 59500 57932 59556 57988
rect 59276 57650 59332 57652
rect 59276 57598 59278 57650
rect 59278 57598 59330 57650
rect 59330 57598 59332 57650
rect 59276 57596 59332 57598
rect 59052 57538 59108 57540
rect 59052 57486 59054 57538
rect 59054 57486 59106 57538
rect 59106 57486 59108 57538
rect 59052 57484 59108 57486
rect 58604 57260 58660 57316
rect 58380 53116 58436 53172
rect 58492 55244 58548 55300
rect 59164 57148 59220 57204
rect 59052 56028 59108 56084
rect 58716 55970 58772 55972
rect 58716 55918 58718 55970
rect 58718 55918 58770 55970
rect 58770 55918 58772 55970
rect 58716 55916 58772 55918
rect 59164 52274 59220 52276
rect 59164 52222 59166 52274
rect 59166 52222 59218 52274
rect 59218 52222 59220 52274
rect 59164 52220 59220 52222
rect 59276 52162 59332 52164
rect 59276 52110 59278 52162
rect 59278 52110 59330 52162
rect 59330 52110 59332 52162
rect 59276 52108 59332 52110
rect 58604 51548 58660 51604
rect 60060 59106 60116 59108
rect 60060 59054 60062 59106
rect 60062 59054 60114 59106
rect 60114 59054 60116 59106
rect 60060 59052 60116 59054
rect 59948 58434 60004 58436
rect 59948 58382 59950 58434
rect 59950 58382 60002 58434
rect 60002 58382 60004 58434
rect 59948 58380 60004 58382
rect 59388 51100 59444 51156
rect 59836 58156 59892 58212
rect 59836 57148 59892 57204
rect 57932 6636 57988 6692
rect 55916 5234 55972 5236
rect 55916 5182 55918 5234
rect 55918 5182 55970 5234
rect 55970 5182 55972 5234
rect 55916 5180 55972 5182
rect 55916 4338 55972 4340
rect 55916 4286 55918 4338
rect 55918 4286 55970 4338
rect 55970 4286 55972 4338
rect 55916 4284 55972 4286
rect 55132 4226 55188 4228
rect 55132 4174 55134 4226
rect 55134 4174 55186 4226
rect 55186 4174 55188 4226
rect 55132 4172 55188 4174
rect 55244 3388 55300 3444
rect 55692 3500 55748 3556
rect 56588 4338 56644 4340
rect 56588 4286 56590 4338
rect 56590 4286 56642 4338
rect 56642 4286 56644 4338
rect 56588 4284 56644 4286
rect 56364 3388 56420 3444
rect 57708 6076 57764 6132
rect 58156 6300 58212 6356
rect 59836 52162 59892 52164
rect 59836 52110 59838 52162
rect 59838 52110 59890 52162
rect 59890 52110 59892 52162
rect 59836 52108 59892 52110
rect 60620 60002 60676 60004
rect 60620 59950 60622 60002
rect 60622 59950 60674 60002
rect 60674 59950 60676 60002
rect 60620 59948 60676 59950
rect 60396 59052 60452 59108
rect 60396 58546 60452 58548
rect 60396 58494 60398 58546
rect 60398 58494 60450 58546
rect 60450 58494 60452 58546
rect 60396 58492 60452 58494
rect 60284 52386 60340 52388
rect 60284 52334 60286 52386
rect 60286 52334 60338 52386
rect 60338 52334 60340 52386
rect 60284 52332 60340 52334
rect 60396 52274 60452 52276
rect 60396 52222 60398 52274
rect 60398 52222 60450 52274
rect 60450 52222 60452 52274
rect 60396 52220 60452 52222
rect 60172 51100 60228 51156
rect 59836 6300 59892 6356
rect 59612 6188 59668 6244
rect 59164 6130 59220 6132
rect 59164 6078 59166 6130
rect 59166 6078 59218 6130
rect 59218 6078 59220 6130
rect 59164 6076 59220 6078
rect 57708 4172 57764 4228
rect 57372 3666 57428 3668
rect 57372 3614 57374 3666
rect 57374 3614 57426 3666
rect 57426 3614 57428 3666
rect 57372 3612 57428 3614
rect 58156 3500 58212 3556
rect 58380 3612 58436 3668
rect 61740 60732 61796 60788
rect 61068 60674 61124 60676
rect 61068 60622 61070 60674
rect 61070 60622 61122 60674
rect 61122 60622 61124 60674
rect 61068 60620 61124 60622
rect 61292 60562 61348 60564
rect 61292 60510 61294 60562
rect 61294 60510 61346 60562
rect 61346 60510 61348 60562
rect 61292 60508 61348 60510
rect 60956 60060 61012 60116
rect 61516 60172 61572 60228
rect 61404 59778 61460 59780
rect 61404 59726 61406 59778
rect 61406 59726 61458 59778
rect 61458 59726 61460 59778
rect 61404 59724 61460 59726
rect 62300 61010 62356 61012
rect 62300 60958 62302 61010
rect 62302 60958 62354 61010
rect 62354 60958 62356 61010
rect 62300 60956 62356 60958
rect 62524 60898 62580 60900
rect 62524 60846 62526 60898
rect 62526 60846 62578 60898
rect 62578 60846 62580 60898
rect 62524 60844 62580 60846
rect 62076 60674 62132 60676
rect 62076 60622 62078 60674
rect 62078 60622 62130 60674
rect 62130 60622 62132 60674
rect 62076 60620 62132 60622
rect 62076 60172 62132 60228
rect 61292 57260 61348 57316
rect 61404 52274 61460 52276
rect 61404 52222 61406 52274
rect 61406 52222 61458 52274
rect 61458 52222 61460 52274
rect 61404 52220 61460 52222
rect 60172 6076 60228 6132
rect 59388 3442 59444 3444
rect 59388 3390 59390 3442
rect 59390 3390 59442 3442
rect 59442 3390 59444 3442
rect 59388 3388 59444 3390
rect 60284 6636 60340 6692
rect 61068 6188 61124 6244
rect 59948 4226 60004 4228
rect 59948 4174 59950 4226
rect 59950 4174 60002 4226
rect 60002 4174 60004 4226
rect 59948 4172 60004 4174
rect 59724 3500 59780 3556
rect 60732 6130 60788 6132
rect 60732 6078 60734 6130
rect 60734 6078 60786 6130
rect 60786 6078 60788 6130
rect 60732 6076 60788 6078
rect 60956 5180 61012 5236
rect 60396 3388 60452 3444
rect 62076 6300 62132 6356
rect 61628 6188 61684 6244
rect 62076 5234 62132 5236
rect 62076 5182 62078 5234
rect 62078 5182 62130 5234
rect 62130 5182 62132 5234
rect 62076 5180 62132 5182
rect 61740 4172 61796 4228
rect 61292 3666 61348 3668
rect 61292 3614 61294 3666
rect 61294 3614 61346 3666
rect 61346 3614 61348 3666
rect 61292 3612 61348 3614
rect 61852 3500 61908 3556
rect 62748 57650 62804 57652
rect 62748 57598 62750 57650
rect 62750 57598 62802 57650
rect 62802 57598 62804 57650
rect 62748 57596 62804 57598
rect 62636 57426 62692 57428
rect 62636 57374 62638 57426
rect 62638 57374 62690 57426
rect 62690 57374 62692 57426
rect 62636 57372 62692 57374
rect 62972 61404 63028 61460
rect 63308 62748 63364 62804
rect 63868 62354 63924 62356
rect 63868 62302 63870 62354
rect 63870 62302 63922 62354
rect 63922 62302 63924 62354
rect 63868 62300 63924 62302
rect 65100 64092 65156 64148
rect 65100 63868 65156 63924
rect 65324 64482 65380 64484
rect 65324 64430 65326 64482
rect 65326 64430 65378 64482
rect 65378 64430 65380 64482
rect 65324 64428 65380 64430
rect 65548 64092 65604 64148
rect 65548 63922 65604 63924
rect 65548 63870 65550 63922
rect 65550 63870 65602 63922
rect 65602 63870 65604 63922
rect 65548 63868 65604 63870
rect 65324 62412 65380 62468
rect 63644 62076 63700 62132
rect 63308 61458 63364 61460
rect 63308 61406 63310 61458
rect 63310 61406 63362 61458
rect 63362 61406 63364 61458
rect 63308 61404 63364 61406
rect 63196 60844 63252 60900
rect 63420 61068 63476 61124
rect 63084 60786 63140 60788
rect 63084 60734 63086 60786
rect 63086 60734 63138 60786
rect 63138 60734 63140 60786
rect 63084 60732 63140 60734
rect 63196 57650 63252 57652
rect 63196 57598 63198 57650
rect 63198 57598 63250 57650
rect 63250 57598 63252 57650
rect 63196 57596 63252 57598
rect 63420 6636 63476 6692
rect 63532 60844 63588 60900
rect 63644 60732 63700 60788
rect 63532 6300 63588 6356
rect 62860 6188 62916 6244
rect 64316 62242 64372 62244
rect 64316 62190 64318 62242
rect 64318 62190 64370 62242
rect 64370 62190 64372 62242
rect 64316 62188 64372 62190
rect 64204 61570 64260 61572
rect 64204 61518 64206 61570
rect 64206 61518 64258 61570
rect 64258 61518 64260 61570
rect 64204 61516 64260 61518
rect 64540 60562 64596 60564
rect 64540 60510 64542 60562
rect 64542 60510 64594 60562
rect 64594 60510 64596 60562
rect 64540 60508 64596 60510
rect 63756 6076 63812 6132
rect 62412 4284 62468 4340
rect 63084 4226 63140 4228
rect 63084 4174 63086 4226
rect 63086 4174 63138 4226
rect 63138 4174 63140 4226
rect 63084 4172 63140 4174
rect 62524 3612 62580 3668
rect 63756 5068 63812 5124
rect 64204 6188 64260 6244
rect 65772 64540 65828 64596
rect 65884 64146 65940 64148
rect 65884 64094 65886 64146
rect 65886 64094 65938 64146
rect 65938 64094 65940 64146
rect 65884 64092 65940 64094
rect 66556 65660 66612 65716
rect 66332 64594 66388 64596
rect 66332 64542 66334 64594
rect 66334 64542 66386 64594
rect 66386 64542 66388 64594
rect 66332 64540 66388 64542
rect 66444 64316 66500 64372
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 66108 62076 66164 62132
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 65436 6188 65492 6244
rect 65772 6300 65828 6356
rect 63868 4338 63924 4340
rect 63868 4286 63870 4338
rect 63870 4286 63922 4338
rect 63922 4286 63924 4338
rect 63868 4284 63924 4286
rect 63756 4172 63812 4228
rect 63308 3442 63364 3444
rect 63308 3390 63310 3442
rect 63310 3390 63362 3442
rect 63362 3390 63364 3442
rect 63308 3388 63364 3390
rect 65324 6130 65380 6132
rect 65324 6078 65326 6130
rect 65326 6078 65378 6130
rect 65378 6078 65380 6130
rect 65324 6076 65380 6078
rect 64316 5122 64372 5124
rect 64316 5070 64318 5122
rect 64318 5070 64370 5122
rect 64370 5070 64372 5122
rect 64316 5068 64372 5070
rect 64540 4338 64596 4340
rect 64540 4286 64542 4338
rect 64542 4286 64594 4338
rect 64594 4286 64596 4338
rect 64540 4284 64596 4286
rect 64428 3500 64484 3556
rect 66108 6636 66164 6692
rect 67004 65772 67060 65828
rect 67788 66050 67844 66052
rect 67788 65998 67790 66050
rect 67790 65998 67842 66050
rect 67842 65998 67844 66050
rect 67788 65996 67844 65998
rect 68572 68012 68628 68068
rect 68236 67058 68292 67060
rect 68236 67006 68238 67058
rect 68238 67006 68290 67058
rect 68290 67006 68292 67058
rect 68236 67004 68292 67006
rect 68348 66668 68404 66724
rect 68124 66444 68180 66500
rect 69580 71932 69636 71988
rect 69468 70194 69524 70196
rect 69468 70142 69470 70194
rect 69470 70142 69522 70194
rect 69522 70142 69524 70194
rect 69468 70140 69524 70142
rect 69356 70028 69412 70084
rect 69692 69298 69748 69300
rect 69692 69246 69694 69298
rect 69694 69246 69746 69298
rect 69746 69246 69748 69298
rect 69692 69244 69748 69246
rect 69468 67954 69524 67956
rect 69468 67902 69470 67954
rect 69470 67902 69522 67954
rect 69522 67902 69524 67954
rect 69468 67900 69524 67902
rect 72156 72546 72212 72548
rect 72156 72494 72158 72546
rect 72158 72494 72210 72546
rect 72210 72494 72212 72546
rect 72156 72492 72212 72494
rect 72492 72492 72548 72548
rect 73052 72546 73108 72548
rect 73052 72494 73054 72546
rect 73054 72494 73106 72546
rect 73106 72494 73108 72546
rect 73052 72492 73108 72494
rect 75068 74898 75124 74900
rect 75068 74846 75070 74898
rect 75070 74846 75122 74898
rect 75122 74846 75124 74898
rect 75068 74844 75124 74846
rect 76076 74508 76132 74564
rect 74060 73948 74116 74004
rect 73836 73442 73892 73444
rect 73836 73390 73838 73442
rect 73838 73390 73890 73442
rect 73890 73390 73892 73442
rect 73836 73388 73892 73390
rect 73612 72604 73668 72660
rect 73724 72492 73780 72548
rect 72492 72268 72548 72324
rect 76860 73948 76916 74004
rect 77308 74002 77364 74004
rect 77308 73950 77310 74002
rect 77310 73950 77362 74002
rect 77362 73950 77364 74002
rect 77308 73948 77364 73950
rect 75068 73330 75124 73332
rect 75068 73278 75070 73330
rect 75070 73278 75122 73330
rect 75122 73278 75124 73330
rect 75068 73276 75124 73278
rect 74172 72658 74228 72660
rect 74172 72606 74174 72658
rect 74174 72606 74226 72658
rect 74226 72606 74228 72658
rect 74172 72604 74228 72606
rect 74620 72658 74676 72660
rect 74620 72606 74622 72658
rect 74622 72606 74674 72658
rect 74674 72606 74676 72658
rect 74620 72604 74676 72606
rect 75068 72546 75124 72548
rect 75068 72494 75070 72546
rect 75070 72494 75122 72546
rect 75122 72494 75124 72546
rect 75068 72492 75124 72494
rect 76076 72492 76132 72548
rect 73836 72380 73892 72436
rect 74060 72380 74116 72436
rect 73388 71986 73444 71988
rect 73388 71934 73390 71986
rect 73390 71934 73442 71986
rect 73442 71934 73444 71986
rect 73388 71932 73444 71934
rect 71148 71874 71204 71876
rect 71148 71822 71150 71874
rect 71150 71822 71202 71874
rect 71202 71822 71204 71874
rect 71148 71820 71204 71822
rect 70700 71762 70756 71764
rect 70700 71710 70702 71762
rect 70702 71710 70754 71762
rect 70754 71710 70756 71762
rect 70700 71708 70756 71710
rect 71484 71762 71540 71764
rect 71484 71710 71486 71762
rect 71486 71710 71538 71762
rect 71538 71710 71540 71762
rect 71484 71708 71540 71710
rect 72268 71762 72324 71764
rect 72268 71710 72270 71762
rect 72270 71710 72322 71762
rect 72322 71710 72324 71762
rect 72268 71708 72324 71710
rect 72828 71708 72884 71764
rect 70588 71596 70644 71652
rect 70140 70754 70196 70756
rect 70140 70702 70142 70754
rect 70142 70702 70194 70754
rect 70194 70702 70196 70754
rect 70140 70700 70196 70702
rect 70924 70700 70980 70756
rect 71932 70866 71988 70868
rect 71932 70814 71934 70866
rect 71934 70814 71986 70866
rect 71986 70814 71988 70866
rect 71932 70812 71988 70814
rect 71820 70700 71876 70756
rect 71260 70588 71316 70644
rect 69916 70306 69972 70308
rect 69916 70254 69918 70306
rect 69918 70254 69970 70306
rect 69970 70254 69972 70306
rect 69916 70252 69972 70254
rect 70252 70194 70308 70196
rect 70252 70142 70254 70194
rect 70254 70142 70306 70194
rect 70306 70142 70308 70194
rect 70252 70140 70308 70142
rect 70924 70194 70980 70196
rect 70924 70142 70926 70194
rect 70926 70142 70978 70194
rect 70978 70142 70980 70194
rect 70924 70140 70980 70142
rect 70252 69298 70308 69300
rect 70252 69246 70254 69298
rect 70254 69246 70306 69298
rect 70306 69246 70308 69298
rect 70252 69244 70308 69246
rect 70588 69298 70644 69300
rect 70588 69246 70590 69298
rect 70590 69246 70642 69298
rect 70642 69246 70644 69298
rect 70588 69244 70644 69246
rect 70028 68012 70084 68068
rect 68796 66444 68852 66500
rect 68684 66332 68740 66388
rect 68572 65996 68628 66052
rect 68348 65660 68404 65716
rect 66668 64316 66724 64372
rect 66332 6636 66388 6692
rect 66668 63980 66724 64036
rect 67788 64482 67844 64484
rect 67788 64430 67790 64482
rect 67790 64430 67842 64482
rect 67842 64430 67844 64482
rect 67788 64428 67844 64430
rect 68012 64428 68068 64484
rect 67676 64146 67732 64148
rect 67676 64094 67678 64146
rect 67678 64094 67730 64146
rect 67730 64094 67732 64146
rect 67676 64092 67732 64094
rect 67452 63980 67508 64036
rect 67004 63868 67060 63924
rect 67340 63922 67396 63924
rect 67340 63870 67342 63922
rect 67342 63870 67394 63922
rect 67394 63870 67396 63922
rect 67340 63868 67396 63870
rect 66332 6188 66388 6244
rect 65884 5852 65940 5908
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 66668 62076 66724 62132
rect 66668 60114 66724 60116
rect 66668 60062 66670 60114
rect 66670 60062 66722 60114
rect 66722 60062 66724 60114
rect 66668 60060 66724 60062
rect 67228 60114 67284 60116
rect 67228 60062 67230 60114
rect 67230 60062 67282 60114
rect 67282 60062 67284 60114
rect 67228 60060 67284 60062
rect 66556 60002 66612 60004
rect 66556 59950 66558 60002
rect 66558 59950 66610 60002
rect 66610 59950 66612 60002
rect 66556 59948 66612 59950
rect 68236 62524 68292 62580
rect 68460 65436 68516 65492
rect 68460 64540 68516 64596
rect 68460 64092 68516 64148
rect 68236 62242 68292 62244
rect 68236 62190 68238 62242
rect 68238 62190 68290 62242
rect 68290 62190 68292 62242
rect 68236 62188 68292 62190
rect 67676 6636 67732 6692
rect 66444 6076 66500 6132
rect 66780 6188 66836 6244
rect 67228 6076 67284 6132
rect 66108 4226 66164 4228
rect 66108 4174 66110 4226
rect 66110 4174 66162 4226
rect 66162 4174 66164 4226
rect 66108 4172 66164 4174
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 65212 3666 65268 3668
rect 65212 3614 65214 3666
rect 65214 3614 65266 3666
rect 65266 3614 65268 3666
rect 65212 3612 65268 3614
rect 65772 3500 65828 3556
rect 67116 5180 67172 5236
rect 67004 3666 67060 3668
rect 67004 3614 67006 3666
rect 67006 3614 67058 3666
rect 67058 3614 67060 3666
rect 67004 3612 67060 3614
rect 66444 3388 66500 3444
rect 68012 49868 68068 49924
rect 68012 49138 68068 49140
rect 68012 49086 68014 49138
rect 68014 49086 68066 49138
rect 68066 49086 68068 49138
rect 68012 49084 68068 49086
rect 68124 48802 68180 48804
rect 68124 48750 68126 48802
rect 68126 48750 68178 48802
rect 68178 48750 68180 48802
rect 68124 48748 68180 48750
rect 68796 65436 68852 65492
rect 68684 64428 68740 64484
rect 69356 66946 69412 66948
rect 69356 66894 69358 66946
rect 69358 66894 69410 66946
rect 69410 66894 69412 66946
rect 69356 66892 69412 66894
rect 69244 66332 69300 66388
rect 69356 64594 69412 64596
rect 69356 64542 69358 64594
rect 69358 64542 69410 64594
rect 69410 64542 69412 64594
rect 69356 64540 69412 64542
rect 68796 62578 68852 62580
rect 68796 62526 68798 62578
rect 68798 62526 68850 62578
rect 68850 62526 68852 62578
rect 68796 62524 68852 62526
rect 68684 50706 68740 50708
rect 68684 50654 68686 50706
rect 68686 50654 68738 50706
rect 68738 50654 68740 50706
rect 68684 50652 68740 50654
rect 68572 49138 68628 49140
rect 68572 49086 68574 49138
rect 68574 49086 68626 49138
rect 68626 49086 68628 49138
rect 68572 49084 68628 49086
rect 68908 49810 68964 49812
rect 68908 49758 68910 49810
rect 68910 49758 68962 49810
rect 68962 49758 68964 49810
rect 68908 49756 68964 49758
rect 70028 50764 70084 50820
rect 69356 50706 69412 50708
rect 69356 50654 69358 50706
rect 69358 50654 69410 50706
rect 69410 50654 69412 50706
rect 69356 50652 69412 50654
rect 69244 49756 69300 49812
rect 69580 49810 69636 49812
rect 69580 49758 69582 49810
rect 69582 49758 69634 49810
rect 69634 49758 69636 49810
rect 69580 49756 69636 49758
rect 69916 49756 69972 49812
rect 70252 49980 70308 50036
rect 69580 49532 69636 49588
rect 68796 48412 68852 48468
rect 70028 49698 70084 49700
rect 70028 49646 70030 49698
rect 70030 49646 70082 49698
rect 70082 49646 70084 49698
rect 70028 49644 70084 49646
rect 69804 48802 69860 48804
rect 69804 48750 69806 48802
rect 69806 48750 69858 48802
rect 69858 48750 69860 48802
rect 69804 48748 69860 48750
rect 69356 48466 69412 48468
rect 69356 48414 69358 48466
rect 69358 48414 69410 48466
rect 69410 48414 69412 48466
rect 69356 48412 69412 48414
rect 69468 48300 69524 48356
rect 69916 48300 69972 48356
rect 68572 6188 68628 6244
rect 69132 6188 69188 6244
rect 68460 6076 68516 6132
rect 69020 6130 69076 6132
rect 69020 6078 69022 6130
rect 69022 6078 69074 6130
rect 69074 6078 69076 6130
rect 69020 6076 69076 6078
rect 68124 5852 68180 5908
rect 68012 5234 68068 5236
rect 68012 5182 68014 5234
rect 68014 5182 68066 5234
rect 68066 5182 68068 5234
rect 68012 5180 68068 5182
rect 67900 4396 67956 4452
rect 67788 4172 67844 4228
rect 67900 3500 67956 3556
rect 69468 6188 69524 6244
rect 69244 5740 69300 5796
rect 69356 6076 69412 6132
rect 69692 5404 69748 5460
rect 68572 3500 68628 3556
rect 69356 3442 69412 3444
rect 69356 3390 69358 3442
rect 69358 3390 69410 3442
rect 69410 3390 69412 3442
rect 69356 3388 69412 3390
rect 70700 50764 70756 50820
rect 70700 49698 70756 49700
rect 70700 49646 70702 49698
rect 70702 49646 70754 49698
rect 70754 49646 70756 49698
rect 70700 49644 70756 49646
rect 71708 70194 71764 70196
rect 71708 70142 71710 70194
rect 71710 70142 71762 70194
rect 71762 70142 71764 70194
rect 71708 70140 71764 70142
rect 71148 69186 71204 69188
rect 71148 69134 71150 69186
rect 71150 69134 71202 69186
rect 71202 69134 71204 69186
rect 71148 69132 71204 69134
rect 72380 70754 72436 70756
rect 72380 70702 72382 70754
rect 72382 70702 72434 70754
rect 72434 70702 72436 70754
rect 72380 70700 72436 70702
rect 73948 71932 74004 71988
rect 76860 72268 76916 72324
rect 76076 71148 76132 71204
rect 75068 70812 75124 70868
rect 76860 70588 76916 70644
rect 76860 69244 76916 69300
rect 76524 69132 76580 69188
rect 77308 69186 77364 69188
rect 77308 69134 77310 69186
rect 77310 69134 77362 69186
rect 77362 69134 77364 69186
rect 77308 69132 77364 69134
rect 76188 68684 76244 68740
rect 75964 68626 76020 68628
rect 75964 68574 75966 68626
rect 75966 68574 76018 68626
rect 76018 68574 76020 68626
rect 75964 68572 76020 68574
rect 76412 68514 76468 68516
rect 76412 68462 76414 68514
rect 76414 68462 76466 68514
rect 76466 68462 76468 68514
rect 76412 68460 76468 68462
rect 77196 68460 77252 68516
rect 76860 67900 76916 67956
rect 77308 67842 77364 67844
rect 77308 67790 77310 67842
rect 77310 67790 77362 67842
rect 77362 67790 77364 67842
rect 77308 67788 77364 67790
rect 70364 4508 70420 4564
rect 69804 4284 69860 4340
rect 69692 4226 69748 4228
rect 69692 4174 69694 4226
rect 69694 4174 69746 4226
rect 69746 4174 69748 4226
rect 69692 4172 69748 4174
rect 70588 3554 70644 3556
rect 70588 3502 70590 3554
rect 70590 3502 70642 3554
rect 70642 3502 70644 3554
rect 70588 3500 70644 3502
rect 70476 3388 70532 3444
rect 71148 4562 71204 4564
rect 71148 4510 71150 4562
rect 71150 4510 71202 4562
rect 71202 4510 71204 4562
rect 71148 4508 71204 4510
rect 71260 4396 71316 4452
rect 70812 4338 70868 4340
rect 70812 4286 70814 4338
rect 70814 4286 70866 4338
rect 70866 4286 70868 4338
rect 70812 4284 70868 4286
rect 71148 4284 71204 4340
rect 70700 3276 70756 3332
rect 71260 3612 71316 3668
rect 72044 4338 72100 4340
rect 72044 4286 72046 4338
rect 72046 4286 72098 4338
rect 72098 4286 72100 4338
rect 72044 4284 72100 4286
rect 72492 4338 72548 4340
rect 72492 4286 72494 4338
rect 72494 4286 72546 4338
rect 72546 4286 72548 4338
rect 72492 4284 72548 4286
rect 73500 4508 73556 4564
rect 74620 47180 74676 47236
rect 74620 45724 74676 45780
rect 74732 45666 74788 45668
rect 74732 45614 74734 45666
rect 74734 45614 74786 45666
rect 74786 45614 74788 45666
rect 74732 45612 74788 45614
rect 74620 44156 74676 44212
rect 74620 41020 74676 41076
rect 74620 39452 74676 39508
rect 74732 39004 74788 39060
rect 74620 37772 74676 37828
rect 74620 36204 74676 36260
rect 74620 34748 74676 34804
rect 74732 34300 74788 34356
rect 74620 33068 74676 33124
rect 74620 31500 74676 31556
rect 74620 30044 74676 30100
rect 74732 29596 74788 29652
rect 74620 28364 74676 28420
rect 74620 26796 74676 26852
rect 74620 25228 74676 25284
rect 74732 25116 74788 25172
rect 74620 23772 74676 23828
rect 74508 23660 74564 23716
rect 74620 22092 74676 22148
rect 74508 20524 74564 20580
rect 74508 20076 74564 20132
rect 74620 19068 74676 19124
rect 74508 18956 74564 19012
rect 74620 17836 74676 17892
rect 74508 17724 74564 17780
rect 74732 16044 74788 16100
rect 74732 15372 74788 15428
rect 74620 15202 74676 15204
rect 74620 15150 74622 15202
rect 74622 15150 74674 15202
rect 74674 15150 74676 15202
rect 74620 15148 74676 15150
rect 75068 15148 75124 15204
rect 74620 13746 74676 13748
rect 74620 13694 74622 13746
rect 74622 13694 74674 13746
rect 74674 13694 74676 13746
rect 74620 13692 74676 13694
rect 75068 13746 75124 13748
rect 75068 13694 75070 13746
rect 75070 13694 75122 13746
rect 75122 13694 75124 13746
rect 75068 13692 75124 13694
rect 74620 11228 74676 11284
rect 74732 10780 74788 10836
rect 74620 9548 74676 9604
rect 74620 7980 74676 8036
rect 74620 6524 74676 6580
rect 74732 6636 74788 6692
rect 74732 5964 74788 6020
rect 74396 5404 74452 5460
rect 73164 3666 73220 3668
rect 73164 3614 73166 3666
rect 73166 3614 73218 3666
rect 73218 3614 73220 3666
rect 73164 3612 73220 3614
rect 72716 3442 72772 3444
rect 72716 3390 72718 3442
rect 72718 3390 72770 3442
rect 72770 3390 72772 3442
rect 72716 3388 72772 3390
rect 72380 3330 72436 3332
rect 72380 3278 72382 3330
rect 72382 3278 72434 3330
rect 72434 3278 72436 3330
rect 72380 3276 72436 3278
rect 73500 4284 73556 4340
rect 74284 4562 74340 4564
rect 74284 4510 74286 4562
rect 74286 4510 74338 4562
rect 74338 4510 74340 4562
rect 74284 4508 74340 4510
rect 74060 4284 74116 4340
rect 74620 4844 74676 4900
rect 74508 4338 74564 4340
rect 74508 4286 74510 4338
rect 74510 4286 74562 4338
rect 74562 4286 74564 4338
rect 74508 4284 74564 4286
rect 77308 67058 77364 67060
rect 77308 67006 77310 67058
rect 77310 67006 77362 67058
rect 77362 67006 77364 67058
rect 77308 67004 77364 67006
rect 77308 66050 77364 66052
rect 77308 65998 77310 66050
rect 77310 65998 77362 66050
rect 77362 65998 77364 66050
rect 77308 65996 77364 65998
rect 77308 65378 77364 65380
rect 77308 65326 77310 65378
rect 77310 65326 77362 65378
rect 77362 65326 77364 65378
rect 77308 65324 77364 65326
rect 76636 64594 76692 64596
rect 76636 64542 76638 64594
rect 76638 64542 76690 64594
rect 76690 64542 76692 64594
rect 76636 64540 76692 64542
rect 76860 64204 76916 64260
rect 77308 64204 77364 64260
rect 77420 63980 77476 64036
rect 76412 63922 76468 63924
rect 76412 63870 76414 63922
rect 76414 63870 76466 63922
rect 76466 63870 76468 63922
rect 76412 63868 76468 63870
rect 77196 63922 77252 63924
rect 77196 63870 77198 63922
rect 77198 63870 77250 63922
rect 77250 63870 77252 63922
rect 77196 63868 77252 63870
rect 77308 63026 77364 63028
rect 77308 62974 77310 63026
rect 77310 62974 77362 63026
rect 77362 62974 77364 63026
rect 77308 62972 77364 62974
rect 77308 62242 77364 62244
rect 77308 62190 77310 62242
rect 77310 62190 77362 62242
rect 77362 62190 77364 62242
rect 77308 62188 77364 62190
rect 77420 61516 77476 61572
rect 77308 61458 77364 61460
rect 77308 61406 77310 61458
rect 77310 61406 77362 61458
rect 77362 61406 77364 61458
rect 77308 61404 77364 61406
rect 77308 60674 77364 60676
rect 77308 60622 77310 60674
rect 77310 60622 77362 60674
rect 77362 60622 77364 60674
rect 77308 60620 77364 60622
rect 76636 59778 76692 59780
rect 76636 59726 76638 59778
rect 76638 59726 76690 59778
rect 76690 59726 76692 59778
rect 76636 59724 76692 59726
rect 76412 59106 76468 59108
rect 76412 59054 76414 59106
rect 76414 59054 76466 59106
rect 76466 59054 76468 59106
rect 76412 59052 76468 59054
rect 77308 59164 77364 59220
rect 77196 59052 77252 59108
rect 76860 58380 76916 58436
rect 77308 58322 77364 58324
rect 77308 58270 77310 58322
rect 77310 58270 77362 58322
rect 77362 58270 77364 58322
rect 77308 58268 77364 58270
rect 77308 57538 77364 57540
rect 77308 57486 77310 57538
rect 77310 57486 77362 57538
rect 77362 57486 77364 57538
rect 77308 57484 77364 57486
rect 77308 56642 77364 56644
rect 77308 56590 77310 56642
rect 77310 56590 77362 56642
rect 77362 56590 77364 56642
rect 77308 56588 77364 56590
rect 77308 55970 77364 55972
rect 77308 55918 77310 55970
rect 77310 55918 77362 55970
rect 77362 55918 77364 55970
rect 77308 55916 77364 55918
rect 78092 74002 78148 74004
rect 78092 73950 78094 74002
rect 78094 73950 78146 74002
rect 78146 73950 78148 74002
rect 78092 73948 78148 73950
rect 77868 73388 77924 73444
rect 77868 71820 77924 71876
rect 77868 70588 77924 70644
rect 77868 69804 77924 69860
rect 77980 68626 78036 68628
rect 77980 68574 77982 68626
rect 77982 68574 78034 68626
rect 78034 68574 78036 68626
rect 77980 68572 78036 68574
rect 77868 68012 77924 68068
rect 77980 67842 78036 67844
rect 77980 67790 77982 67842
rect 77982 67790 78034 67842
rect 78034 67790 78036 67842
rect 77980 67788 78036 67790
rect 77644 66892 77700 66948
rect 77868 67116 77924 67172
rect 78204 67788 78260 67844
rect 78092 67340 78148 67396
rect 78092 67058 78148 67060
rect 78092 67006 78094 67058
rect 78094 67006 78146 67058
rect 78146 67006 78148 67058
rect 78092 67004 78148 67006
rect 77980 66444 78036 66500
rect 77756 66220 77812 66276
rect 77756 65772 77812 65828
rect 78092 65996 78148 66052
rect 77756 64652 77812 64708
rect 77980 65324 78036 65380
rect 78204 65772 78260 65828
rect 78092 65100 78148 65156
rect 77980 64428 78036 64484
rect 78092 64594 78148 64596
rect 78092 64542 78094 64594
rect 78094 64542 78146 64594
rect 78146 64542 78148 64594
rect 78092 64540 78148 64542
rect 77980 64204 78036 64260
rect 77756 64034 77812 64036
rect 77756 63982 77758 64034
rect 77758 63982 77810 64034
rect 77810 63982 77812 64034
rect 77756 63980 77812 63982
rect 77644 62524 77700 62580
rect 77756 62466 77812 62468
rect 77756 62414 77758 62466
rect 77758 62414 77810 62466
rect 77810 62414 77812 62466
rect 77756 62412 77812 62414
rect 78092 63196 78148 63252
rect 77980 62524 78036 62580
rect 78092 63026 78148 63028
rect 78092 62974 78094 63026
rect 78094 62974 78146 63026
rect 78146 62974 78148 63026
rect 78092 62972 78148 62974
rect 77868 61292 77924 61348
rect 77980 62188 78036 62244
rect 78092 61740 78148 61796
rect 78092 61458 78148 61460
rect 78092 61406 78094 61458
rect 78094 61406 78146 61458
rect 78146 61406 78148 61458
rect 78092 61404 78148 61406
rect 77980 61068 78036 61124
rect 77756 60172 77812 60228
rect 78092 60620 78148 60676
rect 77644 60060 77700 60116
rect 78204 60508 78260 60564
rect 78092 59836 78148 59892
rect 77980 59724 78036 59780
rect 77644 58492 77700 58548
rect 77756 58210 77812 58212
rect 77756 58158 77758 58210
rect 77758 58158 77810 58210
rect 77810 58158 77812 58210
rect 77756 58156 77812 58158
rect 77980 58828 78036 58884
rect 78092 59218 78148 59220
rect 78092 59166 78094 59218
rect 78094 59166 78146 59218
rect 78146 59166 78148 59218
rect 78092 59164 78148 59166
rect 77868 57596 77924 57652
rect 77980 58268 78036 58324
rect 78092 57820 78148 57876
rect 77980 57260 78036 57316
rect 78092 57484 78148 57540
rect 77756 56194 77812 56196
rect 77756 56142 77758 56194
rect 77758 56142 77810 56194
rect 77810 56142 77812 56194
rect 77756 56140 77812 56142
rect 77644 56028 77700 56084
rect 76636 55074 76692 55076
rect 76636 55022 76638 55074
rect 76638 55022 76690 55074
rect 76690 55022 76692 55074
rect 76636 55020 76692 55022
rect 76860 54738 76916 54740
rect 76860 54686 76862 54738
rect 76862 54686 76914 54738
rect 76914 54686 76916 54738
rect 76860 54684 76916 54686
rect 76412 54402 76468 54404
rect 76412 54350 76414 54402
rect 76414 54350 76466 54402
rect 76466 54350 76468 54402
rect 76412 54348 76468 54350
rect 77308 54460 77364 54516
rect 77196 54348 77252 54404
rect 77308 53506 77364 53508
rect 77308 53454 77310 53506
rect 77310 53454 77362 53506
rect 77362 53454 77364 53506
rect 77308 53452 77364 53454
rect 77308 52834 77364 52836
rect 77308 52782 77310 52834
rect 77310 52782 77362 52834
rect 77362 52782 77364 52834
rect 77308 52780 77364 52782
rect 77308 51938 77364 51940
rect 77308 51886 77310 51938
rect 77310 51886 77362 51938
rect 77362 51886 77364 51938
rect 77308 51884 77364 51886
rect 77308 51266 77364 51268
rect 77308 51214 77310 51266
rect 77310 51214 77362 51266
rect 77362 51214 77364 51266
rect 77308 51212 77364 51214
rect 77980 56588 78036 56644
rect 78092 56364 78148 56420
rect 77980 55692 78036 55748
rect 78092 55916 78148 55972
rect 78092 55468 78148 55524
rect 77868 54796 77924 54852
rect 77980 55020 78036 55076
rect 77756 54626 77812 54628
rect 77756 54574 77758 54626
rect 77758 54574 77810 54626
rect 77810 54574 77812 54626
rect 77756 54572 77812 54574
rect 78092 54514 78148 54516
rect 78092 54462 78094 54514
rect 78094 54462 78146 54514
rect 78146 54462 78148 54514
rect 78092 54460 78148 54462
rect 77980 53788 78036 53844
rect 77644 53676 77700 53732
rect 78092 53452 78148 53508
rect 77644 52220 77700 52276
rect 77756 52108 77812 52164
rect 77980 52780 78036 52836
rect 77420 50764 77476 50820
rect 77308 50706 77364 50708
rect 77308 50654 77310 50706
rect 77310 50654 77362 50706
rect 77362 50654 77364 50706
rect 77308 50652 77364 50654
rect 78204 53004 78260 53060
rect 78092 52332 78148 52388
rect 77980 51660 78036 51716
rect 78092 51884 78148 51940
rect 77756 51490 77812 51492
rect 77756 51438 77758 51490
rect 77758 51438 77810 51490
rect 77810 51438 77812 51490
rect 77756 51436 77812 51438
rect 77644 50540 77700 50596
rect 77980 51212 78036 51268
rect 78092 50988 78148 51044
rect 77980 50428 78036 50484
rect 78092 50652 78148 50708
rect 77756 50370 77812 50372
rect 77756 50318 77758 50370
rect 77758 50318 77810 50370
rect 77810 50318 77812 50370
rect 77756 50316 77812 50318
rect 77308 49698 77364 49700
rect 77308 49646 77310 49698
rect 77310 49646 77362 49698
rect 77362 49646 77364 49698
rect 77308 49644 77364 49646
rect 77756 48972 77812 49028
rect 78092 49756 78148 49812
rect 77980 49644 78036 49700
rect 77980 48972 78036 49028
rect 77308 48802 77364 48804
rect 77308 48750 77310 48802
rect 77310 48750 77362 48802
rect 77362 48750 77364 48802
rect 77308 48748 77364 48750
rect 77756 48412 77812 48468
rect 78092 48748 78148 48804
rect 78092 48300 78148 48356
rect 76076 47628 76132 47684
rect 77868 47068 77924 47124
rect 76972 46732 77028 46788
rect 76076 46284 76132 46340
rect 75292 45612 75348 45668
rect 76188 45612 76244 45668
rect 76076 44268 76132 44324
rect 77756 44940 77812 44996
rect 77084 44044 77140 44100
rect 76524 43708 76580 43764
rect 77868 43708 77924 43764
rect 77868 42924 77924 42980
rect 76412 42476 76468 42532
rect 76076 41580 76132 41636
rect 77756 41970 77812 41972
rect 77756 41918 77758 41970
rect 77758 41918 77810 41970
rect 77810 41918 77812 41970
rect 77756 41916 77812 41918
rect 76636 40962 76692 40964
rect 76636 40910 76638 40962
rect 76638 40910 76690 40962
rect 76690 40910 76692 40962
rect 76636 40908 76692 40910
rect 77756 40908 77812 40964
rect 76860 40460 76916 40516
rect 75964 40402 76020 40404
rect 75964 40350 75966 40402
rect 75966 40350 76018 40402
rect 76018 40350 76020 40402
rect 75964 40348 76020 40350
rect 77196 40460 77252 40516
rect 77756 39564 77812 39620
rect 75292 39004 75348 39060
rect 76188 38892 76244 38948
rect 76860 39340 76916 39396
rect 76076 38220 76132 38276
rect 77756 37548 77812 37604
rect 76636 37324 76692 37380
rect 76076 36988 76132 37044
rect 76860 37324 76916 37380
rect 77756 36204 77812 36260
rect 76860 35756 76916 35812
rect 77196 35756 77252 35812
rect 76076 35586 76132 35588
rect 76076 35534 76078 35586
rect 76078 35534 76130 35586
rect 76130 35534 76132 35586
rect 76076 35532 76132 35534
rect 77756 34860 77812 34916
rect 75292 34300 75348 34356
rect 76188 34188 76244 34244
rect 76860 34636 76916 34692
rect 76076 33628 76132 33684
rect 77756 32844 77812 32900
rect 76636 32620 76692 32676
rect 76076 32172 76132 32228
rect 77756 31500 77812 31556
rect 76860 31052 76916 31108
rect 77196 31052 77252 31108
rect 76076 30882 76132 30884
rect 76076 30830 76078 30882
rect 76078 30830 76130 30882
rect 76130 30830 76132 30882
rect 76076 30828 76132 30830
rect 77756 30156 77812 30212
rect 75292 29596 75348 29652
rect 76188 29484 76244 29540
rect 76860 29932 76916 29988
rect 76076 28812 76132 28868
rect 77756 28140 77812 28196
rect 76636 27916 76692 27972
rect 76076 27468 76132 27524
rect 76860 27916 76916 27972
rect 77756 26796 77812 26852
rect 76860 26348 76916 26404
rect 77196 26348 77252 26404
rect 76076 26178 76132 26180
rect 76076 26126 76078 26178
rect 76078 26126 76130 26178
rect 76130 26126 76132 26178
rect 76076 26124 76132 26126
rect 77756 25452 77812 25508
rect 75292 25116 75348 25172
rect 76188 24780 76244 24836
rect 76636 24668 76692 24724
rect 76076 24108 76132 24164
rect 76860 24722 76916 24724
rect 76860 24670 76862 24722
rect 76862 24670 76914 24722
rect 76914 24670 76916 24722
rect 76860 24668 76916 24670
rect 77756 23436 77812 23492
rect 76636 23212 76692 23268
rect 76076 22764 76132 22820
rect 76860 23212 76916 23268
rect 77756 22092 77812 22148
rect 76860 21644 76916 21700
rect 77196 21644 77252 21700
rect 76076 21474 76132 21476
rect 76076 21422 76078 21474
rect 76078 21422 76130 21474
rect 76130 21422 76132 21474
rect 76076 21420 76132 21422
rect 76188 20188 76244 20244
rect 75292 20076 75348 20132
rect 77756 20130 77812 20132
rect 77756 20078 77758 20130
rect 77758 20078 77810 20130
rect 77810 20078 77812 20130
rect 77756 20076 77812 20078
rect 76076 19404 76132 19460
rect 76636 19852 76692 19908
rect 76860 19852 76916 19908
rect 76076 18060 76132 18116
rect 77756 18450 77812 18452
rect 77756 18398 77758 18450
rect 77758 18398 77810 18450
rect 77810 18398 77812 18450
rect 77756 18396 77812 18398
rect 76636 17666 76692 17668
rect 76636 17614 76638 17666
rect 76638 17614 76690 17666
rect 76690 17614 76692 17666
rect 76636 17612 76692 17614
rect 77756 17388 77812 17444
rect 76860 16940 76916 16996
rect 75964 16882 76020 16884
rect 75964 16830 75966 16882
rect 75966 16830 76018 16882
rect 76018 16830 76020 16882
rect 75964 16828 76020 16830
rect 77196 16940 77252 16996
rect 75292 16098 75348 16100
rect 75292 16046 75294 16098
rect 75294 16046 75346 16098
rect 75346 16046 75348 16098
rect 75292 16044 75348 16046
rect 77756 16044 77812 16100
rect 76188 15372 76244 15428
rect 76860 15820 76916 15876
rect 76076 14700 76132 14756
rect 77756 14028 77812 14084
rect 76636 13804 76692 13860
rect 76076 13468 76132 13524
rect 76860 13804 76916 13860
rect 77756 12684 77812 12740
rect 76860 12236 76916 12292
rect 77196 12236 77252 12292
rect 76076 12066 76132 12068
rect 76076 12014 76078 12066
rect 76078 12014 76130 12066
rect 76130 12014 76132 12066
rect 76076 12012 76132 12014
rect 77756 11340 77812 11396
rect 75292 10780 75348 10836
rect 76188 10668 76244 10724
rect 76860 11116 76916 11172
rect 76076 10108 76132 10164
rect 77756 9324 77812 9380
rect 76636 9100 76692 9156
rect 76076 8652 76132 8708
rect 77756 7980 77812 8036
rect 76860 7532 76916 7588
rect 77196 7532 77252 7588
rect 76076 7362 76132 7364
rect 76076 7310 76078 7362
rect 76078 7310 76130 7362
rect 76130 7310 76132 7362
rect 76076 7308 76132 7310
rect 75292 6690 75348 6692
rect 75292 6638 75294 6690
rect 75294 6638 75346 6690
rect 75346 6638 75348 6690
rect 75292 6636 75348 6638
rect 77756 6636 77812 6692
rect 76188 5964 76244 6020
rect 76860 6412 76916 6468
rect 76076 5292 76132 5348
rect 73836 3388 73892 3444
rect 74956 3442 75012 3444
rect 74956 3390 74958 3442
rect 74958 3390 75010 3442
rect 75010 3390 75012 3442
rect 74956 3388 75012 3390
<< metal3 >>
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 73714 74844 73724 74900
rect 73780 74844 75068 74900
rect 75124 74844 75134 74900
rect 3042 74732 3052 74788
rect 3108 74732 4060 74788
rect 4116 74732 4844 74788
rect 4900 74732 4910 74788
rect 0 74564 800 74592
rect 79200 74564 80000 74592
rect 0 74508 2044 74564
rect 2100 74508 2110 74564
rect 76066 74508 76076 74564
rect 76132 74508 80000 74564
rect 0 74480 800 74508
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 79200 74480 80000 74508
rect 3042 74060 3052 74116
rect 3108 74060 4284 74116
rect 4340 74060 4350 74116
rect 74050 73948 74060 74004
rect 74116 73948 76860 74004
rect 76916 73948 76926 74004
rect 77298 73948 77308 74004
rect 77364 73948 78092 74004
rect 78148 73948 78158 74004
rect 0 73892 800 73920
rect 78092 73892 78148 73948
rect 79200 73892 80000 73920
rect 0 73836 3612 73892
rect 3668 73836 3678 73892
rect 78092 73836 80000 73892
rect 0 73808 800 73836
rect 79200 73808 80000 73836
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 69346 73388 69356 73444
rect 69412 73388 73836 73444
rect 73892 73388 73902 73444
rect 77858 73388 77868 73444
rect 77924 73388 77934 73444
rect 69122 73276 69132 73332
rect 69188 73276 70028 73332
rect 70084 73276 70094 73332
rect 73266 73276 73276 73332
rect 73332 73276 75068 73332
rect 75124 73276 75134 73332
rect 0 73220 800 73248
rect 77868 73220 77924 73388
rect 79200 73220 80000 73248
rect 0 73164 2156 73220
rect 2212 73164 2222 73220
rect 3042 73164 3052 73220
rect 3108 73164 3612 73220
rect 3668 73164 71820 73220
rect 71876 73164 71886 73220
rect 77868 73164 80000 73220
rect 0 73136 800 73164
rect 79200 73136 80000 73164
rect 4834 73052 4844 73108
rect 4900 73052 69244 73108
rect 69300 73052 69310 73108
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 69794 72604 69804 72660
rect 69860 72604 73612 72660
rect 73668 72604 74172 72660
rect 74228 72604 74620 72660
rect 74676 72604 74686 72660
rect 0 72548 800 72576
rect 79200 72548 80000 72576
rect 0 72492 2044 72548
rect 2100 72492 2110 72548
rect 72146 72492 72156 72548
rect 72212 72492 72492 72548
rect 72548 72492 73052 72548
rect 73108 72492 73724 72548
rect 73780 72492 75068 72548
rect 75124 72492 75134 72548
rect 76066 72492 76076 72548
rect 76132 72492 80000 72548
rect 0 72464 800 72492
rect 79200 72464 80000 72492
rect 4274 72380 4284 72436
rect 4340 72380 69468 72436
rect 69524 72380 69534 72436
rect 73826 72380 73836 72436
rect 73892 72380 74060 72436
rect 74116 72380 74126 72436
rect 72482 72268 72492 72324
rect 72548 72268 76860 72324
rect 76916 72268 76926 72324
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 69570 71932 69580 71988
rect 69636 71932 73388 71988
rect 73444 71932 73948 71988
rect 74004 71932 74014 71988
rect 0 71876 800 71904
rect 79200 71876 80000 71904
rect 0 71820 2156 71876
rect 2212 71820 2222 71876
rect 3490 71820 3500 71876
rect 3556 71820 71148 71876
rect 71204 71820 71214 71876
rect 77858 71820 77868 71876
rect 77924 71820 80000 71876
rect 0 71792 800 71820
rect 79200 71792 80000 71820
rect 70690 71708 70700 71764
rect 70756 71708 71484 71764
rect 71540 71708 72268 71764
rect 72324 71708 72828 71764
rect 72884 71708 72894 71764
rect 3042 71596 3052 71652
rect 3108 71596 3612 71652
rect 3668 71596 70588 71652
rect 70644 71596 70654 71652
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 0 71204 800 71232
rect 79200 71204 80000 71232
rect 0 71148 2044 71204
rect 2100 71148 2110 71204
rect 76066 71148 76076 71204
rect 76132 71148 80000 71204
rect 0 71120 800 71148
rect 79200 71120 80000 71148
rect 71922 70812 71932 70868
rect 71988 70812 75068 70868
rect 75124 70812 75134 70868
rect 70130 70700 70140 70756
rect 70196 70700 70924 70756
rect 70980 70700 71820 70756
rect 71876 70700 72380 70756
rect 72436 70700 72446 70756
rect 71250 70588 71260 70644
rect 71316 70588 76860 70644
rect 76916 70588 76926 70644
rect 77858 70588 77868 70644
rect 77924 70588 77934 70644
rect 0 70532 800 70560
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 77868 70532 77924 70588
rect 79200 70532 80000 70560
rect 0 70476 2156 70532
rect 2212 70476 2222 70532
rect 77868 70476 80000 70532
rect 0 70448 800 70476
rect 79200 70448 80000 70476
rect 3490 70252 3500 70308
rect 3556 70252 69916 70308
rect 69972 70252 69982 70308
rect 69458 70140 69468 70196
rect 69524 70140 70252 70196
rect 70308 70140 70924 70196
rect 70980 70140 71708 70196
rect 71764 70140 71774 70196
rect 3042 70028 3052 70084
rect 3108 70028 3612 70084
rect 3668 70028 69356 70084
rect 69412 70028 69422 70084
rect 0 69860 800 69888
rect 79200 69860 80000 69888
rect 0 69804 2044 69860
rect 2100 69804 2110 69860
rect 77858 69804 77868 69860
rect 77924 69804 80000 69860
rect 0 69776 800 69804
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 79200 69776 80000 69804
rect 1810 69244 1820 69300
rect 1876 69244 3948 69300
rect 4004 69244 4014 69300
rect 69682 69244 69692 69300
rect 69748 69244 70252 69300
rect 70308 69244 70318 69300
rect 70578 69244 70588 69300
rect 70644 69244 76860 69300
rect 76916 69244 76926 69300
rect 0 69188 800 69216
rect 70252 69188 70308 69244
rect 79200 69188 80000 69216
rect 0 69132 2716 69188
rect 2772 69132 3500 69188
rect 3556 69132 3566 69188
rect 70252 69132 71148 69188
rect 71204 69132 71214 69188
rect 76514 69132 76524 69188
rect 76580 69132 77308 69188
rect 77364 69132 80000 69188
rect 0 69104 800 69132
rect 79200 69104 80000 69132
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 3042 68684 3052 68740
rect 3108 68684 67340 68740
rect 67396 68684 67676 68740
rect 67732 68684 67742 68740
rect 68674 68684 68684 68740
rect 68740 68684 76188 68740
rect 76244 68684 76254 68740
rect 1922 68572 1932 68628
rect 1988 68572 3500 68628
rect 3556 68572 3566 68628
rect 75954 68572 75964 68628
rect 76020 68572 77980 68628
rect 78036 68572 78046 68628
rect 0 68516 800 68544
rect 79200 68516 80000 68544
rect 0 68460 2716 68516
rect 2772 68460 2782 68516
rect 3154 68460 3164 68516
rect 3220 68460 66780 68516
rect 66836 68460 67788 68516
rect 67844 68460 67854 68516
rect 76402 68460 76412 68516
rect 76468 68460 77196 68516
rect 77252 68460 80000 68516
rect 0 68432 800 68460
rect 79200 68432 80000 68460
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 68562 68012 68572 68068
rect 68628 68012 70028 68068
rect 70084 68012 77868 68068
rect 77924 68012 77934 68068
rect 1708 67900 1820 67956
rect 1876 67900 1886 67956
rect 69458 67900 69468 67956
rect 69524 67900 76860 67956
rect 76916 67900 76926 67956
rect 0 67844 800 67872
rect 1708 67844 1764 67900
rect 79200 67844 80000 67872
rect 0 67788 1764 67844
rect 2258 67788 2268 67844
rect 2324 67788 66668 67844
rect 66724 67788 67116 67844
rect 67172 67788 67182 67844
rect 77298 67788 77308 67844
rect 77364 67788 77980 67844
rect 78036 67788 78046 67844
rect 78194 67788 78204 67844
rect 78260 67788 80000 67844
rect 0 67760 800 67788
rect 79200 67760 80000 67788
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 78082 67340 78092 67396
rect 78148 67340 78260 67396
rect 1596 67228 1932 67284
rect 1988 67228 1998 67284
rect 0 67172 800 67200
rect 1596 67172 1652 67228
rect 78204 67172 78260 67340
rect 79200 67172 80000 67200
rect 0 67116 1652 67172
rect 1810 67116 1820 67172
rect 1876 67116 3052 67172
rect 3108 67116 3118 67172
rect 67554 67116 67564 67172
rect 67620 67116 77868 67172
rect 77924 67116 77934 67172
rect 78204 67116 80000 67172
rect 0 67088 800 67116
rect 79200 67088 80000 67116
rect 63410 67004 63420 67060
rect 63476 67004 65996 67060
rect 66052 67004 66062 67060
rect 67666 67004 67676 67060
rect 67732 67004 68236 67060
rect 68292 67004 68302 67060
rect 77298 67004 77308 67060
rect 77364 67004 78092 67060
rect 78148 67004 78158 67060
rect 1922 66892 1932 66948
rect 1988 66892 2604 66948
rect 2660 66892 2670 66948
rect 67106 66892 67116 66948
rect 67172 66892 69356 66948
rect 69412 66892 77644 66948
rect 77700 66892 77710 66948
rect 68310 66668 68348 66724
rect 68404 66668 68414 66724
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 0 66500 800 66528
rect 79200 66500 80000 66528
rect 0 66444 1820 66500
rect 1876 66444 1886 66500
rect 68114 66444 68124 66500
rect 68180 66444 68796 66500
rect 68852 66444 68862 66500
rect 77970 66444 77980 66500
rect 78036 66444 80000 66500
rect 0 66416 800 66444
rect 79200 66416 80000 66444
rect 66994 66332 67004 66388
rect 67060 66332 67564 66388
rect 67620 66332 67630 66388
rect 68674 66332 68684 66388
rect 68740 66332 69244 66388
rect 69300 66332 69310 66388
rect 2258 66220 2268 66276
rect 2324 66220 8428 66276
rect 8372 66164 8428 66220
rect 55412 66220 63308 66276
rect 63364 66220 63868 66276
rect 63924 66220 63934 66276
rect 64530 66220 64540 66276
rect 64596 66220 64876 66276
rect 64932 66220 77756 66276
rect 77812 66220 77822 66276
rect 55412 66164 55468 66220
rect 8372 66108 55468 66164
rect 62514 66108 62524 66164
rect 62580 66108 65884 66164
rect 65940 66108 65950 66164
rect 2370 65996 2380 66052
rect 2436 65996 61964 66052
rect 62020 65996 62412 66052
rect 62468 65996 62478 66052
rect 65650 65996 65660 66052
rect 65716 65996 66164 66052
rect 67778 65996 67788 66052
rect 67844 65996 68572 66052
rect 68628 65996 68638 66052
rect 77298 65996 77308 66052
rect 77364 65996 78092 66052
rect 78148 65996 78158 66052
rect 66108 65940 66164 65996
rect 66098 65884 66108 65940
rect 66164 65884 66668 65940
rect 66724 65884 66734 65940
rect 0 65828 800 65856
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 79200 65828 80000 65856
rect 0 65772 1932 65828
rect 1988 65772 1998 65828
rect 65650 65772 65660 65828
rect 65716 65772 66220 65828
rect 66276 65772 66286 65828
rect 66434 65772 66444 65828
rect 66500 65772 67004 65828
rect 67060 65772 77756 65828
rect 77812 65772 77822 65828
rect 78194 65772 78204 65828
rect 78260 65772 80000 65828
rect 0 65744 800 65772
rect 79200 65744 80000 65772
rect 65986 65660 65996 65716
rect 66052 65660 66556 65716
rect 66612 65660 66622 65716
rect 68310 65660 68348 65716
rect 68404 65660 68414 65716
rect 61842 65548 61852 65604
rect 61908 65548 65884 65604
rect 65940 65548 65950 65604
rect 2034 65436 2044 65492
rect 2100 65436 8428 65492
rect 68450 65436 68460 65492
rect 68516 65436 68796 65492
rect 68852 65436 68862 65492
rect 8372 65380 8428 65436
rect 1922 65324 1932 65380
rect 1988 65324 2604 65380
rect 2660 65324 2670 65380
rect 8372 65324 61740 65380
rect 61796 65324 62300 65380
rect 62356 65324 62366 65380
rect 77298 65324 77308 65380
rect 77364 65324 77980 65380
rect 78036 65324 78046 65380
rect 0 65156 800 65184
rect 79200 65156 80000 65184
rect 0 65100 1820 65156
rect 1876 65100 2492 65156
rect 2548 65100 2558 65156
rect 78082 65100 78092 65156
rect 78148 65100 80000 65156
rect 0 65072 800 65100
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 79200 65072 80000 65100
rect 2258 64652 2268 64708
rect 2324 64652 60732 64708
rect 60788 64652 61404 64708
rect 61460 64652 61470 64708
rect 63522 64652 63532 64708
rect 63588 64652 64204 64708
rect 64260 64652 77756 64708
rect 77812 64652 77822 64708
rect 65762 64540 65772 64596
rect 65828 64540 66332 64596
rect 66388 64540 66398 64596
rect 68450 64540 68460 64596
rect 68516 64540 69356 64596
rect 69412 64540 69422 64596
rect 76626 64540 76636 64596
rect 76692 64540 78092 64596
rect 78148 64540 78158 64596
rect 0 64484 800 64512
rect 79200 64484 80000 64512
rect 0 64428 1932 64484
rect 1988 64428 1998 64484
rect 61506 64428 61516 64484
rect 61572 64428 65324 64484
rect 65380 64428 65390 64484
rect 67778 64428 67788 64484
rect 67844 64428 68012 64484
rect 68068 64428 68684 64484
rect 68740 64428 68750 64484
rect 77970 64428 77980 64484
rect 78036 64428 80000 64484
rect 0 64400 800 64428
rect 79200 64400 80000 64428
rect 65090 64316 65100 64372
rect 65156 64316 66444 64372
rect 66500 64316 66668 64372
rect 66724 64316 66734 64372
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 64530 64204 64540 64260
rect 64596 64204 64876 64260
rect 64932 64204 76860 64260
rect 76916 64204 76926 64260
rect 77298 64204 77308 64260
rect 77364 64204 77980 64260
rect 78036 64204 78046 64260
rect 59490 64092 59500 64148
rect 59556 64092 62188 64148
rect 62244 64092 65100 64148
rect 65156 64092 65166 64148
rect 65538 64092 65548 64148
rect 65604 64092 65884 64148
rect 65940 64092 65950 64148
rect 67666 64092 67676 64148
rect 67732 64092 68460 64148
rect 68516 64092 68526 64148
rect 1922 63980 1932 64036
rect 1988 63980 3500 64036
rect 3556 63980 3566 64036
rect 61170 63980 61180 64036
rect 61236 63980 63420 64036
rect 63476 63980 63486 64036
rect 66658 63980 66668 64036
rect 66724 63980 67452 64036
rect 67508 63980 67518 64036
rect 77410 63980 77420 64036
rect 77476 63980 77756 64036
rect 77812 63980 77822 64036
rect 2034 63868 2044 63924
rect 2100 63868 61068 63924
rect 61124 63868 61628 63924
rect 61684 63868 61694 63924
rect 63522 63868 63532 63924
rect 63588 63868 64428 63924
rect 64484 63868 64494 63924
rect 65090 63868 65100 63924
rect 65156 63868 65548 63924
rect 65604 63868 67004 63924
rect 67060 63868 67340 63924
rect 67396 63868 67406 63924
rect 76402 63868 76412 63924
rect 76468 63868 77196 63924
rect 77252 63868 77262 63924
rect 0 63812 800 63840
rect 77196 63812 77252 63868
rect 79200 63812 80000 63840
rect 0 63756 2716 63812
rect 2772 63756 2782 63812
rect 62514 63756 62524 63812
rect 62580 63756 63420 63812
rect 63476 63756 63644 63812
rect 63700 63756 63980 63812
rect 64036 63756 64046 63812
rect 77196 63756 80000 63812
rect 0 63728 800 63756
rect 79200 63728 80000 63756
rect 1698 63644 1708 63700
rect 1764 63644 2604 63700
rect 2660 63644 2670 63700
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 63298 63196 63308 63252
rect 63364 63196 63420 63252
rect 63476 63196 63486 63252
rect 78082 63196 78092 63252
rect 78148 63196 78158 63252
rect 0 63140 800 63168
rect 78092 63140 78148 63196
rect 79200 63140 80000 63168
rect 0 63084 1708 63140
rect 1764 63084 1774 63140
rect 2146 63084 2156 63140
rect 2212 63084 61404 63140
rect 61460 63084 61964 63140
rect 62020 63084 62030 63140
rect 63186 63084 63196 63140
rect 63252 63084 63644 63140
rect 63700 63084 63710 63140
rect 78092 63084 80000 63140
rect 0 63056 800 63084
rect 79200 63056 80000 63084
rect 77298 62972 77308 63028
rect 77364 62972 78092 63028
rect 78148 62972 78158 63028
rect 3154 62860 3164 62916
rect 3220 62860 59276 62916
rect 59332 62860 59836 62916
rect 59892 62860 59902 62916
rect 59378 62748 59388 62804
rect 59444 62748 63308 62804
rect 63364 62748 63374 62804
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 1922 62524 1932 62580
rect 1988 62524 1998 62580
rect 61506 62524 61516 62580
rect 61572 62524 62636 62580
rect 62692 62524 62702 62580
rect 68226 62524 68236 62580
rect 68292 62524 68796 62580
rect 68852 62524 77644 62580
rect 77700 62524 77710 62580
rect 77970 62524 77980 62580
rect 78036 62524 78046 62580
rect 0 62468 800 62496
rect 1932 62468 1988 62524
rect 77980 62468 78036 62524
rect 79200 62468 80000 62496
rect 0 62412 1988 62468
rect 65314 62412 65324 62468
rect 65380 62412 77756 62468
rect 77812 62412 77822 62468
rect 77980 62412 80000 62468
rect 0 62384 800 62412
rect 79200 62384 80000 62412
rect 59826 62300 59836 62356
rect 59892 62300 63868 62356
rect 63924 62300 63934 62356
rect 2370 62188 2380 62244
rect 2436 62188 59724 62244
rect 59780 62188 60284 62244
rect 60340 62188 60350 62244
rect 64306 62188 64316 62244
rect 64372 62188 68236 62244
rect 68292 62188 68302 62244
rect 77298 62188 77308 62244
rect 77364 62188 77980 62244
rect 78036 62188 78046 62244
rect 1922 62076 1932 62132
rect 1988 62076 2604 62132
rect 2660 62076 2670 62132
rect 63634 62076 63644 62132
rect 63700 62076 66108 62132
rect 66164 62076 66668 62132
rect 66724 62076 66734 62132
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 0 61796 800 61824
rect 79200 61796 80000 61824
rect 0 61740 1820 61796
rect 1876 61740 3052 61796
rect 3108 61740 3118 61796
rect 78082 61740 78092 61796
rect 78148 61740 80000 61796
rect 0 61712 800 61740
rect 79200 61712 80000 61740
rect 2258 61516 2268 61572
rect 2324 61516 8428 61572
rect 62738 61516 62748 61572
rect 62804 61516 64204 61572
rect 64260 61516 77420 61572
rect 77476 61516 77486 61572
rect 8372 61460 8428 61516
rect 1810 61404 1820 61460
rect 1876 61404 2604 61460
rect 2660 61404 2670 61460
rect 8372 61404 59724 61460
rect 59780 61404 60172 61460
rect 60228 61404 60238 61460
rect 61394 61404 61404 61460
rect 61460 61404 62076 61460
rect 62132 61348 62188 61460
rect 62962 61404 62972 61460
rect 63028 61404 63308 61460
rect 63364 61404 63374 61460
rect 77298 61404 77308 61460
rect 77364 61404 78092 61460
rect 78148 61404 78158 61460
rect 62132 61292 77868 61348
rect 77924 61292 77934 61348
rect 0 61124 800 61152
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 79200 61124 80000 61152
rect 0 61068 1932 61124
rect 1988 61068 1998 61124
rect 63382 61068 63420 61124
rect 63476 61068 63486 61124
rect 77970 61068 77980 61124
rect 78036 61068 80000 61124
rect 0 61040 800 61068
rect 79200 61040 80000 61068
rect 60274 60956 60284 61012
rect 60340 60956 62300 61012
rect 62356 60956 62366 61012
rect 60610 60844 60620 60900
rect 60676 60844 60956 60900
rect 61012 60844 62524 60900
rect 62580 60844 62590 60900
rect 63186 60844 63196 60900
rect 63252 60844 63532 60900
rect 63588 60844 63598 60900
rect 57586 60732 57596 60788
rect 57652 60732 60844 60788
rect 60900 60732 60910 60788
rect 61730 60732 61740 60788
rect 61796 60732 63084 60788
rect 63140 60732 63644 60788
rect 63700 60732 63710 60788
rect 2034 60620 2044 60676
rect 2100 60620 57484 60676
rect 57540 60620 58044 60676
rect 58100 60620 58110 60676
rect 58370 60620 58380 60676
rect 58436 60620 58828 60676
rect 58884 60620 59388 60676
rect 59444 60620 59454 60676
rect 59714 60620 59724 60676
rect 59780 60620 60396 60676
rect 60452 60620 61068 60676
rect 61124 60620 62076 60676
rect 62132 60620 62142 60676
rect 77298 60620 77308 60676
rect 77364 60620 78092 60676
rect 78148 60620 78158 60676
rect 61282 60508 61292 60564
rect 61348 60508 64540 60564
rect 64596 60508 64606 60564
rect 78194 60508 78204 60564
rect 78260 60508 78270 60564
rect 0 60452 800 60480
rect 78204 60452 78260 60508
rect 79200 60452 80000 60480
rect 0 60396 1708 60452
rect 1764 60396 1774 60452
rect 1922 60396 1932 60452
rect 1988 60396 2604 60452
rect 2660 60396 2670 60452
rect 78204 60396 80000 60452
rect 0 60368 800 60396
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 79200 60368 80000 60396
rect 61506 60172 61516 60228
rect 61572 60172 62076 60228
rect 62132 60172 77756 60228
rect 77812 60172 77822 60228
rect 2258 60060 2268 60116
rect 2324 60060 20188 60116
rect 59938 60060 59948 60116
rect 60004 60060 60956 60116
rect 61012 60060 61022 60116
rect 66658 60060 66668 60116
rect 66724 60060 67228 60116
rect 67284 60060 77644 60116
rect 77700 60060 77710 60116
rect 20132 60004 20188 60060
rect 2146 59948 2156 60004
rect 2212 59948 8428 60004
rect 20132 59948 57372 60004
rect 57428 59948 57932 60004
rect 57988 59948 57998 60004
rect 60610 59948 60620 60004
rect 60676 59948 66556 60004
rect 66612 59948 66622 60004
rect 8372 59892 8428 59948
rect 8372 59836 50428 59892
rect 57474 59836 57484 59892
rect 57540 59836 60172 59892
rect 60228 59836 60238 59892
rect 78082 59836 78092 59892
rect 78148 59836 78260 59892
rect 0 59780 800 59808
rect 50372 59780 50428 59836
rect 78204 59780 78260 59836
rect 79200 59780 80000 59808
rect 0 59724 1932 59780
rect 1988 59724 1998 59780
rect 50372 59724 58716 59780
rect 58772 59724 59276 59780
rect 59332 59724 59342 59780
rect 60274 59724 60284 59780
rect 60340 59724 61404 59780
rect 61460 59724 61470 59780
rect 76626 59724 76636 59780
rect 76692 59724 77980 59780
rect 78036 59724 78046 59780
rect 78204 59724 80000 59780
rect 0 59696 800 59724
rect 79200 59696 80000 59724
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 59602 59276 59612 59332
rect 59668 59276 59948 59332
rect 60004 59276 60014 59332
rect 1922 59164 1932 59220
rect 1988 59164 3500 59220
rect 3556 59164 3566 59220
rect 77298 59164 77308 59220
rect 77364 59164 78092 59220
rect 78148 59164 78158 59220
rect 0 59108 800 59136
rect 79200 59108 80000 59136
rect 0 59052 2716 59108
rect 2772 59052 2782 59108
rect 60050 59052 60060 59108
rect 60116 59052 60396 59108
rect 60452 59052 60462 59108
rect 76402 59052 76412 59108
rect 76468 59052 77196 59108
rect 77252 59052 80000 59108
rect 0 59024 800 59052
rect 79200 59024 80000 59052
rect 77970 58828 77980 58884
rect 78036 58828 78046 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 2146 58604 2156 58660
rect 2212 58604 3276 58660
rect 3332 58604 3342 58660
rect 2258 58492 2268 58548
rect 2324 58492 20188 58548
rect 59378 58492 59388 58548
rect 59444 58492 60396 58548
rect 60452 58492 77644 58548
rect 77700 58492 77710 58548
rect 0 58436 800 58464
rect 20132 58436 20188 58492
rect 77980 58436 78036 58828
rect 79200 58436 80000 58464
rect 0 58380 1708 58436
rect 1764 58380 2604 58436
rect 2660 58380 2670 58436
rect 3042 58380 3052 58436
rect 3108 58380 8428 58436
rect 20132 58380 56140 58436
rect 56196 58380 56700 58436
rect 56756 58380 56766 58436
rect 58482 58380 58492 58436
rect 58548 58380 59948 58436
rect 60004 58380 76860 58436
rect 76916 58380 76926 58436
rect 77980 58380 80000 58436
rect 0 58352 800 58380
rect 8372 58324 8428 58380
rect 79200 58352 80000 58380
rect 8372 58268 57260 58324
rect 57316 58268 57820 58324
rect 57876 58268 57886 58324
rect 77298 58268 77308 58324
rect 77364 58268 77980 58324
rect 78036 58268 78046 58324
rect 59826 58156 59836 58212
rect 59892 58156 77756 58212
rect 77812 58156 77822 58212
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 57586 57932 57596 57988
rect 57652 57932 57932 57988
rect 57988 57932 59500 57988
rect 59556 57932 59566 57988
rect 1922 57820 1932 57876
rect 1988 57820 1998 57876
rect 58482 57820 58492 57876
rect 58548 57820 59276 57876
rect 59332 57820 59342 57876
rect 78082 57820 78092 57876
rect 78148 57820 78260 57876
rect 0 57764 800 57792
rect 1932 57764 1988 57820
rect 78204 57764 78260 57820
rect 79200 57764 80000 57792
rect 0 57708 1988 57764
rect 57362 57708 57372 57764
rect 57428 57708 59332 57764
rect 78204 57708 80000 57764
rect 0 57680 800 57708
rect 59276 57652 59332 57708
rect 79200 57680 80000 57708
rect 55122 57596 55132 57652
rect 55188 57596 57820 57652
rect 57876 57596 57886 57652
rect 59266 57596 59276 57652
rect 59332 57596 59342 57652
rect 62738 57596 62748 57652
rect 62804 57596 63196 57652
rect 63252 57596 77868 57652
rect 77924 57596 77934 57652
rect 3266 57484 3276 57540
rect 3332 57484 55020 57540
rect 55076 57484 55580 57540
rect 55636 57484 55646 57540
rect 58146 57484 58156 57540
rect 58212 57484 59052 57540
rect 59108 57484 59118 57540
rect 77298 57484 77308 57540
rect 77364 57484 78092 57540
rect 78148 57484 78158 57540
rect 58258 57372 58268 57428
rect 58324 57372 62636 57428
rect 62692 57372 62702 57428
rect 58594 57260 58604 57316
rect 58660 57260 61292 57316
rect 61348 57260 61358 57316
rect 77970 57260 77980 57316
rect 78036 57260 78372 57316
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 59154 57148 59164 57204
rect 59220 57148 59836 57204
rect 59892 57148 59902 57204
rect 0 57092 800 57120
rect 78316 57092 78372 57260
rect 79200 57092 80000 57120
rect 0 57036 1820 57092
rect 1876 57036 3052 57092
rect 3108 57036 3118 57092
rect 78316 57036 80000 57092
rect 0 57008 800 57036
rect 79200 57008 80000 57036
rect 1922 56924 1932 56980
rect 1988 56924 2604 56980
rect 2660 56924 2670 56980
rect 56242 56924 56252 56980
rect 56308 56924 58044 56980
rect 58100 56924 58110 56980
rect 2706 56700 2716 56756
rect 2772 56700 56252 56756
rect 56308 56700 56700 56756
rect 56756 56700 56766 56756
rect 1810 56588 1820 56644
rect 1876 56588 2604 56644
rect 2660 56588 2670 56644
rect 77298 56588 77308 56644
rect 77364 56588 77980 56644
rect 78036 56588 78046 56644
rect 0 56420 800 56448
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 79200 56420 80000 56448
rect 0 56364 1932 56420
rect 1988 56364 1998 56420
rect 78082 56364 78092 56420
rect 78148 56364 80000 56420
rect 0 56336 800 56364
rect 79200 56336 80000 56364
rect 56802 56252 56812 56308
rect 56868 56252 57820 56308
rect 57876 56252 57886 56308
rect 56242 56140 56252 56196
rect 56308 56140 77756 56196
rect 77812 56140 77822 56196
rect 52210 56028 52220 56084
rect 52276 56028 55580 56084
rect 55636 56028 55646 56084
rect 58258 56028 58268 56084
rect 58324 56028 59052 56084
rect 59108 56028 59118 56084
rect 62132 56028 77644 56084
rect 77700 56028 77710 56084
rect 62132 55972 62188 56028
rect 2034 55916 2044 55972
rect 2100 55916 52108 55972
rect 52164 55916 52668 55972
rect 52724 55916 52734 55972
rect 56690 55916 56700 55972
rect 56756 55916 58716 55972
rect 58772 55916 62188 55972
rect 77298 55916 77308 55972
rect 77364 55916 78092 55972
rect 78148 55916 78158 55972
rect 0 55748 800 55776
rect 79200 55748 80000 55776
rect 0 55692 1820 55748
rect 1876 55692 1886 55748
rect 77970 55692 77980 55748
rect 78036 55692 80000 55748
rect 0 55664 800 55692
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 79200 55664 80000 55692
rect 78082 55468 78092 55524
rect 78148 55468 79268 55524
rect 79212 55412 79268 55468
rect 2258 55356 2268 55412
rect 2324 55356 50316 55412
rect 50372 55356 50876 55412
rect 50932 55356 50942 55412
rect 78988 55356 79268 55412
rect 52322 55244 52332 55300
rect 52388 55244 54124 55300
rect 54180 55244 54684 55300
rect 54740 55244 56924 55300
rect 56980 55244 56990 55300
rect 57698 55244 57708 55300
rect 57764 55244 58492 55300
rect 58548 55244 58558 55300
rect 54338 55132 54348 55188
rect 54404 55132 55580 55188
rect 55636 55132 55646 55188
rect 57250 55132 57260 55188
rect 57316 55132 58044 55188
rect 58100 55132 58110 55188
rect 0 55076 800 55104
rect 78988 55076 79044 55356
rect 79200 55076 80000 55104
rect 0 55020 1932 55076
rect 1988 55020 2492 55076
rect 2548 55020 2558 55076
rect 50418 55020 50428 55076
rect 50484 55020 55356 55076
rect 55412 55020 55422 55076
rect 56914 55020 56924 55076
rect 56980 55020 57708 55076
rect 57764 55020 57774 55076
rect 76626 55020 76636 55076
rect 76692 55020 77980 55076
rect 78036 55020 78046 55076
rect 78988 55020 80000 55076
rect 0 54992 800 55020
rect 79200 54992 80000 55020
rect 55794 54908 55804 54964
rect 55860 54908 56476 54964
rect 56532 54908 56542 54964
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 56578 54796 56588 54852
rect 56644 54796 57596 54852
rect 57652 54796 77868 54852
rect 77924 54796 77934 54852
rect 2034 54684 2044 54740
rect 2100 54684 52444 54740
rect 52500 54684 52780 54740
rect 52836 54684 52846 54740
rect 53554 54684 53564 54740
rect 53620 54684 53788 54740
rect 53844 54684 76860 54740
rect 76916 54684 76926 54740
rect 3042 54572 3052 54628
rect 3108 54572 51660 54628
rect 51716 54572 52108 54628
rect 52164 54572 52174 54628
rect 56914 54572 56924 54628
rect 56980 54572 77756 54628
rect 77812 54572 77822 54628
rect 1922 54460 1932 54516
rect 1988 54460 3500 54516
rect 3556 54460 3566 54516
rect 52882 54460 52892 54516
rect 52948 54460 54796 54516
rect 54852 54460 54862 54516
rect 55010 54460 55020 54516
rect 55076 54460 55580 54516
rect 55636 54460 55646 54516
rect 77298 54460 77308 54516
rect 77364 54460 78092 54516
rect 78148 54460 78158 54516
rect 0 54404 800 54432
rect 79200 54404 80000 54432
rect 0 54348 2716 54404
rect 2772 54348 2782 54404
rect 54674 54348 54684 54404
rect 54740 54348 55356 54404
rect 55412 54348 55422 54404
rect 76402 54348 76412 54404
rect 76468 54348 77196 54404
rect 77252 54348 80000 54404
rect 0 54320 800 54348
rect 79200 54320 80000 54348
rect 55234 54236 55244 54292
rect 55300 54236 55804 54292
rect 55860 54236 55870 54292
rect 54562 54124 54572 54180
rect 54628 54124 55132 54180
rect 55188 54124 55198 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 77970 53788 77980 53844
rect 78036 53788 78046 53844
rect 0 53732 800 53760
rect 77980 53732 78036 53788
rect 79200 53732 80000 53760
rect 0 53676 1708 53732
rect 1764 53676 2604 53732
rect 2660 53676 2670 53732
rect 52210 53676 52220 53732
rect 52276 53676 54684 53732
rect 54740 53676 54750 53732
rect 54898 53676 54908 53732
rect 54964 53676 55580 53732
rect 55636 53676 55646 53732
rect 55906 53676 55916 53732
rect 55972 53676 56140 53732
rect 56196 53676 57148 53732
rect 57204 53676 57214 53732
rect 62132 53676 77644 53732
rect 77700 53676 77710 53732
rect 77980 53676 80000 53732
rect 0 53648 800 53676
rect 62132 53620 62188 53676
rect 79200 53648 80000 53676
rect 2146 53564 2156 53620
rect 2212 53564 46956 53620
rect 47012 53564 47022 53620
rect 52770 53564 52780 53620
rect 52836 53564 53452 53620
rect 53508 53564 62188 53620
rect 1810 53452 1820 53508
rect 1876 53452 3052 53508
rect 3108 53452 3118 53508
rect 8372 53452 47740 53508
rect 47796 53452 48300 53508
rect 48356 53452 48366 53508
rect 77298 53452 77308 53508
rect 77364 53452 78092 53508
rect 78148 53452 78158 53508
rect 8372 53396 8428 53452
rect 2258 53340 2268 53396
rect 2324 53340 8428 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 1922 53116 1932 53172
rect 1988 53116 1998 53172
rect 52658 53116 52668 53172
rect 52724 53116 53228 53172
rect 53284 53116 54460 53172
rect 54516 53116 54526 53172
rect 57810 53116 57820 53172
rect 57876 53116 58380 53172
rect 58436 53116 58446 53172
rect 0 53060 800 53088
rect 1932 53060 1988 53116
rect 79200 53060 80000 53088
rect 0 53004 1988 53060
rect 2146 53004 2156 53060
rect 2212 53004 48748 53060
rect 48804 53004 48814 53060
rect 50306 53004 50316 53060
rect 50372 53004 54348 53060
rect 54404 53004 54414 53060
rect 78194 53004 78204 53060
rect 78260 53004 80000 53060
rect 0 52976 800 53004
rect 79200 52976 80000 53004
rect 48402 52892 48412 52948
rect 48468 52892 52892 52948
rect 52948 52892 52958 52948
rect 56018 52892 56028 52948
rect 56084 52892 56588 52948
rect 56644 52892 56654 52948
rect 2706 52780 2716 52836
rect 2772 52780 50204 52836
rect 50260 52780 50764 52836
rect 50820 52780 50830 52836
rect 51874 52780 51884 52836
rect 51940 52780 52444 52836
rect 52500 52780 53116 52836
rect 53172 52780 54124 52836
rect 54180 52780 54190 52836
rect 77298 52780 77308 52836
rect 77364 52780 77980 52836
rect 78036 52780 78046 52836
rect 53330 52668 53340 52724
rect 53396 52668 56588 52724
rect 56644 52668 56654 52724
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 0 52388 800 52416
rect 79200 52388 80000 52416
rect 0 52332 1820 52388
rect 1876 52332 1886 52388
rect 52658 52332 52668 52388
rect 52724 52332 60284 52388
rect 60340 52332 60350 52388
rect 78082 52332 78092 52388
rect 78148 52332 80000 52388
rect 0 52304 800 52332
rect 79200 52304 80000 52332
rect 46946 52220 46956 52276
rect 47012 52220 47516 52276
rect 47572 52220 47582 52276
rect 48738 52220 48748 52276
rect 48804 52220 49308 52276
rect 49364 52220 49374 52276
rect 52546 52220 52556 52276
rect 52612 52220 59164 52276
rect 59220 52220 59230 52276
rect 60386 52220 60396 52276
rect 60452 52220 61404 52276
rect 61460 52220 77644 52276
rect 77700 52220 77710 52276
rect 56242 52108 56252 52164
rect 56308 52108 56812 52164
rect 56868 52108 57260 52164
rect 57316 52108 57484 52164
rect 57540 52108 57550 52164
rect 59266 52108 59276 52164
rect 59332 52108 59836 52164
rect 59892 52108 77756 52164
rect 77812 52108 77822 52164
rect 1810 51996 1820 52052
rect 1876 51996 2604 52052
rect 2660 51996 2670 52052
rect 47058 51996 47068 52052
rect 47124 51996 52220 52052
rect 52276 51996 52286 52052
rect 2146 51884 2156 51940
rect 2212 51884 49196 51940
rect 49252 51884 49262 51940
rect 51986 51884 51996 51940
rect 52052 51884 53228 51940
rect 53284 51884 53294 51940
rect 77298 51884 77308 51940
rect 77364 51884 78092 51940
rect 78148 51884 78158 51940
rect 0 51716 800 51744
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 79200 51716 80000 51744
rect 0 51660 1932 51716
rect 1988 51660 1998 51716
rect 77970 51660 77980 51716
rect 78036 51660 80000 51716
rect 0 51632 800 51660
rect 79200 51632 80000 51660
rect 48850 51548 48860 51604
rect 48916 51548 52164 51604
rect 53666 51548 53676 51604
rect 53732 51548 56140 51604
rect 56196 51548 56206 51604
rect 57810 51548 57820 51604
rect 57876 51548 58604 51604
rect 58660 51548 58670 51604
rect 52108 51492 52164 51548
rect 52098 51436 52108 51492
rect 52164 51436 52174 51492
rect 52658 51436 52668 51492
rect 52724 51436 77756 51492
rect 77812 51436 77822 51492
rect 55682 51324 55692 51380
rect 55748 51324 56364 51380
rect 56420 51324 57148 51380
rect 57204 51324 57484 51380
rect 57540 51324 57550 51380
rect 77298 51212 77308 51268
rect 77364 51212 77980 51268
rect 78036 51212 78046 51268
rect 59378 51100 59388 51156
rect 59444 51100 60172 51156
rect 60228 51100 60238 51156
rect 0 51044 800 51072
rect 79200 51044 80000 51072
rect 0 50988 1820 51044
rect 1876 50988 1886 51044
rect 78082 50988 78092 51044
rect 78148 50988 80000 51044
rect 0 50960 800 50988
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 79200 50960 80000 50988
rect 70018 50764 70028 50820
rect 70084 50764 70700 50820
rect 70756 50764 77420 50820
rect 77476 50764 77486 50820
rect 4162 50652 4172 50708
rect 4228 50652 68684 50708
rect 68740 50652 69356 50708
rect 69412 50652 69422 50708
rect 77298 50652 77308 50708
rect 77364 50652 78092 50708
rect 78148 50652 78158 50708
rect 51762 50540 51772 50596
rect 51828 50540 52332 50596
rect 52388 50540 77644 50596
rect 77700 50540 77710 50596
rect 49746 50428 49756 50484
rect 49812 50428 50652 50484
rect 50708 50428 50718 50484
rect 77970 50428 77980 50484
rect 78036 50428 78046 50484
rect 0 50372 800 50400
rect 77980 50372 78036 50428
rect 79200 50372 80000 50400
rect 0 50316 1932 50372
rect 1988 50316 1998 50372
rect 50530 50316 50540 50372
rect 50596 50316 51772 50372
rect 51828 50316 51838 50372
rect 55412 50316 77756 50372
rect 77812 50316 77822 50372
rect 77980 50316 80000 50372
rect 0 50288 800 50316
rect 1698 50204 1708 50260
rect 1764 50204 3052 50260
rect 3108 50204 3118 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 50978 50092 50988 50148
rect 51044 50092 53452 50148
rect 53508 50092 53518 50148
rect 55412 50036 55468 50316
rect 79200 50288 80000 50316
rect 46610 49980 46620 50036
rect 46676 49980 51212 50036
rect 51268 49980 51278 50036
rect 51986 49980 51996 50036
rect 52052 49980 55468 50036
rect 70242 49980 70252 50036
rect 70308 49980 70318 50036
rect 2146 49868 2156 49924
rect 2212 49868 51716 49924
rect 3042 49756 3052 49812
rect 3108 49756 47964 49812
rect 48020 49756 48030 49812
rect 0 49700 800 49728
rect 51660 49700 51716 49868
rect 52108 49868 68012 49924
rect 68068 49868 68078 49924
rect 52108 49700 52164 49868
rect 68898 49756 68908 49812
rect 68964 49756 69244 49812
rect 69300 49756 69580 49812
rect 69636 49756 69916 49812
rect 69972 49756 69982 49812
rect 70252 49700 70308 49980
rect 78082 49756 78092 49812
rect 78148 49756 78260 49812
rect 78204 49700 78260 49756
rect 79200 49700 80000 49728
rect 0 49644 2716 49700
rect 2772 49644 2782 49700
rect 2930 49644 2940 49700
rect 2996 49644 46508 49700
rect 46564 49644 47068 49700
rect 47124 49644 47134 49700
rect 49746 49644 49756 49700
rect 49812 49644 50876 49700
rect 50932 49644 51436 49700
rect 51492 49644 51502 49700
rect 51660 49644 52164 49700
rect 69580 49644 70028 49700
rect 70084 49644 70700 49700
rect 70756 49644 70766 49700
rect 77298 49644 77308 49700
rect 77364 49644 77980 49700
rect 78036 49644 78046 49700
rect 78204 49644 80000 49700
rect 0 49616 800 49644
rect 69580 49588 69636 49644
rect 79200 49616 80000 49644
rect 1810 49532 1820 49588
rect 1876 49532 3500 49588
rect 3556 49532 3566 49588
rect 49186 49532 49196 49588
rect 49252 49532 50428 49588
rect 50484 49532 50988 49588
rect 51044 49532 51054 49588
rect 51650 49532 51660 49588
rect 51716 49532 52220 49588
rect 52276 49532 52286 49588
rect 69570 49532 69580 49588
rect 69636 49532 69646 49588
rect 50306 49420 50316 49476
rect 50372 49420 51996 49476
rect 52052 49420 52062 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 48066 49196 48076 49252
rect 48132 49196 49980 49252
rect 50036 49196 50046 49252
rect 47954 49084 47964 49140
rect 48020 49084 48524 49140
rect 48580 49084 48590 49140
rect 68002 49084 68012 49140
rect 68068 49084 68572 49140
rect 68628 49084 68638 49140
rect 0 49028 800 49056
rect 79200 49028 80000 49056
rect 0 48972 1708 49028
rect 1764 48972 1774 49028
rect 49858 48972 49868 49028
rect 49924 48972 50428 49028
rect 50484 48972 50494 49028
rect 55412 48972 77756 49028
rect 77812 48972 77822 49028
rect 77970 48972 77980 49028
rect 78036 48972 80000 49028
rect 0 48944 800 48972
rect 55412 48804 55468 48972
rect 79200 48944 80000 48972
rect 48626 48748 48636 48804
rect 48692 48748 49420 48804
rect 49476 48748 49486 48804
rect 49858 48748 49868 48804
rect 49924 48748 50316 48804
rect 50372 48748 50382 48804
rect 50530 48748 50540 48804
rect 50596 48748 51100 48804
rect 51156 48748 55468 48804
rect 68114 48748 68124 48804
rect 68180 48748 69804 48804
rect 69860 48748 69870 48804
rect 77298 48748 77308 48804
rect 77364 48748 78092 48804
rect 78148 48748 78158 48804
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 68786 48412 68796 48468
rect 68852 48412 69356 48468
rect 69412 48412 77756 48468
rect 77812 48412 77822 48468
rect 0 48356 800 48384
rect 79200 48356 80000 48384
rect 0 48300 1820 48356
rect 1876 48300 1886 48356
rect 69458 48300 69468 48356
rect 69524 48300 69916 48356
rect 69972 48300 69982 48356
rect 78082 48300 78092 48356
rect 78148 48300 80000 48356
rect 0 48272 800 48300
rect 79200 48272 80000 48300
rect 3042 48188 3052 48244
rect 3108 48188 3612 48244
rect 3668 48188 3678 48244
rect 2258 48076 2268 48132
rect 2324 48076 47292 48132
rect 47348 48076 48412 48132
rect 48468 48076 48478 48132
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 0 47684 800 47712
rect 79200 47684 80000 47712
rect 0 47628 2156 47684
rect 2212 47628 2222 47684
rect 76066 47628 76076 47684
rect 76132 47628 80000 47684
rect 0 47600 800 47628
rect 79200 47600 80000 47628
rect 47506 47292 47516 47348
rect 47572 47292 47852 47348
rect 47908 47292 48188 47348
rect 48244 47292 48972 47348
rect 49028 47292 49038 47348
rect 3602 47180 3612 47236
rect 3668 47180 47180 47236
rect 47236 47180 47246 47236
rect 48514 47180 48524 47236
rect 48580 47180 74620 47236
rect 74676 47180 74686 47236
rect 77858 47068 77868 47124
rect 77924 47068 77934 47124
rect 0 47012 800 47040
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 77868 47012 77924 47068
rect 79200 47012 80000 47040
rect 0 46956 2044 47012
rect 2100 46956 2110 47012
rect 77868 46956 80000 47012
rect 0 46928 800 46956
rect 79200 46928 80000 46956
rect 3714 46732 3724 46788
rect 3780 46732 46508 46788
rect 46564 46732 46574 46788
rect 47842 46732 47852 46788
rect 47908 46732 76972 46788
rect 77028 46732 77038 46788
rect 3042 46620 3052 46676
rect 3108 46620 3612 46676
rect 3668 46620 3678 46676
rect 46050 46508 46060 46564
rect 46116 46508 46844 46564
rect 46900 46508 47628 46564
rect 47684 46508 48300 46564
rect 48356 46508 48366 46564
rect 0 46340 800 46368
rect 79200 46340 80000 46368
rect 0 46284 2156 46340
rect 2212 46284 2222 46340
rect 76066 46284 76076 46340
rect 76132 46284 80000 46340
rect 0 46256 800 46284
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 79200 46256 80000 46284
rect 3490 45836 3500 45892
rect 3556 45836 3566 45892
rect 46844 45836 47740 45892
rect 47796 45836 48076 45892
rect 48132 45836 48142 45892
rect 0 45668 800 45696
rect 3500 45668 3556 45836
rect 46844 45780 46900 45836
rect 46162 45724 46172 45780
rect 46228 45724 46844 45780
rect 46900 45724 46910 45780
rect 47170 45724 47180 45780
rect 47236 45724 74620 45780
rect 74676 45724 74686 45780
rect 79200 45668 80000 45696
rect 0 45612 2044 45668
rect 2100 45612 2110 45668
rect 3500 45612 45836 45668
rect 45892 45612 45902 45668
rect 46498 45612 46508 45668
rect 46564 45612 74732 45668
rect 74788 45612 75292 45668
rect 75348 45612 75358 45668
rect 76178 45612 76188 45668
rect 76244 45612 80000 45668
rect 0 45584 800 45612
rect 79200 45584 80000 45612
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 3490 45276 3500 45332
rect 3556 45276 44380 45332
rect 44436 45276 44446 45332
rect 3602 45164 3612 45220
rect 3668 45164 45276 45220
rect 45332 45164 45342 45220
rect 43922 45052 43932 45108
rect 43988 45052 44604 45108
rect 44660 45052 44670 45108
rect 45602 45052 45612 45108
rect 45668 45052 46284 45108
rect 46340 45052 46956 45108
rect 47012 45052 47022 45108
rect 0 44996 800 45024
rect 44604 44996 44660 45052
rect 79200 44996 80000 45024
rect 0 44940 2156 44996
rect 2212 44940 2222 44996
rect 3042 44940 3052 44996
rect 3108 44940 3612 44996
rect 3668 44940 43708 44996
rect 43764 44940 43774 44996
rect 44604 44940 46396 44996
rect 46452 44940 46462 44996
rect 77746 44940 77756 44996
rect 77812 44940 80000 44996
rect 0 44912 800 44940
rect 79200 44912 80000 44940
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 0 44324 800 44352
rect 79200 44324 80000 44352
rect 0 44268 2044 44324
rect 2100 44268 2110 44324
rect 76066 44268 76076 44324
rect 76132 44268 80000 44324
rect 0 44240 800 44268
rect 79200 44240 80000 44268
rect 44034 44156 44044 44212
rect 44100 44156 44604 44212
rect 44660 44156 45276 44212
rect 45332 44156 45500 44212
rect 45556 44156 45566 44212
rect 45826 44156 45836 44212
rect 45892 44156 74620 44212
rect 74676 44156 74686 44212
rect 3042 44044 3052 44100
rect 3108 44044 3500 44100
rect 3556 44044 42924 44100
rect 42980 44044 42990 44100
rect 46722 44044 46732 44100
rect 46788 44044 77084 44100
rect 77140 44044 77150 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 44370 43708 44380 43764
rect 44436 43708 76524 43764
rect 76580 43708 76590 43764
rect 77858 43708 77868 43764
rect 77924 43708 77934 43764
rect 0 43652 800 43680
rect 77868 43652 77924 43708
rect 79200 43652 80000 43680
rect 0 43596 2156 43652
rect 2212 43596 2222 43652
rect 77868 43596 80000 43652
rect 0 43568 800 43596
rect 79200 43568 80000 43596
rect 3042 43372 3052 43428
rect 3108 43372 3612 43428
rect 3668 43372 42252 43428
rect 42308 43372 42318 43428
rect 42466 43372 42476 43428
rect 42532 43372 43260 43428
rect 43316 43372 44268 43428
rect 44324 43372 44828 43428
rect 44884 43372 44894 43428
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 0 42980 800 43008
rect 79200 42980 80000 43008
rect 0 42924 2044 42980
rect 2100 42924 2110 42980
rect 77858 42924 77868 42980
rect 77924 42924 80000 42980
rect 0 42896 800 42924
rect 79200 42896 80000 42924
rect 41906 42700 41916 42756
rect 41972 42700 42588 42756
rect 42644 42700 43372 42756
rect 43428 42700 43708 42756
rect 43652 42644 43708 42700
rect 43652 42588 44044 42644
rect 44100 42588 44110 42644
rect 3042 42476 3052 42532
rect 3108 42476 3500 42532
rect 3556 42476 41692 42532
rect 41748 42476 41758 42532
rect 43698 42476 43708 42532
rect 43764 42476 76412 42532
rect 76468 42476 76478 42532
rect 0 42308 800 42336
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 79200 42308 80000 42336
rect 0 42252 2156 42308
rect 2212 42252 2222 42308
rect 77868 42252 80000 42308
rect 0 42224 800 42252
rect 77868 41972 77924 42252
rect 79200 42224 80000 42252
rect 77746 41916 77756 41972
rect 77812 41916 77924 41972
rect 3042 41804 3052 41860
rect 3108 41804 3612 41860
rect 3668 41804 41020 41860
rect 41076 41804 41086 41860
rect 42018 41804 42028 41860
rect 42084 41804 42924 41860
rect 42980 41804 43484 41860
rect 43540 41804 43932 41860
rect 43988 41804 43998 41860
rect 0 41636 800 41664
rect 79200 41636 80000 41664
rect 0 41580 2044 41636
rect 2100 41580 2110 41636
rect 76066 41580 76076 41636
rect 76132 41580 80000 41636
rect 0 41552 800 41580
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 79200 41552 80000 41580
rect 42354 41020 42364 41076
rect 42420 41020 74620 41076
rect 74676 41020 74686 41076
rect 0 40964 800 40992
rect 79200 40964 80000 40992
rect 0 40908 2156 40964
rect 2212 40908 2222 40964
rect 3042 40908 3052 40964
rect 3108 40908 3500 40964
rect 3556 40908 40236 40964
rect 40292 40908 40302 40964
rect 40562 40908 40572 40964
rect 40628 40908 41356 40964
rect 41412 40908 42140 40964
rect 42196 40908 42812 40964
rect 42868 40908 42878 40964
rect 43026 40908 43036 40964
rect 43092 40908 76636 40964
rect 76692 40908 76702 40964
rect 77746 40908 77756 40964
rect 77812 40908 80000 40964
rect 0 40880 800 40908
rect 79200 40880 80000 40908
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 41906 40460 41916 40516
rect 41972 40460 76860 40516
rect 76916 40460 77196 40516
rect 77252 40460 77262 40516
rect 3042 40348 3052 40404
rect 3108 40348 3612 40404
rect 3668 40348 39340 40404
rect 39396 40348 39406 40404
rect 40562 40348 40572 40404
rect 40628 40348 41580 40404
rect 41636 40348 42364 40404
rect 42420 40348 42430 40404
rect 75954 40348 75964 40404
rect 76020 40348 76030 40404
rect 0 40292 800 40320
rect 75964 40292 76020 40348
rect 79200 40292 80000 40320
rect 0 40236 2044 40292
rect 2100 40236 2110 40292
rect 75964 40236 80000 40292
rect 0 40208 800 40236
rect 79200 40208 80000 40236
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 0 39620 800 39648
rect 79200 39620 80000 39648
rect 0 39564 2156 39620
rect 2212 39564 2222 39620
rect 77746 39564 77756 39620
rect 77812 39564 80000 39620
rect 0 39536 800 39564
rect 79200 39536 80000 39564
rect 3042 39452 3052 39508
rect 3108 39452 3612 39508
rect 3668 39452 38780 39508
rect 38836 39452 38846 39508
rect 39106 39452 39116 39508
rect 39172 39452 39676 39508
rect 39732 39452 39742 39508
rect 40898 39452 40908 39508
rect 40964 39452 74620 39508
rect 74676 39452 74686 39508
rect 39116 39396 39172 39452
rect 38322 39340 38332 39396
rect 38388 39340 38892 39396
rect 38948 39340 39172 39396
rect 40002 39340 40012 39396
rect 40068 39340 76860 39396
rect 76916 39340 76926 39396
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 74722 39004 74732 39060
rect 74788 39004 75292 39060
rect 75348 39004 75358 39060
rect 0 38948 800 38976
rect 74732 38948 74788 39004
rect 79200 38948 80000 38976
rect 0 38892 2156 38948
rect 2212 38892 2222 38948
rect 39778 38892 39788 38948
rect 39844 38892 74788 38948
rect 76178 38892 76188 38948
rect 76244 38892 80000 38948
rect 0 38864 800 38892
rect 79200 38864 80000 38892
rect 3042 38780 3052 38836
rect 3108 38780 3612 38836
rect 3668 38780 38332 38836
rect 38388 38780 38398 38836
rect 38658 38780 38668 38836
rect 38724 38780 39564 38836
rect 39620 38780 40684 38836
rect 40740 38780 40750 38836
rect 38668 38724 38724 38780
rect 37874 38668 37884 38724
rect 37940 38668 38724 38724
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 0 38276 800 38304
rect 79200 38276 80000 38304
rect 0 38220 2044 38276
rect 2100 38220 2110 38276
rect 76066 38220 76076 38276
rect 76132 38220 80000 38276
rect 0 38192 800 38220
rect 79200 38192 80000 38220
rect 37986 37884 37996 37940
rect 38052 37884 38668 37940
rect 38724 37884 39452 37940
rect 39508 37884 39518 37940
rect 3042 37772 3052 37828
rect 3108 37772 3612 37828
rect 3668 37772 37660 37828
rect 37716 37772 37726 37828
rect 38994 37772 39004 37828
rect 39060 37772 74620 37828
rect 74676 37772 74686 37828
rect 0 37604 800 37632
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 79200 37604 80000 37632
rect 0 37548 2156 37604
rect 2212 37548 2222 37604
rect 77746 37548 77756 37604
rect 77812 37548 80000 37604
rect 0 37520 800 37548
rect 79200 37520 80000 37548
rect 38322 37324 38332 37380
rect 38388 37324 76636 37380
rect 76692 37324 76860 37380
rect 76916 37324 76926 37380
rect 36530 37100 36540 37156
rect 36596 37100 37212 37156
rect 37268 37100 37996 37156
rect 38052 37100 38332 37156
rect 38388 37100 38398 37156
rect 3042 36988 3052 37044
rect 3108 36988 3612 37044
rect 3668 36988 36988 37044
rect 37044 36988 37054 37044
rect 76066 36988 76076 37044
rect 76132 36988 76142 37044
rect 0 36932 800 36960
rect 76076 36932 76132 36988
rect 79200 36932 80000 36960
rect 0 36876 2044 36932
rect 2100 36876 2110 36932
rect 76076 36876 80000 36932
rect 0 36848 800 36876
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 79200 36848 80000 36876
rect 35858 36316 35868 36372
rect 35924 36316 36652 36372
rect 36708 36316 37548 36372
rect 37604 36316 38780 36372
rect 38836 36316 38846 36372
rect 0 36260 800 36288
rect 79200 36260 80000 36288
rect 0 36204 2156 36260
rect 2212 36204 2222 36260
rect 3042 36204 3052 36260
rect 3108 36204 3612 36260
rect 3668 36204 36316 36260
rect 36372 36204 36382 36260
rect 37874 36204 37884 36260
rect 37940 36204 74620 36260
rect 74676 36204 74686 36260
rect 77746 36204 77756 36260
rect 77812 36204 80000 36260
rect 0 36176 800 36204
rect 79200 36176 80000 36204
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 3042 35756 3052 35812
rect 3108 35756 3612 35812
rect 3668 35756 35532 35812
rect 35588 35756 35598 35812
rect 35858 35756 35868 35812
rect 35924 35756 36764 35812
rect 36820 35756 36830 35812
rect 36978 35756 36988 35812
rect 37044 35756 76860 35812
rect 76916 35756 77196 35812
rect 77252 35756 77262 35812
rect 36764 35700 36820 35756
rect 34962 35644 34972 35700
rect 35028 35644 35308 35700
rect 35364 35644 36092 35700
rect 36148 35644 36158 35700
rect 36764 35644 37436 35700
rect 37492 35644 37502 35700
rect 0 35588 800 35616
rect 79200 35588 80000 35616
rect 0 35532 2044 35588
rect 2100 35532 2110 35588
rect 4834 35532 4844 35588
rect 4900 35532 5404 35588
rect 5460 35532 34188 35588
rect 34244 35532 34254 35588
rect 76066 35532 76076 35588
rect 76132 35532 80000 35588
rect 0 35504 800 35532
rect 79200 35504 80000 35532
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 0 34916 800 34944
rect 79200 34916 80000 34944
rect 0 34860 3836 34916
rect 3892 34860 3902 34916
rect 33730 34860 33740 34916
rect 33796 34860 34524 34916
rect 34580 34860 35196 34916
rect 35252 34860 35262 34916
rect 77746 34860 77756 34916
rect 77812 34860 80000 34916
rect 0 34832 800 34860
rect 79200 34832 80000 34860
rect 36306 34748 36316 34804
rect 36372 34748 74620 34804
rect 74676 34748 74686 34804
rect 3042 34636 3052 34692
rect 3108 34636 4060 34692
rect 4116 34636 34636 34692
rect 34692 34636 34702 34692
rect 35410 34636 35420 34692
rect 35476 34636 76860 34692
rect 76916 34636 76926 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 74722 34300 74732 34356
rect 74788 34300 75292 34356
rect 75348 34300 75358 34356
rect 0 34244 800 34272
rect 74732 34244 74788 34300
rect 79200 34244 80000 34272
rect 0 34188 2156 34244
rect 2212 34188 2222 34244
rect 35074 34188 35084 34244
rect 35140 34188 74788 34244
rect 76178 34188 76188 34244
rect 76244 34188 80000 34244
rect 0 34160 800 34188
rect 79200 34160 80000 34188
rect 32946 34076 32956 34132
rect 33012 34076 33964 34132
rect 34020 34076 34860 34132
rect 34916 34076 34926 34132
rect 3042 33852 3052 33908
rect 3108 33852 3612 33908
rect 3668 33852 33628 33908
rect 33684 33852 33694 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 76066 33628 76076 33684
rect 76132 33628 76142 33684
rect 0 33572 800 33600
rect 76076 33572 76132 33628
rect 79200 33572 80000 33600
rect 0 33516 2044 33572
rect 2100 33516 2110 33572
rect 76076 33516 80000 33572
rect 0 33488 800 33516
rect 79200 33488 80000 33516
rect 32498 33292 32508 33348
rect 32564 33292 33180 33348
rect 33236 33292 34076 33348
rect 34132 33292 34142 33348
rect 3042 33068 3052 33124
rect 3108 33068 3612 33124
rect 3668 33068 32956 33124
rect 33012 33068 33022 33124
rect 34402 33068 34412 33124
rect 34468 33068 74620 33124
rect 74676 33068 74686 33124
rect 0 32900 800 32928
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 79200 32900 80000 32928
rect 0 32844 2156 32900
rect 2212 32844 2222 32900
rect 77746 32844 77756 32900
rect 77812 32844 80000 32900
rect 0 32816 800 32844
rect 79200 32816 80000 32844
rect 33954 32620 33964 32676
rect 34020 32620 76636 32676
rect 76692 32620 76702 32676
rect 31892 32508 32508 32564
rect 32564 32508 33404 32564
rect 33460 32508 33628 32564
rect 33684 32508 33694 32564
rect 31892 32452 31948 32508
rect 31714 32396 31724 32452
rect 31780 32396 31948 32452
rect 3042 32284 3052 32340
rect 3108 32284 3612 32340
rect 3668 32284 32172 32340
rect 32228 32284 32238 32340
rect 0 32228 800 32256
rect 79200 32228 80000 32256
rect 0 32172 2044 32228
rect 2100 32172 2110 32228
rect 76066 32172 76076 32228
rect 76132 32172 80000 32228
rect 0 32144 800 32172
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 79200 32144 80000 32172
rect 31154 31612 31164 31668
rect 31220 31612 31948 31668
rect 32004 31612 32620 31668
rect 32676 31612 33852 31668
rect 33908 31612 33918 31668
rect 0 31556 800 31584
rect 79200 31556 80000 31584
rect 0 31500 2156 31556
rect 2212 31500 2222 31556
rect 3042 31500 3052 31556
rect 3108 31500 3612 31556
rect 3668 31500 31612 31556
rect 31668 31500 31678 31556
rect 32946 31500 32956 31556
rect 33012 31500 74620 31556
rect 74676 31500 74686 31556
rect 77746 31500 77756 31556
rect 77812 31500 80000 31556
rect 0 31472 800 31500
rect 79200 31472 80000 31500
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 3042 31052 3052 31108
rect 3108 31052 3612 31108
rect 3668 31052 30940 31108
rect 30996 31052 31006 31108
rect 32274 31052 32284 31108
rect 32340 31052 76860 31108
rect 76916 31052 77196 31108
rect 77252 31052 77262 31108
rect 31266 30940 31276 30996
rect 31332 30940 32060 30996
rect 32116 30940 32732 30996
rect 32788 30940 32798 30996
rect 0 30884 800 30912
rect 79200 30884 80000 30912
rect 0 30828 2156 30884
rect 2212 30828 2222 30884
rect 4834 30828 4844 30884
rect 4900 30828 5404 30884
rect 5460 30828 29596 30884
rect 29652 30828 29662 30884
rect 76066 30828 76076 30884
rect 76132 30828 80000 30884
rect 0 30800 800 30828
rect 79200 30800 80000 30828
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 0 30212 800 30240
rect 79200 30212 80000 30240
rect 0 30156 3836 30212
rect 3892 30156 3902 30212
rect 77746 30156 77756 30212
rect 77812 30156 80000 30212
rect 0 30128 800 30156
rect 79200 30128 80000 30156
rect 31602 30044 31612 30100
rect 31668 30044 74620 30100
rect 74676 30044 74686 30100
rect 3042 29932 3052 29988
rect 3108 29932 4060 29988
rect 4116 29932 30044 29988
rect 30100 29932 30110 29988
rect 30706 29932 30716 29988
rect 30772 29932 76860 29988
rect 76916 29932 76926 29988
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 74722 29596 74732 29652
rect 74788 29596 75292 29652
rect 75348 29596 75358 29652
rect 0 29540 800 29568
rect 74732 29540 74788 29596
rect 79200 29540 80000 29568
rect 0 29484 2156 29540
rect 2212 29484 2222 29540
rect 30818 29484 30828 29540
rect 30884 29484 74788 29540
rect 76178 29484 76188 29540
rect 76244 29484 80000 29540
rect 0 29456 800 29484
rect 79200 29456 80000 29484
rect 29922 29372 29932 29428
rect 29988 29372 30380 29428
rect 30436 29372 30604 29428
rect 30660 29372 30670 29428
rect 28242 29260 28252 29316
rect 28308 29260 29036 29316
rect 29092 29260 29102 29316
rect 3042 29148 3052 29204
rect 3108 29148 3612 29204
rect 3668 29148 28700 29204
rect 28756 29148 28766 29204
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 0 28868 800 28896
rect 79200 28868 80000 28896
rect 0 28812 2044 28868
rect 2100 28812 2110 28868
rect 76066 28812 76076 28868
rect 76132 28812 80000 28868
rect 0 28784 800 28812
rect 79200 28784 80000 28812
rect 3042 28588 3052 28644
rect 3108 28588 3612 28644
rect 3668 28588 28252 28644
rect 28308 28588 28318 28644
rect 29026 28588 29036 28644
rect 29092 28588 29708 28644
rect 29764 28588 30380 28644
rect 30436 28588 30446 28644
rect 27794 28476 27804 28532
rect 27860 28476 28588 28532
rect 28644 28476 29372 28532
rect 29428 28476 29438 28532
rect 29922 28364 29932 28420
rect 29988 28364 74620 28420
rect 74676 28364 74686 28420
rect 0 28196 800 28224
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 79200 28196 80000 28224
rect 0 28140 2156 28196
rect 2212 28140 2222 28196
rect 77746 28140 77756 28196
rect 77812 28140 80000 28196
rect 0 28112 800 28140
rect 79200 28112 80000 28140
rect 28914 27916 28924 27972
rect 28980 27916 76636 27972
rect 76692 27916 76860 27972
rect 76916 27916 76926 27972
rect 27122 27804 27132 27860
rect 27188 27804 27916 27860
rect 27972 27804 28476 27860
rect 28532 27804 29820 27860
rect 29876 27804 29886 27860
rect 3042 27692 3052 27748
rect 3108 27692 3612 27748
rect 3668 27692 27580 27748
rect 27636 27692 27646 27748
rect 0 27524 800 27552
rect 79200 27524 80000 27552
rect 0 27468 2044 27524
rect 2100 27468 2110 27524
rect 76066 27468 76076 27524
rect 76132 27468 80000 27524
rect 0 27440 800 27468
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 79200 27440 80000 27468
rect 3042 27020 3052 27076
rect 3108 27020 3612 27076
rect 3668 27020 26908 27076
rect 26964 27020 26974 27076
rect 26450 26908 26460 26964
rect 26516 26908 27244 26964
rect 27300 26908 28028 26964
rect 28084 26908 28812 26964
rect 28868 26908 28878 26964
rect 0 26852 800 26880
rect 79200 26852 80000 26880
rect 0 26796 2156 26852
rect 2212 26796 2222 26852
rect 28354 26796 28364 26852
rect 28420 26796 74620 26852
rect 74676 26796 74686 26852
rect 77746 26796 77756 26852
rect 77812 26796 80000 26852
rect 0 26768 800 26796
rect 79200 26768 80000 26796
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 27682 26348 27692 26404
rect 27748 26348 76860 26404
rect 76916 26348 77196 26404
rect 77252 26348 77262 26404
rect 0 26180 800 26208
rect 79200 26180 80000 26208
rect 0 26124 2044 26180
rect 2100 26124 2110 26180
rect 4834 26124 4844 26180
rect 4900 26124 5404 26180
rect 5460 26124 24332 26180
rect 24388 26124 24398 26180
rect 25778 26124 25788 26180
rect 25844 26124 26460 26180
rect 26516 26124 26526 26180
rect 76066 26124 76076 26180
rect 76132 26124 80000 26180
rect 0 26096 800 26124
rect 79200 26096 80000 26124
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 0 25508 800 25536
rect 79200 25508 80000 25536
rect 0 25452 3836 25508
rect 3892 25452 3902 25508
rect 25554 25452 25564 25508
rect 25620 25452 26348 25508
rect 26404 25452 27580 25508
rect 27636 25452 27646 25508
rect 77746 25452 77756 25508
rect 77812 25452 80000 25508
rect 0 25424 800 25452
rect 79200 25424 80000 25452
rect 3042 25340 3052 25396
rect 3108 25340 4060 25396
rect 4116 25340 25228 25396
rect 25284 25340 25294 25396
rect 26450 25340 26460 25396
rect 26516 25340 27132 25396
rect 27188 25340 27356 25396
rect 27412 25340 27422 25396
rect 2930 25228 2940 25284
rect 2996 25228 3612 25284
rect 3668 25228 26236 25284
rect 26292 25228 26302 25284
rect 26674 25228 26684 25284
rect 26740 25228 74620 25284
rect 74676 25228 74686 25284
rect 74722 25116 74732 25172
rect 74788 25116 75292 25172
rect 75348 25116 75358 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 0 24836 800 24864
rect 79200 24836 80000 24864
rect 0 24780 2156 24836
rect 2212 24780 2222 24836
rect 26114 24780 26124 24836
rect 26180 24780 55468 24836
rect 76178 24780 76188 24836
rect 76244 24780 80000 24836
rect 0 24752 800 24780
rect 55412 24724 55468 24780
rect 79200 24752 80000 24780
rect 55412 24668 76636 24724
rect 76692 24668 76860 24724
rect 76916 24668 76926 24724
rect 3042 24556 3052 24612
rect 3108 24556 3612 24612
rect 3668 24556 24108 24612
rect 24164 24556 24174 24612
rect 24882 24556 24892 24612
rect 24948 24556 25900 24612
rect 25956 24556 27020 24612
rect 27076 24556 27086 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 0 24164 800 24192
rect 79200 24164 80000 24192
rect 0 24108 2044 24164
rect 2100 24108 2110 24164
rect 76066 24108 76076 24164
rect 76132 24108 80000 24164
rect 0 24080 800 24108
rect 79200 24080 80000 24108
rect 26674 23772 26684 23828
rect 26740 23772 74620 23828
rect 74676 23772 74686 23828
rect 3042 23660 3052 23716
rect 3108 23660 3612 23716
rect 3668 23660 23660 23716
rect 23716 23660 23726 23716
rect 24658 23660 24668 23716
rect 24724 23660 25564 23716
rect 25620 23660 25630 23716
rect 25778 23660 25788 23716
rect 25844 23660 74508 23716
rect 74564 23660 74574 23716
rect 23986 23548 23996 23604
rect 24052 23548 26012 23604
rect 26068 23548 26348 23604
rect 26404 23548 26414 23604
rect 0 23492 800 23520
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 79200 23492 80000 23520
rect 0 23436 2156 23492
rect 2212 23436 2222 23492
rect 77746 23436 77756 23492
rect 77812 23436 80000 23492
rect 0 23408 800 23436
rect 79200 23408 80000 23436
rect 23874 23212 23884 23268
rect 23940 23212 76636 23268
rect 76692 23212 76860 23268
rect 76916 23212 76926 23268
rect 22754 23100 22764 23156
rect 22820 23100 23100 23156
rect 23156 23100 23660 23156
rect 23716 23100 24780 23156
rect 24836 23100 24846 23156
rect 3042 22988 3052 23044
rect 3108 22988 3612 23044
rect 3668 22988 22428 23044
rect 22484 22988 22494 23044
rect 0 22820 800 22848
rect 79200 22820 80000 22848
rect 0 22764 2044 22820
rect 2100 22764 2110 22820
rect 76066 22764 76076 22820
rect 76132 22764 80000 22820
rect 0 22736 800 22764
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 79200 22736 80000 22764
rect 3042 22204 3052 22260
rect 3108 22204 3612 22260
rect 3668 22204 22092 22260
rect 22148 22204 22158 22260
rect 22418 22204 22428 22260
rect 22484 22204 22988 22260
rect 23044 22204 23054 22260
rect 0 22148 800 22176
rect 22428 22148 22484 22204
rect 79200 22148 80000 22176
rect 0 22092 2156 22148
rect 2212 22092 2222 22148
rect 21634 22092 21644 22148
rect 21700 22092 22484 22148
rect 23314 22092 23324 22148
rect 23380 22092 74620 22148
rect 74676 22092 74686 22148
rect 77746 22092 77756 22148
rect 77812 22092 80000 22148
rect 0 22064 800 22092
rect 79200 22064 80000 22092
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 23986 21644 23996 21700
rect 24052 21644 76860 21700
rect 76916 21644 77196 21700
rect 77252 21644 77262 21700
rect 0 21476 800 21504
rect 79200 21476 80000 21504
rect 0 21420 2044 21476
rect 2100 21420 2110 21476
rect 4834 21420 4844 21476
rect 4900 21420 5404 21476
rect 5460 21420 19628 21476
rect 19684 21420 19694 21476
rect 76066 21420 76076 21476
rect 76132 21420 80000 21476
rect 0 21392 800 21420
rect 79200 21392 80000 21420
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 0 20804 800 20832
rect 79200 20804 80000 20832
rect 0 20748 3836 20804
rect 3892 20748 3902 20804
rect 77868 20748 80000 20804
rect 0 20720 800 20748
rect 3042 20636 3052 20692
rect 3108 20636 4060 20692
rect 4116 20636 21644 20692
rect 21700 20636 21710 20692
rect 2930 20524 2940 20580
rect 2996 20524 3612 20580
rect 3668 20524 21532 20580
rect 21588 20524 21598 20580
rect 21858 20524 21868 20580
rect 21924 20524 22428 20580
rect 22484 20524 23100 20580
rect 23156 20524 23166 20580
rect 23538 20524 23548 20580
rect 23604 20524 74508 20580
rect 74564 20524 74574 20580
rect 23100 20468 23156 20524
rect 23100 20412 23660 20468
rect 23716 20412 23726 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 76178 20188 76188 20244
rect 76244 20188 76468 20244
rect 0 20132 800 20160
rect 0 20076 2156 20132
rect 2212 20076 2222 20132
rect 74498 20076 74508 20132
rect 74564 20076 75292 20132
rect 75348 20076 75358 20132
rect 0 20048 800 20076
rect 76412 20020 76468 20188
rect 77868 20132 77924 20748
rect 79200 20720 80000 20748
rect 79200 20132 80000 20160
rect 77746 20076 77756 20132
rect 77812 20076 77924 20132
rect 77980 20076 80000 20132
rect 77980 20020 78036 20076
rect 79200 20048 80000 20076
rect 19506 19964 19516 20020
rect 19572 19964 20300 20020
rect 20356 19964 20636 20020
rect 20692 19964 20860 20020
rect 20916 19964 20926 20020
rect 21186 19964 21196 20020
rect 21252 19964 55468 20020
rect 76412 19964 78036 20020
rect 55412 19908 55468 19964
rect 3042 19852 3052 19908
rect 3108 19852 3612 19908
rect 3668 19852 19404 19908
rect 19460 19852 19470 19908
rect 22194 19852 22204 19908
rect 22260 19852 22876 19908
rect 22932 19852 22942 19908
rect 55412 19852 76636 19908
rect 76692 19852 76860 19908
rect 76916 19852 76926 19908
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 0 19460 800 19488
rect 79200 19460 80000 19488
rect 0 19404 2044 19460
rect 2100 19404 2110 19460
rect 76066 19404 76076 19460
rect 76132 19404 80000 19460
rect 0 19376 800 19404
rect 79200 19376 80000 19404
rect 19842 19068 19852 19124
rect 19908 19068 20524 19124
rect 20580 19068 20590 19124
rect 21970 19068 21980 19124
rect 22036 19068 74620 19124
rect 74676 19068 74686 19124
rect 20738 18956 20748 19012
rect 20804 18956 74508 19012
rect 74564 18956 74574 19012
rect 3042 18844 3052 18900
rect 3108 18844 3612 18900
rect 3668 18844 18620 18900
rect 18676 18844 18686 18900
rect 20514 18844 20524 18900
rect 20580 18844 21756 18900
rect 21812 18844 21980 18900
rect 22036 18844 22046 18900
rect 0 18788 800 18816
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 79200 18788 80000 18816
rect 0 18732 2156 18788
rect 2212 18732 2222 18788
rect 77868 18732 80000 18788
rect 0 18704 800 18732
rect 18162 18620 18172 18676
rect 18228 18620 18956 18676
rect 19012 18620 20860 18676
rect 20916 18620 21532 18676
rect 21588 18620 21598 18676
rect 20066 18508 20076 18564
rect 20132 18508 20412 18564
rect 20468 18508 20478 18564
rect 54786 18508 54796 18564
rect 54852 18508 55580 18564
rect 55636 18508 55646 18564
rect 77868 18452 77924 18732
rect 79200 18704 80000 18732
rect 54562 18396 54572 18452
rect 54628 18396 56028 18452
rect 56084 18396 56094 18452
rect 77746 18396 77756 18452
rect 77812 18396 77924 18452
rect 3042 18284 3052 18340
rect 3108 18284 3612 18340
rect 3668 18284 18620 18340
rect 18676 18284 18686 18340
rect 55010 18284 55020 18340
rect 55076 18284 55804 18340
rect 55860 18284 55870 18340
rect 0 18116 800 18144
rect 79200 18116 80000 18144
rect 0 18060 2044 18116
rect 2100 18060 2110 18116
rect 76066 18060 76076 18116
rect 76132 18060 80000 18116
rect 0 18032 800 18060
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 79200 18032 80000 18060
rect 18946 17836 18956 17892
rect 19012 17836 74620 17892
rect 74676 17836 74686 17892
rect 19618 17724 19628 17780
rect 19684 17724 74508 17780
rect 74564 17724 74574 17780
rect 21074 17612 21084 17668
rect 21140 17612 76636 17668
rect 76692 17612 76702 17668
rect 20290 17500 20300 17556
rect 20356 17500 21532 17556
rect 21588 17500 21598 17556
rect 25442 17500 25452 17556
rect 25508 17500 25788 17556
rect 25844 17500 27020 17556
rect 27076 17500 27086 17556
rect 0 17444 800 17472
rect 79200 17444 80000 17472
rect 0 17388 2156 17444
rect 2212 17388 2222 17444
rect 3042 17388 3052 17444
rect 3108 17388 3612 17444
rect 3668 17388 17724 17444
rect 17780 17388 17790 17444
rect 20066 17388 20076 17444
rect 20132 17388 20636 17444
rect 20692 17388 20702 17444
rect 26002 17388 26012 17444
rect 26068 17388 26236 17444
rect 26292 17388 26572 17444
rect 26628 17388 26638 17444
rect 54002 17388 54012 17444
rect 54068 17388 55468 17444
rect 55524 17388 56028 17444
rect 56084 17388 56588 17444
rect 56644 17388 56654 17444
rect 77746 17388 77756 17444
rect 77812 17388 80000 17444
rect 0 17360 800 17388
rect 79200 17360 80000 17388
rect 23202 17276 23212 17332
rect 23268 17276 31948 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 20850 17164 20860 17220
rect 20916 17164 26012 17220
rect 26068 17164 26078 17220
rect 31892 17108 31948 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 54562 17164 54572 17220
rect 54628 17164 55132 17220
rect 55188 17164 55198 17220
rect 19394 17052 19404 17108
rect 19460 17052 20300 17108
rect 20356 17052 20366 17108
rect 24322 17052 24332 17108
rect 24388 17052 24892 17108
rect 24948 17052 25788 17108
rect 25844 17052 25854 17108
rect 31892 17052 53564 17108
rect 53620 17052 55020 17108
rect 55076 17052 55086 17108
rect 3042 16940 3052 16996
rect 3108 16940 3612 16996
rect 3668 16940 16604 16996
rect 16660 16940 16670 16996
rect 18610 16940 18620 16996
rect 18676 16940 76860 16996
rect 76916 16940 77196 16996
rect 77252 16940 77262 16996
rect 4834 16828 4844 16884
rect 4900 16828 5404 16884
rect 5460 16828 15596 16884
rect 15652 16828 15662 16884
rect 17042 16828 17052 16884
rect 17108 16828 18060 16884
rect 18116 16828 18508 16884
rect 18564 16828 18574 16884
rect 21522 16828 21532 16884
rect 21588 16828 22428 16884
rect 22484 16828 22652 16884
rect 22708 16828 22988 16884
rect 23044 16828 23054 16884
rect 24434 16828 24444 16884
rect 24500 16828 25676 16884
rect 25732 16828 25742 16884
rect 26674 16828 26684 16884
rect 26740 16828 54460 16884
rect 54516 16828 55244 16884
rect 55300 16828 55310 16884
rect 75954 16828 75964 16884
rect 76020 16828 76030 16884
rect 0 16772 800 16800
rect 75964 16772 76020 16828
rect 79200 16772 80000 16800
rect 0 16716 2044 16772
rect 2100 16716 2110 16772
rect 19618 16716 19628 16772
rect 19684 16716 20748 16772
rect 20804 16716 20814 16772
rect 22306 16716 22316 16772
rect 22372 16716 23324 16772
rect 23380 16716 23390 16772
rect 75964 16716 80000 16772
rect 0 16688 800 16716
rect 79200 16688 80000 16716
rect 23090 16604 23100 16660
rect 23156 16604 23884 16660
rect 23940 16604 23950 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 17602 16156 17612 16212
rect 17668 16156 18956 16212
rect 19012 16156 19404 16212
rect 19460 16156 19470 16212
rect 0 16100 800 16128
rect 79200 16100 80000 16128
rect 0 16044 3836 16100
rect 3892 16044 3902 16100
rect 19058 16044 19068 16100
rect 19124 16044 22652 16100
rect 22708 16044 22718 16100
rect 74722 16044 74732 16100
rect 74788 16044 75292 16100
rect 75348 16044 75358 16100
rect 77746 16044 77756 16100
rect 77812 16044 80000 16100
rect 0 16016 800 16044
rect 79200 16016 80000 16044
rect 3042 15820 3052 15876
rect 3108 15820 4060 15876
rect 4116 15820 15820 15876
rect 15876 15820 15886 15876
rect 16034 15820 16044 15876
rect 16100 15820 17276 15876
rect 17332 15820 18732 15876
rect 18788 15820 19292 15876
rect 19348 15820 19628 15876
rect 19684 15820 19694 15876
rect 19954 15820 19964 15876
rect 20020 15820 76860 15876
rect 76916 15820 76926 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 0 15428 800 15456
rect 79200 15428 80000 15456
rect 0 15372 2156 15428
rect 2212 15372 2222 15428
rect 55906 15372 55916 15428
rect 55972 15372 74732 15428
rect 74788 15372 74798 15428
rect 76178 15372 76188 15428
rect 76244 15372 80000 15428
rect 0 15344 800 15372
rect 79200 15344 80000 15372
rect 15474 15260 15484 15316
rect 15540 15260 53900 15316
rect 53956 15260 54796 15316
rect 54852 15260 55020 15316
rect 55076 15260 55580 15316
rect 55636 15260 55646 15316
rect 3042 15148 3052 15204
rect 3108 15148 3612 15204
rect 3668 15148 14700 15204
rect 14756 15148 14766 15204
rect 15922 15148 15932 15204
rect 15988 15148 16380 15204
rect 16436 15148 17724 15204
rect 17780 15148 17790 15204
rect 56130 15148 56140 15204
rect 56196 15148 74620 15204
rect 74676 15148 75068 15204
rect 75124 15148 75134 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 0 14756 800 14784
rect 79200 14756 80000 14784
rect 0 14700 2044 14756
rect 2100 14700 2110 14756
rect 76066 14700 76076 14756
rect 76132 14700 80000 14756
rect 0 14672 800 14700
rect 79200 14672 80000 14700
rect 55412 14476 55916 14532
rect 55972 14476 56588 14532
rect 56644 14476 56654 14532
rect 55412 14420 55468 14476
rect 14354 14364 14364 14420
rect 14420 14364 14812 14420
rect 14868 14364 53452 14420
rect 53508 14364 55020 14420
rect 55076 14364 55468 14420
rect 3042 14252 3052 14308
rect 3108 14252 3612 14308
rect 3668 14252 14028 14308
rect 14084 14252 14094 14308
rect 54572 14252 54796 14308
rect 54852 14252 54862 14308
rect 54572 14196 54628 14252
rect 54562 14140 54572 14196
rect 54628 14140 54638 14196
rect 0 14084 800 14112
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 79200 14084 80000 14112
rect 0 14028 2156 14084
rect 2212 14028 2222 14084
rect 77746 14028 77756 14084
rect 77812 14028 80000 14084
rect 0 14000 800 14028
rect 79200 14000 80000 14028
rect 55570 13804 55580 13860
rect 55636 13804 76636 13860
rect 76692 13804 76860 13860
rect 76916 13804 76926 13860
rect 12002 13692 12012 13748
rect 12068 13692 12796 13748
rect 12852 13692 13916 13748
rect 13972 13692 15148 13748
rect 15092 13636 15148 13692
rect 55412 13636 55468 13748
rect 55524 13692 56700 13748
rect 56756 13692 57484 13748
rect 57540 13692 57550 13748
rect 57810 13692 57820 13748
rect 57876 13692 74620 13748
rect 74676 13692 75068 13748
rect 75124 13692 75134 13748
rect 3042 13580 3052 13636
rect 3108 13580 3612 13636
rect 3668 13580 13356 13636
rect 13412 13580 13422 13636
rect 15092 13580 55468 13636
rect 13682 13468 13692 13524
rect 13748 13468 14140 13524
rect 14196 13468 54348 13524
rect 54404 13468 54908 13524
rect 54964 13468 55244 13524
rect 55300 13468 55310 13524
rect 76066 13468 76076 13524
rect 76132 13468 76142 13524
rect 0 13412 800 13440
rect 76076 13412 76132 13468
rect 79200 13412 80000 13440
rect 0 13356 2044 13412
rect 2100 13356 2110 13412
rect 76076 13356 80000 13412
rect 0 13328 800 13356
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 79200 13328 80000 13356
rect 0 12740 800 12768
rect 79200 12740 80000 12768
rect 0 12684 2156 12740
rect 2212 12684 2222 12740
rect 3042 12684 3052 12740
rect 3108 12684 3612 12740
rect 3668 12684 12460 12740
rect 12516 12684 12526 12740
rect 77746 12684 77756 12740
rect 77812 12684 80000 12740
rect 0 12656 800 12684
rect 79200 12656 80000 12684
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 3042 12236 3052 12292
rect 3108 12236 3612 12292
rect 3668 12236 12236 12292
rect 12292 12236 12302 12292
rect 13570 12236 13580 12292
rect 13636 12236 76860 12292
rect 76916 12236 77196 12292
rect 77252 12236 77262 12292
rect 12674 12124 12684 12180
rect 12740 12124 13020 12180
rect 13076 12124 13244 12180
rect 13300 12124 14028 12180
rect 14084 12124 14094 12180
rect 0 12068 800 12096
rect 79200 12068 80000 12096
rect 0 12012 2044 12068
rect 2100 12012 2110 12068
rect 76066 12012 76076 12068
rect 76132 12012 80000 12068
rect 0 11984 800 12012
rect 79200 11984 80000 12012
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 3042 11452 3052 11508
rect 3108 11452 4060 11508
rect 4116 11452 11340 11508
rect 11396 11452 11406 11508
rect 0 11396 800 11424
rect 79200 11396 80000 11424
rect 0 11340 3836 11396
rect 3892 11340 3902 11396
rect 77746 11340 77756 11396
rect 77812 11340 80000 11396
rect 0 11312 800 11340
rect 79200 11312 80000 11340
rect 4834 11228 4844 11284
rect 4900 11228 10780 11284
rect 10836 11228 10846 11284
rect 12898 11228 12908 11284
rect 12964 11228 74620 11284
rect 74676 11228 74686 11284
rect 12002 11116 12012 11172
rect 12068 11116 76860 11172
rect 76916 11116 76926 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 74722 10780 74732 10836
rect 74788 10780 75292 10836
rect 75348 10780 75358 10836
rect 0 10724 800 10752
rect 74732 10724 74788 10780
rect 79200 10724 80000 10752
rect 0 10668 2156 10724
rect 2212 10668 2222 10724
rect 3042 10668 3052 10724
rect 3108 10668 10108 10724
rect 10164 10668 10174 10724
rect 11442 10668 11452 10724
rect 11508 10668 74788 10724
rect 76178 10668 76188 10724
rect 76244 10668 80000 10724
rect 0 10640 800 10668
rect 79200 10640 80000 10668
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 76066 10108 76076 10164
rect 76132 10108 76142 10164
rect 0 10052 800 10080
rect 76076 10052 76132 10108
rect 79200 10052 80000 10080
rect 0 9996 2044 10052
rect 2100 9996 2110 10052
rect 76076 9996 80000 10052
rect 0 9968 800 9996
rect 79200 9968 80000 9996
rect 3042 9660 3052 9716
rect 3108 9660 9436 9716
rect 9492 9660 9502 9716
rect 9650 9660 9660 9716
rect 9716 9660 10556 9716
rect 10612 9660 10622 9716
rect 11554 9660 11564 9716
rect 11620 9660 11900 9716
rect 11956 9660 11966 9716
rect 10882 9548 10892 9604
rect 10948 9548 74620 9604
rect 74676 9548 74686 9604
rect 0 9380 800 9408
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 79200 9380 80000 9408
rect 0 9324 2156 9380
rect 2212 9324 2222 9380
rect 77746 9324 77756 9380
rect 77812 9324 80000 9380
rect 0 9296 800 9324
rect 79200 9296 80000 9324
rect 15698 9212 15708 9268
rect 15764 9212 16268 9268
rect 16324 9212 16334 9268
rect 3042 9100 3052 9156
rect 3108 9100 8652 9156
rect 8708 9100 8718 9156
rect 10210 9100 10220 9156
rect 10276 9100 76636 9156
rect 76692 9100 76702 9156
rect 8978 8988 8988 9044
rect 9044 8988 9884 9044
rect 9940 8988 9950 9044
rect 0 8708 800 8736
rect 79200 8708 80000 8736
rect 0 8652 2044 8708
rect 2100 8652 2110 8708
rect 76066 8652 76076 8708
rect 76132 8652 80000 8708
rect 0 8624 800 8652
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 79200 8624 80000 8652
rect 3042 8092 3052 8148
rect 3108 8092 7980 8148
rect 8036 8092 8046 8148
rect 8306 8092 8316 8148
rect 8372 8092 9100 8148
rect 9156 8092 9772 8148
rect 9828 8092 9838 8148
rect 0 8036 800 8064
rect 79200 8036 80000 8064
rect 0 7980 2156 8036
rect 2212 7980 2222 8036
rect 9426 7980 9436 8036
rect 9492 7980 74620 8036
rect 74676 7980 74686 8036
rect 77746 7980 77756 8036
rect 77812 7980 80000 8036
rect 0 7952 800 7980
rect 79200 7952 80000 7980
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 3042 7532 3052 7588
rect 3108 7532 7420 7588
rect 7476 7532 7486 7588
rect 8754 7532 8764 7588
rect 8820 7532 76860 7588
rect 76916 7532 77196 7588
rect 77252 7532 77262 7588
rect 7634 7420 7644 7476
rect 7700 7420 8428 7476
rect 8484 7420 8494 7476
rect 0 7364 800 7392
rect 79200 7364 80000 7392
rect 0 7308 2156 7364
rect 2212 7308 2222 7364
rect 76066 7308 76076 7364
rect 76132 7308 80000 7364
rect 0 7280 800 7308
rect 79200 7280 80000 7308
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 3042 6748 3052 6804
rect 3108 6748 6524 6804
rect 6580 6748 6590 6804
rect 0 6692 800 6720
rect 79200 6692 80000 6720
rect 0 6636 3836 6692
rect 3892 6636 3902 6692
rect 6962 6636 6972 6692
rect 7028 6636 7756 6692
rect 7812 6636 7822 6692
rect 57922 6636 57932 6692
rect 57988 6636 60284 6692
rect 60340 6636 60350 6692
rect 63410 6636 63420 6692
rect 63476 6636 66108 6692
rect 66164 6636 66174 6692
rect 66322 6636 66332 6692
rect 66388 6636 67676 6692
rect 67732 6636 67742 6692
rect 74722 6636 74732 6692
rect 74788 6636 75292 6692
rect 75348 6636 75358 6692
rect 77746 6636 77756 6692
rect 77812 6636 80000 6692
rect 0 6608 800 6636
rect 79200 6608 80000 6636
rect 4834 6524 4844 6580
rect 4900 6524 5964 6580
rect 6020 6524 6030 6580
rect 6290 6524 6300 6580
rect 6356 6524 6860 6580
rect 6916 6524 6926 6580
rect 8082 6524 8092 6580
rect 8148 6524 74620 6580
rect 74676 6524 74686 6580
rect 7186 6412 7196 6468
rect 7252 6412 76860 6468
rect 76916 6412 76926 6468
rect 56466 6300 56476 6356
rect 56532 6300 58156 6356
rect 58212 6300 58222 6356
rect 59826 6300 59836 6356
rect 59892 6300 62076 6356
rect 62132 6300 62142 6356
rect 63522 6300 63532 6356
rect 63588 6300 65772 6356
rect 65828 6300 65838 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 54562 6188 54572 6244
rect 54628 6188 57372 6244
rect 57428 6188 57438 6244
rect 59602 6188 59612 6244
rect 59668 6188 61068 6244
rect 61124 6188 61628 6244
rect 61684 6188 61694 6244
rect 62850 6188 62860 6244
rect 62916 6188 64204 6244
rect 64260 6188 64270 6244
rect 65426 6188 65436 6244
rect 65492 6188 66332 6244
rect 66388 6188 66780 6244
rect 66836 6188 66846 6244
rect 68562 6188 68572 6244
rect 68628 6188 69132 6244
rect 69188 6188 69468 6244
rect 69524 6188 69534 6244
rect 52658 6076 52668 6132
rect 52724 6076 54236 6132
rect 54292 6076 54684 6132
rect 54740 6076 54750 6132
rect 54898 6076 54908 6132
rect 54964 6076 56364 6132
rect 56420 6076 56430 6132
rect 57698 6076 57708 6132
rect 57764 6076 59164 6132
rect 59220 6076 59230 6132
rect 60162 6076 60172 6132
rect 60228 6076 60732 6132
rect 60788 6076 60798 6132
rect 63746 6076 63756 6132
rect 63812 6076 65324 6132
rect 65380 6076 65390 6132
rect 66434 6076 66444 6132
rect 66500 6076 67228 6132
rect 67284 6076 67294 6132
rect 68450 6076 68460 6132
rect 68516 6076 69020 6132
rect 69076 6076 69356 6132
rect 69412 6076 69422 6132
rect 0 6020 800 6048
rect 79200 6020 80000 6048
rect 0 5964 2156 6020
rect 2212 5964 2222 6020
rect 3042 5964 3052 6020
rect 3108 5964 5292 6020
rect 5348 5964 5358 6020
rect 6738 5964 6748 6020
rect 6804 5964 74732 6020
rect 74788 5964 74798 6020
rect 76178 5964 76188 6020
rect 76244 5964 80000 6020
rect 0 5936 800 5964
rect 79200 5936 80000 5964
rect 50306 5852 50316 5908
rect 50372 5852 55468 5908
rect 65874 5852 65884 5908
rect 65940 5852 68124 5908
rect 68180 5852 68190 5908
rect 55412 5796 55468 5852
rect 55412 5740 69244 5796
rect 69300 5740 69310 5796
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 69682 5404 69692 5460
rect 69748 5404 74396 5460
rect 74452 5404 74462 5460
rect 0 5348 800 5376
rect 79200 5348 80000 5376
rect 0 5292 2044 5348
rect 2100 5292 2110 5348
rect 52322 5292 52332 5348
rect 52388 5292 53116 5348
rect 53172 5292 53182 5348
rect 76066 5292 76076 5348
rect 76132 5292 80000 5348
rect 0 5264 800 5292
rect 79200 5264 80000 5292
rect 49970 5180 49980 5236
rect 50036 5180 50876 5236
rect 50932 5180 50942 5236
rect 51762 5180 51772 5236
rect 51828 5180 52668 5236
rect 52724 5180 52734 5236
rect 53554 5180 53564 5236
rect 53620 5180 54124 5236
rect 54180 5180 54190 5236
rect 55010 5180 55020 5236
rect 55076 5180 55916 5236
rect 55972 5180 55982 5236
rect 60946 5180 60956 5236
rect 61012 5180 62076 5236
rect 62132 5180 62142 5236
rect 67106 5180 67116 5236
rect 67172 5180 68012 5236
rect 68068 5180 68078 5236
rect 63746 5068 63756 5124
rect 63812 5068 64316 5124
rect 64372 5068 64382 5124
rect 3042 4956 3052 5012
rect 3108 4956 4620 5012
rect 4676 4956 4686 5012
rect 4946 4956 4956 5012
rect 5012 4956 5740 5012
rect 5796 4956 5806 5012
rect 6066 4844 6076 4900
rect 6132 4844 74620 4900
rect 74676 4844 74686 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 70354 4508 70364 4564
rect 70420 4508 71148 4564
rect 71204 4508 71214 4564
rect 73490 4508 73500 4564
rect 73556 4508 74284 4564
rect 74340 4508 74350 4564
rect 67890 4396 67900 4452
rect 67956 4396 71260 4452
rect 71316 4396 71326 4452
rect 6402 4284 6412 4340
rect 6468 4284 7084 4340
rect 7140 4284 7150 4340
rect 8978 4284 8988 4340
rect 9044 4284 9996 4340
rect 10052 4284 10062 4340
rect 15138 4284 15148 4340
rect 15204 4284 15372 4340
rect 15428 4284 15596 4340
rect 15652 4284 15662 4340
rect 17042 4284 17052 4340
rect 17108 4284 17388 4340
rect 17444 4284 17724 4340
rect 17780 4284 17790 4340
rect 19842 4284 19852 4340
rect 19908 4284 20300 4340
rect 20356 4284 20366 4340
rect 21186 4284 21196 4340
rect 21252 4284 21420 4340
rect 21476 4284 21644 4340
rect 21700 4284 21710 4340
rect 23874 4284 23884 4340
rect 23940 4284 24108 4340
rect 24164 4284 24332 4340
rect 24388 4284 24398 4340
rect 25890 4284 25900 4340
rect 25956 4284 26124 4340
rect 26180 4284 26348 4340
rect 26404 4284 26414 4340
rect 30146 4284 30156 4340
rect 30212 4284 30380 4340
rect 30436 4284 30446 4340
rect 31938 4284 31948 4340
rect 32004 4284 32396 4340
rect 32452 4284 32462 4340
rect 38658 4284 38668 4340
rect 38724 4284 38892 4340
rect 38948 4284 39116 4340
rect 39172 4284 39182 4340
rect 40898 4284 40908 4340
rect 40964 4284 41580 4340
rect 41636 4284 41646 4340
rect 46050 4284 46060 4340
rect 46116 4284 46508 4340
rect 46564 4284 46574 4340
rect 54450 4284 54460 4340
rect 54516 4284 55916 4340
rect 55972 4284 56588 4340
rect 56644 4284 56654 4340
rect 62402 4284 62412 4340
rect 62468 4284 63868 4340
rect 63924 4284 64540 4340
rect 64596 4284 64606 4340
rect 69794 4284 69804 4340
rect 69860 4284 70812 4340
rect 70868 4284 70878 4340
rect 71138 4284 71148 4340
rect 71204 4284 72044 4340
rect 72100 4284 72492 4340
rect 72548 4284 72558 4340
rect 73490 4284 73500 4340
rect 73556 4284 74060 4340
rect 74116 4284 74508 4340
rect 74564 4284 74574 4340
rect 47954 4172 47964 4228
rect 48020 4172 48636 4228
rect 48692 4172 48702 4228
rect 48962 4172 48972 4228
rect 49028 4172 50204 4228
rect 50260 4172 50270 4228
rect 53666 4172 53676 4228
rect 53732 4172 55132 4228
rect 55188 4172 55198 4228
rect 57698 4172 57708 4228
rect 57764 4172 59948 4228
rect 60004 4172 60014 4228
rect 61730 4172 61740 4228
rect 61796 4172 63084 4228
rect 63140 4172 63150 4228
rect 63746 4172 63756 4228
rect 63812 4172 66108 4228
rect 66164 4172 66174 4228
rect 67778 4172 67788 4228
rect 67844 4172 69692 4228
rect 69748 4172 69758 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 51650 3724 51660 3780
rect 51716 3724 53788 3780
rect 53844 3724 53854 3780
rect 50978 3612 50988 3668
rect 51044 3612 53452 3668
rect 53508 3612 53518 3668
rect 54338 3612 54348 3668
rect 54404 3612 57372 3668
rect 57428 3612 57438 3668
rect 58370 3612 58380 3668
rect 58436 3612 61292 3668
rect 61348 3612 61358 3668
rect 62514 3612 62524 3668
rect 62580 3612 65212 3668
rect 65268 3612 65278 3668
rect 65436 3612 67004 3668
rect 67060 3612 67070 3668
rect 71250 3612 71260 3668
rect 71316 3612 73164 3668
rect 73220 3612 73230 3668
rect 65436 3556 65492 3612
rect 21634 3500 21644 3556
rect 21700 3500 22092 3556
rect 22148 3500 22428 3556
rect 22484 3500 22494 3556
rect 42914 3500 42924 3556
rect 42980 3500 43596 3556
rect 43652 3500 43662 3556
rect 44258 3500 44268 3556
rect 44324 3500 44940 3556
rect 44996 3500 45006 3556
rect 46946 3500 46956 3556
rect 47012 3500 47964 3556
rect 48020 3500 48030 3556
rect 50306 3500 50316 3556
rect 50372 3500 52108 3556
rect 52164 3500 52174 3556
rect 55682 3500 55692 3556
rect 55748 3500 58156 3556
rect 58212 3500 58222 3556
rect 59714 3500 59724 3556
rect 59780 3500 61852 3556
rect 61908 3500 61918 3556
rect 64418 3500 64428 3556
rect 64484 3500 65492 3556
rect 65762 3500 65772 3556
rect 65828 3500 67900 3556
rect 67956 3500 67966 3556
rect 68562 3500 68572 3556
rect 68628 3500 70588 3556
rect 70644 3500 70654 3556
rect 5058 3388 5068 3444
rect 5124 3388 5964 3444
rect 6020 3388 6030 3444
rect 8530 3388 8540 3444
rect 8596 3388 9324 3444
rect 9380 3388 9390 3444
rect 45042 3388 45052 3444
rect 45108 3388 45612 3444
rect 45668 3388 45678 3444
rect 45938 3388 45948 3444
rect 46004 3388 47068 3444
rect 47124 3388 47134 3444
rect 48290 3388 48300 3444
rect 48356 3388 49196 3444
rect 49252 3388 49262 3444
rect 49634 3388 49644 3444
rect 49700 3388 51548 3444
rect 51604 3388 51614 3444
rect 52322 3388 52332 3444
rect 52388 3388 55244 3444
rect 55300 3388 55310 3444
rect 56354 3388 56364 3444
rect 56420 3388 59388 3444
rect 59444 3388 59454 3444
rect 60386 3388 60396 3444
rect 60452 3388 63308 3444
rect 63364 3388 63374 3444
rect 66434 3388 66444 3444
rect 66500 3388 69356 3444
rect 69412 3388 69422 3444
rect 70466 3388 70476 3444
rect 70532 3388 72716 3444
rect 72772 3388 72782 3444
rect 73826 3388 73836 3444
rect 73892 3388 74956 3444
rect 75012 3388 75022 3444
rect 35074 3276 35084 3332
rect 35140 3276 36092 3332
rect 36148 3276 36158 3332
rect 70690 3276 70700 3332
rect 70756 3276 72380 3332
rect 72436 3276 72446 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 68348 66668 68404 66724
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 68348 65660 68404 65716
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 63420 63196 63476 63252
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 63420 61068 63476 61124
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 51996 49980 52052 50036
rect 51996 49420 52052 49476
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 76076 4768 76892
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 76860 20128 76892
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 76076 35488 76892
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 76860 50848 76892
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 65888 76076 66208 76892
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 68348 66724 68404 66734
rect 68348 65716 68404 66668
rect 68348 65650 68404 65660
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 63420 63252 63476 63262
rect 63420 61124 63476 63196
rect 63420 61058 63476 61068
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 51996 50036 52052 50046
rect 51996 49476 52052 49980
rect 51996 49410 52052 49420
rect 65888 49420 66208 50932
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__I dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 68768 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A1
timestamp 1666464484
transform 1 0 20720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A2
timestamp 1666464484
transform 1 0 20272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A3
timestamp 1666464484
transform 1 0 21504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A4
timestamp 1666464484
transform 1 0 21952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__A1
timestamp 1666464484
transform 1 0 26544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__A2
timestamp 1666464484
transform 1 0 26992 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__A1
timestamp 1666464484
transform 1 0 24416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__A2
timestamp 1666464484
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__A1
timestamp 1666464484
transform 1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__A2
timestamp 1666464484
transform 1 0 17248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__A3
timestamp 1666464484
transform -1 0 17136 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__A4
timestamp 1666464484
transform 1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__A1
timestamp 1666464484
transform 1 0 21840 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__A2
timestamp 1666464484
transform 1 0 22288 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__A3
timestamp 1666464484
transform 1 0 23856 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__A4
timestamp 1666464484
transform -1 0 21616 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__A1
timestamp 1666464484
transform 1 0 53872 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__A2
timestamp 1666464484
transform 1 0 53424 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__A3
timestamp 1666464484
transform 1 0 54320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__A1
timestamp 1666464484
transform 1 0 53984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__A2
timestamp 1666464484
transform 1 0 54432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__A3
timestamp 1666464484
transform 1 0 53536 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__I
timestamp 1666464484
transform 1 0 57120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__I
timestamp 1666464484
transform -1 0 67312 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__I
timestamp 1666464484
transform 1 0 56560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__A2
timestamp 1666464484
transform 1 0 54544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__A3
timestamp 1666464484
transform 1 0 54992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__I
timestamp 1666464484
transform 1 0 57232 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__I
timestamp 1666464484
transform 1 0 66976 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__I
timestamp 1666464484
transform -1 0 70784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__A2
timestamp 1666464484
transform 1 0 68880 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__B1
timestamp 1666464484
transform 1 0 70672 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I
timestamp 1666464484
transform 1 0 68544 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__I
timestamp 1666464484
transform 1 0 69328 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__A2
timestamp 1666464484
transform -1 0 70000 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__B1
timestamp 1666464484
transform -1 0 70784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__I
timestamp 1666464484
transform 1 0 47264 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I
timestamp 1666464484
transform 1 0 55552 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__I
timestamp 1666464484
transform 1 0 56784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__I
timestamp 1666464484
transform 1 0 51296 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1666464484
transform -1 0 51184 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__I
timestamp 1666464484
transform 1 0 48496 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__I
timestamp 1666464484
transform 1 0 50288 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I
timestamp 1666464484
transform 1 0 47040 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__I
timestamp 1666464484
transform 1 0 52752 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__I
timestamp 1666464484
transform -1 0 49280 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__I
timestamp 1666464484
transform -1 0 52416 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__I
timestamp 1666464484
transform 1 0 49280 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__I
timestamp 1666464484
transform 1 0 52080 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__I
timestamp 1666464484
transform -1 0 59920 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__I
timestamp 1666464484
transform 1 0 47488 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__I
timestamp 1666464484
transform -1 0 61488 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__146__I
timestamp 1666464484
transform 1 0 47712 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__I
timestamp 1666464484
transform 1 0 56896 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__I
timestamp 1666464484
transform 1 0 50736 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__I
timestamp 1666464484
transform -1 0 52864 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__I
timestamp 1666464484
transform -1 0 51744 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I
timestamp 1666464484
transform -1 0 54768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__155__I
timestamp 1666464484
transform -1 0 53648 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__I
timestamp 1666464484
transform 1 0 52416 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__I
timestamp 1666464484
transform 1 0 56224 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__I
timestamp 1666464484
transform 1 0 50848 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__I
timestamp 1666464484
transform -1 0 57568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__I
timestamp 1666464484
transform 1 0 52640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__I
timestamp 1666464484
transform 1 0 58688 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__I
timestamp 1666464484
transform -1 0 56336 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__I
timestamp 1666464484
transform 1 0 57680 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__I
timestamp 1666464484
transform -1 0 59808 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__I
timestamp 1666464484
transform 1 0 55552 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I
timestamp 1666464484
transform 1 0 63168 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__I
timestamp 1666464484
transform 1 0 56672 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I
timestamp 1666464484
transform -1 0 60480 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__I
timestamp 1666464484
transform 1 0 57792 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1666464484
transform -1 0 60032 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I
timestamp 1666464484
transform 1 0 59248 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1666464484
transform 1 0 61824 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I
timestamp 1666464484
transform 1 0 58800 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I
timestamp 1666464484
transform -1 0 62160 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I
timestamp 1666464484
transform 1 0 57904 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1666464484
transform -1 0 67312 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__I
timestamp 1666464484
transform 1 0 58016 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I
timestamp 1666464484
transform 1 0 65296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__I
timestamp 1666464484
transform -1 0 59808 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__I
timestamp 1666464484
transform -1 0 62160 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__I
timestamp 1666464484
transform 1 0 61936 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__I
timestamp 1666464484
transform 1 0 63056 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__I
timestamp 1666464484
transform -1 0 62160 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I
timestamp 1666464484
transform -1 0 64288 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__I
timestamp 1666464484
transform 1 0 60256 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__I
timestamp 1666464484
transform 1 0 68768 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__I
timestamp 1666464484
transform 1 0 59808 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I
timestamp 1666464484
transform -1 0 64960 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__I
timestamp 1666464484
transform 1 0 61600 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I
timestamp 1666464484
transform -1 0 64288 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__I
timestamp 1666464484
transform -1 0 60816 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I
timestamp 1666464484
transform 1 0 66080 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__I
timestamp 1666464484
transform 1 0 65184 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__I
timestamp 1666464484
transform -1 0 67088 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__I
timestamp 1666464484
transform 1 0 62272 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__I
timestamp 1666464484
transform 1 0 64848 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__I
timestamp 1666464484
transform -1 0 62048 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__I
timestamp 1666464484
transform 1 0 67536 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__I
timestamp 1666464484
transform 1 0 63840 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__I
timestamp 1666464484
transform 1 0 69328 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__I
timestamp 1666464484
transform -1 0 66752 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__I
timestamp 1666464484
transform -1 0 70112 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__I
timestamp 1666464484
transform -1 0 67424 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__I
timestamp 1666464484
transform 1 0 66752 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__I
timestamp 1666464484
transform 1 0 73696 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__A2
timestamp 1666464484
transform 1 0 74592 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__I
timestamp 1666464484
transform 1 0 74368 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__A2
timestamp 1666464484
transform -1 0 73472 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__A2
timestamp 1666464484
transform -1 0 68768 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__A2
timestamp 1666464484
transform -1 0 70112 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__I
timestamp 1666464484
transform 1 0 12208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__I
timestamp 1666464484
transform -1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__I
timestamp 1666464484
transform 1 0 56672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__I
timestamp 1666464484
transform 1 0 54880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__I
timestamp 1666464484
transform 1 0 56560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__I
timestamp 1666464484
transform 1 0 54992 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__I
timestamp 1666464484
transform 1 0 19264 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__I
timestamp 1666464484
transform 1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__I
timestamp 1666464484
transform 1 0 17696 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__I
timestamp 1666464484
transform 1 0 17136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__I
timestamp 1666464484
transform 1 0 19600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__I
timestamp 1666464484
transform 1 0 21504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__I
timestamp 1666464484
transform -1 0 21840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__I
timestamp 1666464484
transform -1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__I
timestamp 1666464484
transform 1 0 22848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__I
timestamp 1666464484
transform 1 0 23072 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__I
timestamp 1666464484
transform 1 0 22624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__I
timestamp 1666464484
transform 1 0 24752 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__I
timestamp 1666464484
transform 1 0 25984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__I
timestamp 1666464484
transform 1 0 25536 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__I
timestamp 1666464484
transform 1 0 26992 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__I
timestamp 1666464484
transform 1 0 27552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__I
timestamp 1666464484
transform -1 0 12096 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__280__I
timestamp 1666464484
transform 1 0 14000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__I
timestamp 1666464484
transform -1 0 12096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__I
timestamp 1666464484
transform 1 0 14112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__283__I
timestamp 1666464484
transform 1 0 14784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__I
timestamp 1666464484
transform 1 0 15456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__I
timestamp 1666464484
transform 1 0 16240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__I
timestamp 1666464484
transform -1 0 16464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__I
timestamp 1666464484
transform 1 0 16800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__288__I
timestamp 1666464484
transform -1 0 18256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__I
timestamp 1666464484
transform 1 0 19376 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__I
timestamp 1666464484
transform -1 0 18256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__291__I
timestamp 1666464484
transform 1 0 20048 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__I
timestamp 1666464484
transform -1 0 19600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__I
timestamp 1666464484
transform 1 0 22176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__I
timestamp 1666464484
transform 1 0 22400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__I
timestamp 1666464484
transform -1 0 21728 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__I
timestamp 1666464484
transform -1 0 23184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__I
timestamp 1666464484
transform 1 0 24304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__I
timestamp 1666464484
transform 1 0 24640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__I
timestamp 1666464484
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__I
timestamp 1666464484
transform 1 0 26544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__I
timestamp 1666464484
transform 1 0 27104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__I
timestamp 1666464484
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__I
timestamp 1666464484
transform 1 0 29792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__I
timestamp 1666464484
transform 1 0 29344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__I
timestamp 1666464484
transform 1 0 30352 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__I
timestamp 1666464484
transform -1 0 30016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__I
timestamp 1666464484
transform 1 0 31248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__I
timestamp 1666464484
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__I
timestamp 1666464484
transform 1 0 33824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__I
timestamp 1666464484
transform 1 0 33376 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__I
timestamp 1666464484
transform 1 0 34384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__I
timestamp 1666464484
transform 1 0 34832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__I
timestamp 1666464484
transform 1 0 35616 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__314__I
timestamp 1666464484
transform 1 0 36064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__I
timestamp 1666464484
transform 1 0 37408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__I
timestamp 1666464484
transform 1 0 38752 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__I
timestamp 1666464484
transform 1 0 38304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__318__I
timestamp 1666464484
transform 1 0 39424 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__I
timestamp 1666464484
transform 1 0 40656 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__I
timestamp 1666464484
transform -1 0 38416 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__321__I
timestamp 1666464484
transform 1 0 40208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__I
timestamp 1666464484
transform 1 0 42336 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__323__I
timestamp 1666464484
transform 1 0 42784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__I
timestamp 1666464484
transform 1 0 43904 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__I
timestamp 1666464484
transform 1 0 44128 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__I
timestamp 1666464484
transform 1 0 44800 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__I
timestamp 1666464484
transform 1 0 45248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__I
timestamp 1666464484
transform 1 0 46032 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__I
timestamp 1666464484
transform 1 0 47376 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__I
timestamp 1666464484
transform 1 0 48048 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__I
timestamp 1666464484
transform 1 0 48272 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__332__I
timestamp 1666464484
transform 1 0 48944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__I
timestamp 1666464484
transform -1 0 25872 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__I
timestamp 1666464484
transform -1 0 26544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__I
timestamp 1666464484
transform -1 0 27216 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__I
timestamp 1666464484
transform -1 0 27888 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__I
timestamp 1666464484
transform -1 0 28336 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__I
timestamp 1666464484
transform 1 0 30800 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__I
timestamp 1666464484
transform -1 0 30800 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__I
timestamp 1666464484
transform 1 0 32032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__I
timestamp 1666464484
transform -1 0 31248 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__I
timestamp 1666464484
transform -1 0 31808 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__I
timestamp 1666464484
transform -1 0 32592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__I
timestamp 1666464484
transform -1 0 33040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__I
timestamp 1666464484
transform -1 0 33824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__I
timestamp 1666464484
transform -1 0 35392 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__I
timestamp 1666464484
transform 1 0 36736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__I
timestamp 1666464484
transform -1 0 35952 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__I
timestamp 1666464484
transform -1 0 36624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__I
timestamp 1666464484
transform 1 0 38752 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__I
timestamp 1666464484
transform -1 0 37968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__I
timestamp 1666464484
transform -1 0 38976 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__I
timestamp 1666464484
transform -1 0 40096 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__I
timestamp 1666464484
transform 1 0 41328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__I
timestamp 1666464484
transform -1 0 40656 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__I
timestamp 1666464484
transform 1 0 43456 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__I
timestamp 1666464484
transform -1 0 42000 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__I
timestamp 1666464484
transform -1 0 42560 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__I
timestamp 1666464484
transform -1 0 44688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__I
timestamp 1666464484
transform -1 0 44016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__I
timestamp 1666464484
transform 1 0 46928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__I
timestamp 1666464484
transform -1 0 47824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__I
timestamp 1666464484
transform -1 0 46144 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__I
timestamp 1666464484
transform -1 0 47936 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__I
timestamp 1666464484
transform 1 0 71680 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__I
timestamp 1666464484
transform 1 0 72352 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__I
timestamp 1666464484
transform 1 0 72800 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__I
timestamp 1666464484
transform 1 0 75040 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__I
timestamp 1666464484
transform -1 0 69552 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__I
timestamp 1666464484
transform -1 0 70224 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__I
timestamp 1666464484
transform -1 0 70784 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__372__I
timestamp 1666464484
transform -1 0 72576 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__I
timestamp 1666464484
transform -1 0 71232 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__374__I
timestamp 1666464484
transform 1 0 69888 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1666464484
transform -1 0 77392 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1666464484
transform -1 0 3696 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1666464484
transform -1 0 5152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1666464484
transform 1 0 12096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1666464484
transform -1 0 12768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1666464484
transform -1 0 13216 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1666464484
transform 1 0 14224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1666464484
transform -1 0 14784 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1666464484
transform -1 0 15232 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1666464484
transform 1 0 16016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1666464484
transform -1 0 16688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1666464484
transform -1 0 17136 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1666464484
transform 1 0 18144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1666464484
transform -1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1666464484
transform 1 0 18816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1666464484
transform -1 0 19488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1666464484
transform -1 0 19936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1666464484
transform 1 0 20832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1666464484
transform -1 0 21280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1666464484
transform 1 0 22400 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1666464484
transform 1 0 22848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1666464484
transform -1 0 23520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1666464484
transform -1 0 23968 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1666464484
transform 1 0 24752 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1666464484
transform -1 0 6496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1666464484
transform 1 0 25984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1666464484
transform -1 0 25984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1666464484
transform 1 0 7616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1666464484
transform 1 0 8064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1666464484
transform 1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1666464484
transform -1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1666464484
transform 1 0 10304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1666464484
transform -1 0 10752 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1666464484
transform -1 0 11200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1666464484
transform -1 0 75040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1666464484
transform -1 0 77392 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1666464484
transform -1 0 77392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1666464484
transform -1 0 77392 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1666464484
transform -1 0 77392 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1666464484
transform -1 0 77392 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1666464484
transform -1 0 77392 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1666464484
transform -1 0 76720 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1666464484
transform -1 0 76496 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1666464484
transform -1 0 77392 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1666464484
transform -1 0 77392 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1666464484
transform -1 0 77392 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1666464484
transform -1 0 77392 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1666464484
transform -1 0 77392 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1666464484
transform -1 0 77392 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1666464484
transform -1 0 76720 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1666464484
transform -1 0 76496 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1666464484
transform -1 0 77392 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1666464484
transform -1 0 77392 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1666464484
transform -1 0 77392 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1666464484
transform -1 0 77392 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1666464484
transform -1 0 76048 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1666464484
transform -1 0 78288 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1666464484
transform -1 0 77392 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1666464484
transform -1 0 76496 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1666464484
transform -1 0 77392 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1666464484
transform -1 0 77392 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1666464484
transform -1 0 77392 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1666464484
transform -1 0 77392 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1666464484
transform -1 0 77392 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1666464484
transform -1 0 77392 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1666464484
transform -1 0 76720 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1666464484
transform -1 0 76496 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1666464484
transform 1 0 3472 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1666464484
transform 1 0 2576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1666464484
transform 1 0 2576 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1666464484
transform 1 0 2576 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1666464484
transform 1 0 3024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1666464484
transform 1 0 3472 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1666464484
transform 1 0 2576 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1666464484
transform -1 0 2800 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1666464484
transform 1 0 2576 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1666464484
transform 1 0 2576 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1666464484
transform 1 0 2576 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1666464484
transform 1 0 3024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1666464484
transform 1 0 3024 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1666464484
transform 1 0 3472 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1666464484
transform 1 0 2576 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1666464484
transform -1 0 2800 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input84_I
timestamp 1666464484
transform 1 0 2576 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input85_I
timestamp 1666464484
transform 1 0 2576 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input86_I
timestamp 1666464484
transform 1 0 2576 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input87_I
timestamp 1666464484
transform 1 0 3024 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input88_I
timestamp 1666464484
transform 1 0 3472 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input89_I
timestamp 1666464484
transform 1 0 3920 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input90_I
timestamp 1666464484
transform -1 0 2800 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input91_I
timestamp 1666464484
transform -1 0 2800 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input92_I
timestamp 1666464484
transform 1 0 3472 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input93_I
timestamp 1666464484
transform 1 0 2576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input94_I
timestamp 1666464484
transform 1 0 2576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input95_I
timestamp 1666464484
transform 1 0 2576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input96_I
timestamp 1666464484
transform 1 0 3024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input97_I
timestamp 1666464484
transform 1 0 3472 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input98_I
timestamp 1666464484
transform 1 0 2576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input99_I
timestamp 1666464484
transform -1 0 2800 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input100_I
timestamp 1666464484
transform 1 0 27104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input101_I
timestamp 1666464484
transform 1 0 33600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input102_I
timestamp 1666464484
transform -1 0 34272 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input103_I
timestamp 1666464484
transform -1 0 34720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input104_I
timestamp 1666464484
transform 1 0 35616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input105_I
timestamp 1666464484
transform -1 0 36288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input106_I
timestamp 1666464484
transform -1 0 36736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input107_I
timestamp 1666464484
transform 1 0 37744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input108_I
timestamp 1666464484
transform -1 0 38304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input109_I
timestamp 1666464484
transform -1 0 38752 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input110_I
timestamp 1666464484
transform 1 0 39872 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input111_I
timestamp 1666464484
transform 1 0 27552 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input112_I
timestamp 1666464484
transform 1 0 40320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input113_I
timestamp 1666464484
transform -1 0 40992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input114_I
timestamp 1666464484
transform -1 0 41440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input115_I
timestamp 1666464484
transform -1 0 42560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input116_I
timestamp 1666464484
transform -1 0 43008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input117_I
timestamp 1666464484
transform -1 0 43456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input118_I
timestamp 1666464484
transform -1 0 44800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input119_I
timestamp 1666464484
transform -1 0 45696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input120_I
timestamp 1666464484
transform 1 0 47264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input121_I
timestamp 1666464484
transform -1 0 46144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input122_I
timestamp 1666464484
transform -1 0 28224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input123_I
timestamp 1666464484
transform 1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input124_I
timestamp 1666464484
transform -1 0 47712 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input125_I
timestamp 1666464484
transform -1 0 28672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input126_I
timestamp 1666464484
transform 1 0 29904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input127_I
timestamp 1666464484
transform -1 0 30016 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input128_I
timestamp 1666464484
transform 1 0 30800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input129_I
timestamp 1666464484
transform -1 0 31584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input130_I
timestamp 1666464484
transform -1 0 32032 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input131_I
timestamp 1666464484
transform -1 0 32816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input132_I
timestamp 1666464484
transform 1 0 72800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input133_I
timestamp 1666464484
transform 1 0 72464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input134_I
timestamp 1666464484
transform -1 0 71680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input135_I
timestamp 1666464484
transform -1 0 73472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input136_I
timestamp 1666464484
transform -1 0 74144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input137_I
timestamp 1666464484
transform 1 0 71008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output138_I
timestamp 1666464484
transform 1 0 74368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output139_I
timestamp 1666464484
transform -1 0 74704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output140_I
timestamp 1666464484
transform -1 0 74704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output141_I
timestamp 1666464484
transform 1 0 77168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output142_I
timestamp 1666464484
transform -1 0 74704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output143_I
timestamp 1666464484
transform -1 0 76720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output144_I
timestamp 1666464484
transform -1 0 74704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output145_I
timestamp 1666464484
transform 1 0 74704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output146_I
timestamp 1666464484
transform -1 0 76720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output147_I
timestamp 1666464484
transform -1 0 74704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output148_I
timestamp 1666464484
transform 1 0 77168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output149_I
timestamp 1666464484
transform -1 0 74704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output150_I
timestamp 1666464484
transform 1 0 74704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output151_I
timestamp 1666464484
transform -1 0 76720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output152_I
timestamp 1666464484
transform -1 0 74704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output153_I
timestamp 1666464484
transform 1 0 74704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output154_I
timestamp 1666464484
transform -1 0 76720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output155_I
timestamp 1666464484
transform -1 0 74704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output156_I
timestamp 1666464484
transform 1 0 77168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output157_I
timestamp 1666464484
transform -1 0 74704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output158_I
timestamp 1666464484
transform -1 0 76720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output159_I
timestamp 1666464484
transform -1 0 74704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output160_I
timestamp 1666464484
transform 1 0 74704 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output161_I
timestamp 1666464484
transform -1 0 76720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output162_I
timestamp 1666464484
transform -1 0 76720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output163_I
timestamp 1666464484
transform -1 0 74704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output164_I
timestamp 1666464484
transform -1 0 74704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output165_I
timestamp 1666464484
transform 1 0 77168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output166_I
timestamp 1666464484
transform -1 0 74704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output167_I
timestamp 1666464484
transform -1 0 76720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output168_I
timestamp 1666464484
transform -1 0 74704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output169_I
timestamp 1666464484
transform 1 0 74704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output170_I
timestamp 1666464484
transform -1 0 76720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output172_I
timestamp 1666464484
transform -1 0 4144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output173_I
timestamp 1666464484
transform -1 0 3696 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output174_I
timestamp 1666464484
transform -1 0 3696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output175_I
timestamp 1666464484
transform -1 0 3696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output176_I
timestamp 1666464484
transform -1 0 3696 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output177_I
timestamp 1666464484
transform -1 0 3696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output178_I
timestamp 1666464484
transform -1 0 5488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output179_I
timestamp 1666464484
transform -1 0 4144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output180_I
timestamp 1666464484
transform -1 0 3696 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output181_I
timestamp 1666464484
transform -1 0 3696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output183_I
timestamp 1666464484
transform -1 0 3696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output184_I
timestamp 1666464484
transform -1 0 3696 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output185_I
timestamp 1666464484
transform -1 0 3696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output186_I
timestamp 1666464484
transform -1 0 5488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output187_I
timestamp 1666464484
transform -1 0 4144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output188_I
timestamp 1666464484
transform -1 0 3696 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output189_I
timestamp 1666464484
transform -1 0 3696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output190_I
timestamp 1666464484
transform -1 0 3696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output191_I
timestamp 1666464484
transform -1 0 3696 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output192_I
timestamp 1666464484
transform -1 0 3696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output194_I
timestamp 1666464484
transform -1 0 5488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output195_I
timestamp 1666464484
transform -1 0 4144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output204_I
timestamp 1666464484
transform -1 0 4144 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output205_I
timestamp 1666464484
transform 1 0 50288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output206_I
timestamp 1666464484
transform -1 0 55104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output207_I
timestamp 1666464484
transform 1 0 57344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output208_I
timestamp 1666464484
transform 1 0 58128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output209_I
timestamp 1666464484
transform 1 0 58688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output210_I
timestamp 1666464484
transform 1 0 59136 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output211_I
timestamp 1666464484
transform 1 0 60256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output212_I
timestamp 1666464484
transform 1 0 60704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output213_I
timestamp 1666464484
transform 1 0 61600 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output214_I
timestamp 1666464484
transform 1 0 62048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output215_I
timestamp 1666464484
transform 1 0 61152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output216_I
timestamp 1666464484
transform -1 0 49392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output217_I
timestamp 1666464484
transform 1 0 64512 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output218_I
timestamp 1666464484
transform 1 0 64176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output219_I
timestamp 1666464484
transform 1 0 65296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output220_I
timestamp 1666464484
transform 1 0 65744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output221_I
timestamp 1666464484
transform 1 0 66192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output222_I
timestamp 1666464484
transform 1 0 66752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output223_I
timestamp 1666464484
transform 1 0 67648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output224_I
timestamp 1666464484
transform 1 0 68096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output225_I
timestamp 1666464484
transform 1 0 67200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output226_I
timestamp 1666464484
transform 1 0 69440 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output227_I
timestamp 1666464484
transform -1 0 50064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output228_I
timestamp 1666464484
transform 1 0 73136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output229_I
timestamp 1666464484
transform 1 0 68992 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output230_I
timestamp 1666464484
transform -1 0 51184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output231_I
timestamp 1666464484
transform 1 0 51744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output232_I
timestamp 1666464484
transform -1 0 52416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output233_I
timestamp 1666464484
transform 1 0 54208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output234_I
timestamp 1666464484
transform -1 0 52864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output235_I
timestamp 1666464484
transform 1 0 56560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output236_I
timestamp 1666464484
transform 1 0 56336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output237_I
timestamp 1666464484
transform 1 0 77168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output238_I
timestamp 1666464484
transform -1 0 74704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output239_I
timestamp 1666464484
transform 1 0 74704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output240_I
timestamp 1666464484
transform -1 0 76720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output241_I
timestamp 1666464484
transform -1 0 74704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output242_I
timestamp 1666464484
transform 1 0 77168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output243_I
timestamp 1666464484
transform -1 0 74704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output244_I
timestamp 1666464484
transform -1 0 76720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output245_I
timestamp 1666464484
transform -1 0 74704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output246_I
timestamp 1666464484
transform 1 0 74704 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output247_I
timestamp 1666464484
transform -1 0 76720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output248_I
timestamp 1666464484
transform -1 0 74704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output249_I
timestamp 1666464484
transform -1 0 74704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output250_I
timestamp 1666464484
transform 1 0 77168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output251_I
timestamp 1666464484
transform -1 0 74704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output252_I
timestamp 1666464484
transform -1 0 76720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output253_I
timestamp 1666464484
transform -1 0 76496 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output254_I
timestamp 1666464484
transform 1 0 76496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output255_I
timestamp 1666464484
transform -1 0 74704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output256_I
timestamp 1666464484
transform -1 0 76720 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output257_I
timestamp 1666464484
transform 1 0 74704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output258_I
timestamp 1666464484
transform -1 0 74704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output259_I
timestamp 1666464484
transform -1 0 76720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output260_I
timestamp 1666464484
transform -1 0 76720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output261_I
timestamp 1666464484
transform -1 0 74704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output262_I
timestamp 1666464484
transform -1 0 74704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output263_I
timestamp 1666464484
transform 1 0 74704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output264_I
timestamp 1666464484
transform -1 0 76720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output265_I
timestamp 1666464484
transform -1 0 74704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output266_I
timestamp 1666464484
transform 1 0 77168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output267_I
timestamp 1666464484
transform -1 0 74704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output268_I
timestamp 1666464484
transform -1 0 76720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output269_I
timestamp 1666464484
transform -1 0 3696 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output270_I
timestamp 1666464484
transform -1 0 3696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output271_I
timestamp 1666464484
transform -1 0 3696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output272_I
timestamp 1666464484
transform -1 0 5488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output273_I
timestamp 1666464484
transform -1 0 4144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output274_I
timestamp 1666464484
transform -1 0 3696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output275_I
timestamp 1666464484
transform -1 0 3696 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output276_I
timestamp 1666464484
transform -1 0 3696 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output277_I
timestamp 1666464484
transform -1 0 3696 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output278_I
timestamp 1666464484
transform -1 0 3696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output279_I
timestamp 1666464484
transform -1 0 3696 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output280_I
timestamp 1666464484
transform -1 0 3696 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output281_I
timestamp 1666464484
transform -1 0 3696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output282_I
timestamp 1666464484
transform 1 0 3472 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output283_I
timestamp 1666464484
transform -1 0 3696 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output284_I
timestamp 1666464484
transform 1 0 3472 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output285_I
timestamp 1666464484
transform -1 0 3696 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output286_I
timestamp 1666464484
transform 1 0 3472 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output287_I
timestamp 1666464484
transform -1 0 3696 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output288_I
timestamp 1666464484
transform 1 0 3472 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output289_I
timestamp 1666464484
transform -1 0 3696 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output290_I
timestamp 1666464484
transform 1 0 3472 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output291_I
timestamp 1666464484
transform -1 0 3696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output292_I
timestamp 1666464484
transform -1 0 3696 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output293_I
timestamp 1666464484
transform 1 0 3472 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output294_I
timestamp 1666464484
transform -1 0 3696 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output295_I
timestamp 1666464484
transform -1 0 3696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output296_I
timestamp 1666464484
transform -1 0 5488 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output297_I
timestamp 1666464484
transform -1 0 4144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output298_I
timestamp 1666464484
transform -1 0 3696 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output299_I
timestamp 1666464484
transform -1 0 3696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output300_I
timestamp 1666464484
transform -1 0 3696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output305_I
timestamp 1666464484
transform 1 0 3472 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output306_I
timestamp 1666464484
transform -1 0 3696 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output307_I
timestamp 1666464484
transform 1 0 3472 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output308_I
timestamp 1666464484
transform -1 0 3696 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output310_I
timestamp 1666464484
transform 1 0 4368 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output312_I
timestamp 1666464484
transform -1 0 3696 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 3360 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 4256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 4704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37
timestamp 1666464484
transform 1 0 5488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45
timestamp 1666464484
transform 1 0 6384 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53
timestamp 1666464484
transform 1 0 7280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61
timestamp 1666464484
transform 1 0 8176 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1666464484
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72
timestamp 1666464484
transform 1 0 9408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80
timestamp 1666464484
transform 1 0 10304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88
timestamp 1666464484
transform 1 0 11200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96
timestamp 1666464484
transform 1 0 12096 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1666464484
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107
timestamp 1666464484
transform 1 0 13328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115
timestamp 1666464484
transform 1 0 14224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123
timestamp 1666464484
transform 1 0 15120 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131
timestamp 1666464484
transform 1 0 16016 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1666464484
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1666464484
transform 1 0 17248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_150
timestamp 1666464484
transform 1 0 18144 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_158
timestamp 1666464484
transform 1 0 19040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_166
timestamp 1666464484
transform 1 0 19936 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1666464484
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_177
timestamp 1666464484
transform 1 0 21168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_185
timestamp 1666464484
transform 1 0 22064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_193
timestamp 1666464484
transform 1 0 22960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_201
timestamp 1666464484
transform 1 0 23856 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1666464484
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_212
timestamp 1666464484
transform 1 0 25088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_220
timestamp 1666464484
transform 1 0 25984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_228
timestamp 1666464484
transform 1 0 26880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_236
timestamp 1666464484
transform 1 0 27776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1666464484
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_247
timestamp 1666464484
transform 1 0 29008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_255
timestamp 1666464484
transform 1 0 29904 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_263
timestamp 1666464484
transform 1 0 30800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_271
timestamp 1666464484
transform 1 0 31696 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1666464484
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_282
timestamp 1666464484
transform 1 0 32928 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_290
timestamp 1666464484
transform 1 0 33824 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_298
timestamp 1666464484
transform 1 0 34720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_306
timestamp 1666464484
transform 1 0 35616 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1666464484
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_317
timestamp 1666464484
transform 1 0 36848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_325
timestamp 1666464484
transform 1 0 37744 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_333
timestamp 1666464484
transform 1 0 38640 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_341
timestamp 1666464484
transform 1 0 39536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1666464484
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_352
timestamp 1666464484
transform 1 0 40768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_358
timestamp 1666464484
transform 1 0 41440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_366
timestamp 1666464484
transform 1 0 42336 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_374
timestamp 1666464484
transform 1 0 43232 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_382
timestamp 1666464484
transform 1 0 44128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1666464484
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1666464484
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_394
timestamp 1666464484
transform 1 0 45472 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_402
timestamp 1666464484
transform 1 0 46368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_410
timestamp 1666464484
transform 1 0 47264 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_418
timestamp 1666464484
transform 1 0 48160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1666464484
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_437
timestamp 1666464484
transform 1 0 50288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_453
timestamp 1666464484
transform 1 0 52080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1666464484
transform 1 0 52528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_472
timestamp 1666464484
transform 1 0 54208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_488
timestamp 1666464484
transform 1 0 56000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1666464484
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_507
timestamp 1666464484
transform 1 0 58128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_523
timestamp 1666464484
transform 1 0 59920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_527
timestamp 1666464484
transform 1 0 60368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_542
timestamp 1666464484
transform 1 0 62048 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_558
timestamp 1666464484
transform 1 0 63840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_562
timestamp 1666464484
transform 1 0 64288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_577
timestamp 1666464484
transform 1 0 65968 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_593
timestamp 1666464484
transform 1 0 67760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1666464484
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_612
timestamp 1666464484
transform 1 0 69888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_628
timestamp 1666464484
transform 1 0 71680 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_632
timestamp 1666464484
transform 1 0 72128 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_639
timestamp 1666464484
transform 1 0 72912 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_643
timestamp 1666464484
transform 1 0 73360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_647
timestamp 1666464484
transform 1 0 73808 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_662
timestamp 1666464484
transform 1 0 75488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1666464484
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_667
timestamp 1666464484
transform 1 0 76048 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_683
timestamp 1666464484
transform 1 0 77840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_687
timestamp 1666464484
transform 1 0 78288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_2
timestamp 1666464484
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_18
timestamp 1666464484
transform 1 0 3360 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_26
timestamp 1666464484
transform 1 0 4256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_30
timestamp 1666464484
transform 1 0 4704 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_34
timestamp 1666464484
transform 1 0 5152 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_42
timestamp 1666464484
transform 1 0 6048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_46
timestamp 1666464484
transform 1 0 6496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_54
timestamp 1666464484
transform 1 0 7392 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_58
timestamp 1666464484
transform 1 0 7840 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_62
timestamp 1666464484
transform 1 0 8288 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_66
timestamp 1666464484
transform 1 0 8736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1666464484
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1666464484
transform 1 0 9520 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_80
timestamp 1666464484
transform 1 0 10304 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_84
timestamp 1666464484
transform 1 0 10752 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_88
timestamp 1666464484
transform 1 0 11200 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_96
timestamp 1666464484
transform 1 0 12096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_102
timestamp 1666464484
transform 1 0 12768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_106
timestamp 1666464484
transform 1 0 13216 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_114
timestamp 1666464484
transform 1 0 14112 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_120
timestamp 1666464484
transform 1 0 14784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_124
timestamp 1666464484
transform 1 0 15232 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_132
timestamp 1666464484
transform 1 0 16128 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_134
timestamp 1666464484
transform 1 0 16352 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_137
timestamp 1666464484
transform 1 0 16688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1666464484
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1666464484
transform 1 0 17472 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_151
timestamp 1666464484
transform 1 0 18256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_155
timestamp 1666464484
transform 1 0 18704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_158
timestamp 1666464484
transform 1 0 19040 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_162
timestamp 1666464484
transform 1 0 19488 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_166
timestamp 1666464484
transform 1 0 19936 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_174
timestamp 1666464484
transform 1 0 20832 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_178
timestamp 1666464484
transform 1 0 21280 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_186
timestamp 1666464484
transform 1 0 22176 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_190
timestamp 1666464484
transform 1 0 22624 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_194
timestamp 1666464484
transform 1 0 23072 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_198
timestamp 1666464484
transform 1 0 23520 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_202
timestamp 1666464484
transform 1 0 23968 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_210
timestamp 1666464484
transform 1 0 24864 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1666464484
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_215
timestamp 1666464484
transform 1 0 25424 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_217
timestamp 1666464484
transform 1 0 25648 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_220
timestamp 1666464484
transform 1 0 25984 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_228
timestamp 1666464484
transform 1 0 26880 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_232
timestamp 1666464484
transform 1 0 27328 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_236
timestamp 1666464484
transform 1 0 27776 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_240
timestamp 1666464484
transform 1 0 28224 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_244
timestamp 1666464484
transform 1 0 28672 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_252
timestamp 1666464484
transform 1 0 29568 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_256
timestamp 1666464484
transform 1 0 30016 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_264
timestamp 1666464484
transform 1 0 30912 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_270
timestamp 1666464484
transform 1 0 31584 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_274
timestamp 1666464484
transform 1 0 32032 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_282
timestamp 1666464484
transform 1 0 32928 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_286
timestamp 1666464484
transform 1 0 33376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_290
timestamp 1666464484
transform 1 0 33824 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_294
timestamp 1666464484
transform 1 0 34272 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_298
timestamp 1666464484
transform 1 0 34720 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_306
timestamp 1666464484
transform 1 0 35616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_312
timestamp 1666464484
transform 1 0 36288 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_316
timestamp 1666464484
transform 1 0 36736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_324
timestamp 1666464484
transform 1 0 37632 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_330
timestamp 1666464484
transform 1 0 38304 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_334
timestamp 1666464484
transform 1 0 38752 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_342
timestamp 1666464484
transform 1 0 39648 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_346
timestamp 1666464484
transform 1 0 40096 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_350
timestamp 1666464484
transform 1 0 40544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1666464484
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_357
timestamp 1666464484
transform 1 0 41328 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_364
timestamp 1666464484
transform 1 0 42112 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_368
timestamp 1666464484
transform 1 0 42560 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_372
timestamp 1666464484
transform 1 0 43008 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_376
timestamp 1666464484
transform 1 0 43456 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_384
timestamp 1666464484
transform 1 0 44352 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_388
timestamp 1666464484
transform 1 0 44800 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_392
timestamp 1666464484
transform 1 0 45248 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_396
timestamp 1666464484
transform 1 0 45696 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_400
timestamp 1666464484
transform 1 0 46144 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_408
timestamp 1666464484
transform 1 0 47040 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_412
timestamp 1666464484
transform 1 0 47488 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_420
timestamp 1666464484
transform 1 0 48384 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_424
timestamp 1666464484
transform 1 0 48832 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1666464484
transform 1 0 49280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_443
timestamp 1666464484
transform 1 0 50960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_459
timestamp 1666464484
transform 1 0 52752 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_475
timestamp 1666464484
transform 1 0 54544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_491
timestamp 1666464484
transform 1 0 56336 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_495
timestamp 1666464484
transform 1 0 56784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_499
timestamp 1666464484
transform 1 0 57232 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_514
timestamp 1666464484
transform 1 0 58912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_530
timestamp 1666464484
transform 1 0 60704 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_546
timestamp 1666464484
transform 1 0 62496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_562
timestamp 1666464484
transform 1 0 64288 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_566
timestamp 1666464484
transform 1 0 64736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1666464484
transform 1 0 65184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_585
timestamp 1666464484
transform 1 0 66864 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_601
timestamp 1666464484
transform 1 0 68656 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_617
timestamp 1666464484
transform 1 0 70448 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_625
timestamp 1666464484
transform 1 0 71344 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_633
timestamp 1666464484
transform 1 0 72240 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_637
timestamp 1666464484
transform 1 0 72688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1666464484
transform 1 0 73136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_648
timestamp 1666464484
transform 1 0 73920 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_656
timestamp 1666464484
transform 1 0 74816 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_664
timestamp 1666464484
transform 1 0 75712 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_680
timestamp 1666464484
transform 1 0 77504 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1666464484
transform 1 0 1568 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_17
timestamp 1666464484
transform 1 0 3248 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_25
timestamp 1666464484
transform 1 0 4144 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 4368 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1666464484
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1666464484
transform 1 0 5488 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_44 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 6272 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_76
timestamp 1666464484
transform 1 0 9856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_82
timestamp 1666464484
transform 1 0 10528 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_90
timestamp 1666464484
transform 1 0 11424 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_94
timestamp 1666464484
transform 1 0 11872 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_98
timestamp 1666464484
transform 1 0 12320 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_108
timestamp 1666464484
transform 1 0 13440 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_112
timestamp 1666464484
transform 1 0 13888 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_114
timestamp 1666464484
transform 1 0 14112 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_117
timestamp 1666464484
transform 1 0 14448 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_125
timestamp 1666464484
transform 1 0 15344 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_129
timestamp 1666464484
transform 1 0 15792 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_133
timestamp 1666464484
transform 1 0 16240 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_149
timestamp 1666464484
transform 1 0 18032 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_152
timestamp 1666464484
transform 1 0 18368 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_168
timestamp 1666464484
transform 1 0 20160 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_172
timestamp 1666464484
transform 1 0 20608 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1666464484
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_179
timestamp 1666464484
transform 1 0 21392 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_195
timestamp 1666464484
transform 1 0 23184 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_203
timestamp 1666464484
transform 1 0 24080 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_207
timestamp 1666464484
transform 1 0 24528 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_211
timestamp 1666464484
transform 1 0 24976 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_219
timestamp 1666464484
transform 1 0 25872 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_222
timestamp 1666464484
transform 1 0 26208 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_238
timestamp 1666464484
transform 1 0 28000 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_246
timestamp 1666464484
transform 1 0 28896 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_250
timestamp 1666464484
transform 1 0 29344 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_254
timestamp 1666464484
transform 1 0 29792 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_257
timestamp 1666464484
transform 1 0 30128 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_261
timestamp 1666464484
transform 1 0 30576 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_265
timestamp 1666464484
transform 1 0 31024 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_273
timestamp 1666464484
transform 1 0 31920 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_277
timestamp 1666464484
transform 1 0 32368 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_281
timestamp 1666464484
transform 1 0 32816 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_297
timestamp 1666464484
transform 1 0 34608 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_305
timestamp 1666464484
transform 1 0 35504 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_308
timestamp 1666464484
transform 1 0 35840 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_316
timestamp 1666464484
transform 1 0 36736 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1666464484
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_321
timestamp 1666464484
transform 1 0 37296 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_327
timestamp 1666464484
transform 1 0 37968 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_359
timestamp 1666464484
transform 1 0 41552 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_375
timestamp 1666464484
transform 1 0 43344 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_383
timestamp 1666464484
transform 1 0 44240 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_387
timestamp 1666464484
transform 1 0 44688 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1666464484
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_392
timestamp 1666464484
transform 1 0 45248 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_408
timestamp 1666464484
transform 1 0 47040 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_414
timestamp 1666464484
transform 1 0 47712 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_422
timestamp 1666464484
transform 1 0 48608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_426
timestamp 1666464484
transform 1 0 49056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_429
timestamp 1666464484
transform 1 0 49392 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_435
timestamp 1666464484
transform 1 0 50064 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_439
timestamp 1666464484
transform 1 0 50512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_445
timestamp 1666464484
transform 1 0 51184 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_449
timestamp 1666464484
transform 1 0 51632 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_452
timestamp 1666464484
transform 1 0 51968 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_456
timestamp 1666464484
transform 1 0 52416 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1666464484
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_463
timestamp 1666464484
transform 1 0 53200 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_478
timestamp 1666464484
transform 1 0 54880 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_494
timestamp 1666464484
transform 1 0 56672 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_512
timestamp 1666464484
transform 1 0 58688 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_530
timestamp 1666464484
transform 1 0 60704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_534
timestamp 1666464484
transform 1 0 61152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_549
timestamp 1666464484
transform 1 0 62832 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_551
timestamp 1666464484
transform 1 0 63056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_566
timestamp 1666464484
transform 1 0 64736 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_584
timestamp 1666464484
transform 1 0 66752 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_602
timestamp 1666464484
transform 1 0 68768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1666464484
transform 1 0 69104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_620
timestamp 1666464484
transform 1 0 70784 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_624
timestamp 1666464484
transform 1 0 71232 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_628
timestamp 1666464484
transform 1 0 71680 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_636
timestamp 1666464484
transform 1 0 72576 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_640
timestamp 1666464484
transform 1 0 73024 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_644
timestamp 1666464484
transform 1 0 73472 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_650
timestamp 1666464484
transform 1 0 74144 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_654
timestamp 1666464484
transform 1 0 74592 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_658
timestamp 1666464484
transform 1 0 75040 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_666
timestamp 1666464484
transform 1 0 75936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_670
timestamp 1666464484
transform 1 0 76384 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1666464484
transform 1 0 76720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_676
timestamp 1666464484
transform 1 0 77056 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_684
timestamp 1666464484
transform 1 0 77952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1666464484
transform 1 0 1568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_17
timestamp 1666464484
transform 1 0 3248 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_33
timestamp 1666464484
transform 1 0 5040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_40
timestamp 1666464484
transform 1 0 5824 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_50
timestamp 1666464484
transform 1 0 6944 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1666464484
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1666464484
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1666464484
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1666464484
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1666464484
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1666464484
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1666464484
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1666464484
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1666464484
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1666464484
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1666464484
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1666464484
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1666464484
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1666464484
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1666464484
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1666464484
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_428
timestamp 1666464484
transform 1 0 49280 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_460
timestamp 1666464484
transform 1 0 52864 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_468
timestamp 1666464484
transform 1 0 53760 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_474
timestamp 1666464484
transform 1 0 54432 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_480
timestamp 1666464484
transform 1 0 55104 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_488
timestamp 1666464484
transform 1 0 56000 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_490
timestamp 1666464484
transform 1 0 56224 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_493
timestamp 1666464484
transform 1 0 56560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_499
timestamp 1666464484
transform 1 0 57232 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_502
timestamp 1666464484
transform 1 0 57568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_506
timestamp 1666464484
transform 1 0 58016 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_509
timestamp 1666464484
transform 1 0 58352 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_511
timestamp 1666464484
transform 1 0 58576 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_514
timestamp 1666464484
transform 1 0 58912 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_518
timestamp 1666464484
transform 1 0 59360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_528
timestamp 1666464484
transform 1 0 60480 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_532
timestamp 1666464484
transform 1 0 60928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_536
timestamp 1666464484
transform 1 0 61376 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_540
timestamp 1666464484
transform 1 0 61824 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_544
timestamp 1666464484
transform 1 0 62272 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_560
timestamp 1666464484
transform 1 0 64064 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_563
timestamp 1666464484
transform 1 0 64400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1666464484
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_570
timestamp 1666464484
transform 1 0 65184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_573
timestamp 1666464484
transform 1 0 65520 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_577
timestamp 1666464484
transform 1 0 65968 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_581
timestamp 1666464484
transform 1 0 66416 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_583
timestamp 1666464484
transform 1 0 66640 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_586
timestamp 1666464484
transform 1 0 66976 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_590
timestamp 1666464484
transform 1 0 67424 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_594
timestamp 1666464484
transform 1 0 67872 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_598
timestamp 1666464484
transform 1 0 68320 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_602
timestamp 1666464484
transform 1 0 68768 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_606
timestamp 1666464484
transform 1 0 69216 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_610
timestamp 1666464484
transform 1 0 69664 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_626
timestamp 1666464484
transform 1 0 71456 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_634
timestamp 1666464484
transform 1 0 72352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1666464484
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_641
timestamp 1666464484
transform 1 0 73136 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_649
timestamp 1666464484
transform 1 0 74032 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_655
timestamp 1666464484
transform 1 0 74704 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_671
timestamp 1666464484
transform 1 0 76496 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_687
timestamp 1666464484
transform 1 0 78288 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_2
timestamp 1666464484
transform 1 0 1568 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_17
timestamp 1666464484
transform 1 0 3248 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_33
timestamp 1666464484
transform 1 0 5040 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_37
timestamp 1666464484
transform 1 0 5488 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_39
timestamp 1666464484
transform 1 0 5712 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_46
timestamp 1666464484
transform 1 0 6496 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_54
timestamp 1666464484
transform 1 0 7392 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_62
timestamp 1666464484
transform 1 0 8288 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_94
timestamp 1666464484
transform 1 0 11872 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_102
timestamp 1666464484
transform 1 0 12768 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1666464484
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1666464484
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1666464484
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1666464484
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1666464484
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1666464484
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1666464484
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1666464484
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1666464484
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1666464484
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1666464484
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1666464484
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1666464484
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1666464484
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1666464484
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_463
timestamp 1666464484
transform 1 0 53200 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1666464484
transform 1 0 60368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1666464484
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_534
timestamp 1666464484
transform 1 0 61152 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_598
timestamp 1666464484
transform 1 0 68320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1666464484
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_605
timestamp 1666464484
transform 1 0 69104 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_637
timestamp 1666464484
transform 1 0 72688 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_653
timestamp 1666464484
transform 1 0 74480 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_657
timestamp 1666464484
transform 1 0 74928 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1666464484
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_676
timestamp 1666464484
transform 1 0 77056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_679
timestamp 1666464484
transform 1 0 77392 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_687
timestamp 1666464484
transform 1 0 78288 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1666464484
transform 1 0 1568 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_17
timestamp 1666464484
transform 1 0 3248 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_33
timestamp 1666464484
transform 1 0 5040 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_41
timestamp 1666464484
transform 1 0 5936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_51
timestamp 1666464484
transform 1 0 7056 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_59
timestamp 1666464484
transform 1 0 7952 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_61
timestamp 1666464484
transform 1 0 8176 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_68
timestamp 1666464484
transform 1 0 8960 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1666464484
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1666464484
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1666464484
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1666464484
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1666464484
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1666464484
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1666464484
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1666464484
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1666464484
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1666464484
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1666464484
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1666464484
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1666464484
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1666464484
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1666464484
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1666464484
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1666464484
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1666464484
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1666464484
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_499
timestamp 1666464484
transform 1 0 57232 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_563
timestamp 1666464484
transform 1 0 64400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1666464484
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_570
timestamp 1666464484
transform 1 0 65184 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_634
timestamp 1666464484
transform 1 0 72352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1666464484
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_641
timestamp 1666464484
transform 1 0 73136 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_649
timestamp 1666464484
transform 1 0 74032 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_655
timestamp 1666464484
transform 1 0 74704 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_671
timestamp 1666464484
transform 1 0 76496 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_687
timestamp 1666464484
transform 1 0 78288 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1666464484
transform 1 0 1568 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_17
timestamp 1666464484
transform 1 0 3248 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_33
timestamp 1666464484
transform 1 0 5040 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1666464484
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_53
timestamp 1666464484
transform 1 0 7280 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_57
timestamp 1666464484
transform 1 0 7728 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_64
timestamp 1666464484
transform 1 0 8512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_74
timestamp 1666464484
transform 1 0 9632 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1666464484
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1666464484
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1666464484
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1666464484
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1666464484
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1666464484
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1666464484
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1666464484
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1666464484
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1666464484
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1666464484
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1666464484
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1666464484
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1666464484
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1666464484
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1666464484
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1666464484
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_534
timestamp 1666464484
transform 1 0 61152 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_598
timestamp 1666464484
transform 1 0 68320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1666464484
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1666464484
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_669
timestamp 1666464484
transform 1 0 76272 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1666464484
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_676
timestamp 1666464484
transform 1 0 77056 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_684
timestamp 1666464484
transform 1 0 77952 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1666464484
transform 1 0 1568 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_17
timestamp 1666464484
transform 1 0 3248 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_49
timestamp 1666464484
transform 1 0 6832 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_57
timestamp 1666464484
transform 1 0 7728 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_61
timestamp 1666464484
transform 1 0 8176 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_63
timestamp 1666464484
transform 1 0 8400 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1666464484
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_73
timestamp 1666464484
transform 1 0 9520 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_81
timestamp 1666464484
transform 1 0 10416 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_113
timestamp 1666464484
transform 1 0 14000 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_129
timestamp 1666464484
transform 1 0 15792 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1666464484
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1666464484
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1666464484
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1666464484
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1666464484
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1666464484
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1666464484
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1666464484
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1666464484
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1666464484
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1666464484
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1666464484
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1666464484
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1666464484
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1666464484
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1666464484
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1666464484
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_499
timestamp 1666464484
transform 1 0 57232 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_563
timestamp 1666464484
transform 1 0 64400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1666464484
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_570
timestamp 1666464484
transform 1 0 65184 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_634
timestamp 1666464484
transform 1 0 72352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1666464484
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_641
timestamp 1666464484
transform 1 0 73136 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_649
timestamp 1666464484
transform 1 0 74032 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_655
timestamp 1666464484
transform 1 0 74704 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_671
timestamp 1666464484
transform 1 0 76496 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_687
timestamp 1666464484
transform 1 0 78288 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_2
timestamp 1666464484
transform 1 0 1568 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_17
timestamp 1666464484
transform 1 0 3248 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_33
timestamp 1666464484
transform 1 0 5040 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_37
timestamp 1666464484
transform 1 0 5488 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_69
timestamp 1666464484
transform 1 0 9072 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_77
timestamp 1666464484
transform 1 0 9968 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_87
timestamp 1666464484
transform 1 0 11088 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_103
timestamp 1666464484
transform 1 0 12880 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1666464484
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1666464484
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1666464484
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1666464484
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1666464484
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1666464484
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1666464484
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1666464484
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1666464484
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1666464484
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1666464484
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1666464484
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1666464484
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1666464484
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1666464484
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1666464484
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1666464484
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1666464484
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1666464484
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1666464484
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_598
timestamp 1666464484
transform 1 0 68320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1666464484
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1666464484
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_669
timestamp 1666464484
transform 1 0 76272 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1666464484
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_676
timestamp 1666464484
transform 1 0 77056 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_684
timestamp 1666464484
transform 1 0 77952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_2
timestamp 1666464484
transform 1 0 1568 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_17
timestamp 1666464484
transform 1 0 3248 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_49
timestamp 1666464484
transform 1 0 6832 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_65
timestamp 1666464484
transform 1 0 8624 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_69
timestamp 1666464484
transform 1 0 9072 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_73
timestamp 1666464484
transform 1 0 9520 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_83
timestamp 1666464484
transform 1 0 10640 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_85
timestamp 1666464484
transform 1 0 10864 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_92
timestamp 1666464484
transform 1 0 11648 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_96
timestamp 1666464484
transform 1 0 12096 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_99
timestamp 1666464484
transform 1 0 12432 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_131
timestamp 1666464484
transform 1 0 16016 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_139
timestamp 1666464484
transform 1 0 16912 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1666464484
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1666464484
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1666464484
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1666464484
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1666464484
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1666464484
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1666464484
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1666464484
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1666464484
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1666464484
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1666464484
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1666464484
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1666464484
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1666464484
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1666464484
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1666464484
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1666464484
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_563
timestamp 1666464484
transform 1 0 64400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1666464484
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1666464484
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1666464484
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1666464484
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_641
timestamp 1666464484
transform 1 0 73136 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_649
timestamp 1666464484
transform 1 0 74032 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_655
timestamp 1666464484
transform 1 0 74704 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_671
timestamp 1666464484
transform 1 0 76496 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_687
timestamp 1666464484
transform 1 0 78288 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_2
timestamp 1666464484
transform 1 0 1568 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_17
timestamp 1666464484
transform 1 0 3248 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_21
timestamp 1666464484
transform 1 0 3696 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_25
timestamp 1666464484
transform 1 0 4144 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_33
timestamp 1666464484
transform 1 0 5040 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_37
timestamp 1666464484
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_69
timestamp 1666464484
transform 1 0 9072 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_77
timestamp 1666464484
transform 1 0 9968 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_81
timestamp 1666464484
transform 1 0 10416 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_89
timestamp 1666464484
transform 1 0 11312 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_97
timestamp 1666464484
transform 1 0 12208 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1666464484
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1666464484
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1666464484
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1666464484
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1666464484
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1666464484
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1666464484
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1666464484
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1666464484
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1666464484
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1666464484
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1666464484
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1666464484
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1666464484
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1666464484
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1666464484
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1666464484
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1666464484
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1666464484
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1666464484
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_598
timestamp 1666464484
transform 1 0 68320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1666464484
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_605
timestamp 1666464484
transform 1 0 69104 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_637
timestamp 1666464484
transform 1 0 72688 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_653
timestamp 1666464484
transform 1 0 74480 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_657
timestamp 1666464484
transform 1 0 74928 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1666464484
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_676
timestamp 1666464484
transform 1 0 77056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_679
timestamp 1666464484
transform 1 0 77392 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_687
timestamp 1666464484
transform 1 0 78288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1666464484
transform 1 0 1568 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_17
timestamp 1666464484
transform 1 0 3248 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_33
timestamp 1666464484
transform 1 0 5040 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_65
timestamp 1666464484
transform 1 0 8624 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_69
timestamp 1666464484
transform 1 0 9072 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_73
timestamp 1666464484
transform 1 0 9520 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_81
timestamp 1666464484
transform 1 0 10416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_85
timestamp 1666464484
transform 1 0 10864 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_87
timestamp 1666464484
transform 1 0 11088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_94
timestamp 1666464484
transform 1 0 11872 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_102
timestamp 1666464484
transform 1 0 12768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_104
timestamp 1666464484
transform 1 0 12992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_111
timestamp 1666464484
transform 1 0 13776 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_115
timestamp 1666464484
transform 1 0 14224 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_131
timestamp 1666464484
transform 1 0 16016 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_139
timestamp 1666464484
transform 1 0 16912 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1666464484
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1666464484
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1666464484
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1666464484
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1666464484
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1666464484
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1666464484
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1666464484
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1666464484
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1666464484
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1666464484
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1666464484
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1666464484
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1666464484
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1666464484
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1666464484
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1666464484
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_563
timestamp 1666464484
transform 1 0 64400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1666464484
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1666464484
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1666464484
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1666464484
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_641
timestamp 1666464484
transform 1 0 73136 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_649
timestamp 1666464484
transform 1 0 74032 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_655
timestamp 1666464484
transform 1 0 74704 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_671
timestamp 1666464484
transform 1 0 76496 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_687
timestamp 1666464484
transform 1 0 78288 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_2
timestamp 1666464484
transform 1 0 1568 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_17
timestamp 1666464484
transform 1 0 3248 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_21
timestamp 1666464484
transform 1 0 3696 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_29
timestamp 1666464484
transform 1 0 4592 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_33
timestamp 1666464484
transform 1 0 5040 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_37
timestamp 1666464484
transform 1 0 5488 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_69
timestamp 1666464484
transform 1 0 9072 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_85
timestamp 1666464484
transform 1 0 10864 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_93
timestamp 1666464484
transform 1 0 11760 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_96
timestamp 1666464484
transform 1 0 12096 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_100
timestamp 1666464484
transform 1 0 12544 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_102
timestamp 1666464484
transform 1 0 12768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1666464484
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1666464484
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1666464484
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1666464484
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1666464484
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1666464484
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1666464484
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1666464484
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1666464484
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1666464484
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1666464484
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1666464484
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1666464484
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1666464484
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1666464484
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1666464484
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_463
timestamp 1666464484
transform 1 0 53200 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_471
timestamp 1666464484
transform 1 0 54096 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_475
timestamp 1666464484
transform 1 0 54544 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_477
timestamp 1666464484
transform 1 0 54768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_480
timestamp 1666464484
transform 1 0 55104 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_512
timestamp 1666464484
transform 1 0 58688 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_528
timestamp 1666464484
transform 1 0 60480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1666464484
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_598
timestamp 1666464484
transform 1 0 68320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1666464484
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1666464484
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_669
timestamp 1666464484
transform 1 0 76272 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1666464484
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_676
timestamp 1666464484
transform 1 0 77056 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_684
timestamp 1666464484
transform 1 0 77952 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_2
timestamp 1666464484
transform 1 0 1568 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_17
timestamp 1666464484
transform 1 0 3248 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_21
timestamp 1666464484
transform 1 0 3696 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_53
timestamp 1666464484
transform 1 0 7280 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_69
timestamp 1666464484
transform 1 0 9072 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_73
timestamp 1666464484
transform 1 0 9520 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_89
timestamp 1666464484
transform 1 0 11312 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_93
timestamp 1666464484
transform 1 0 11760 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_96
timestamp 1666464484
transform 1 0 12096 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_104
timestamp 1666464484
transform 1 0 12992 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_112
timestamp 1666464484
transform 1 0 13888 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_116
timestamp 1666464484
transform 1 0 14336 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_132
timestamp 1666464484
transform 1 0 16128 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_140
timestamp 1666464484
transform 1 0 17024 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1666464484
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1666464484
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1666464484
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1666464484
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1666464484
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1666464484
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1666464484
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1666464484
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1666464484
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1666464484
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1666464484
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1666464484
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_428
timestamp 1666464484
transform 1 0 49280 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_460
timestamp 1666464484
transform 1 0 52864 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_468
timestamp 1666464484
transform 1 0 53760 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_472
timestamp 1666464484
transform 1 0 54208 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_475
timestamp 1666464484
transform 1 0 54544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_479
timestamp 1666464484
transform 1 0 54992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_486
timestamp 1666464484
transform 1 0 55776 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1666464484
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_499
timestamp 1666464484
transform 1 0 57232 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_506
timestamp 1666464484
transform 1 0 58016 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_538
timestamp 1666464484
transform 1 0 61600 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_554
timestamp 1666464484
transform 1 0 63392 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_562
timestamp 1666464484
transform 1 0 64288 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_566
timestamp 1666464484
transform 1 0 64736 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1666464484
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1666464484
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1666464484
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_641
timestamp 1666464484
transform 1 0 73136 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_649
timestamp 1666464484
transform 1 0 74032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_655
timestamp 1666464484
transform 1 0 74704 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_671
timestamp 1666464484
transform 1 0 76496 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_687
timestamp 1666464484
transform 1 0 78288 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_2
timestamp 1666464484
transform 1 0 1568 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_17
timestamp 1666464484
transform 1 0 3248 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_21
timestamp 1666464484
transform 1 0 3696 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_29
timestamp 1666464484
transform 1 0 4592 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_33
timestamp 1666464484
transform 1 0 5040 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1666464484
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1666464484
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1666464484
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_108
timestamp 1666464484
transform 1 0 13440 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_118
timestamp 1666464484
transform 1 0 14560 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_122
timestamp 1666464484
transform 1 0 15008 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_154
timestamp 1666464484
transform 1 0 18592 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_170
timestamp 1666464484
transform 1 0 20384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_174
timestamp 1666464484
transform 1 0 20832 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1666464484
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1666464484
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1666464484
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1666464484
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1666464484
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1666464484
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1666464484
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1666464484
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1666464484
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1666464484
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1666464484
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1666464484
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1666464484
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_463
timestamp 1666464484
transform 1 0 53200 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_467
timestamp 1666464484
transform 1 0 53648 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_471
timestamp 1666464484
transform 1 0 54096 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_483
timestamp 1666464484
transform 1 0 55440 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_491
timestamp 1666464484
transform 1 0 56336 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_495
timestamp 1666464484
transform 1 0 56784 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1666464484
transform 1 0 60368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1666464484
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1666464484
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1666464484
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1666464484
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1666464484
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_669
timestamp 1666464484
transform 1 0 76272 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1666464484
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_676
timestamp 1666464484
transform 1 0 77056 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_684
timestamp 1666464484
transform 1 0 77952 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_2
timestamp 1666464484
transform 1 0 1568 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_17
timestamp 1666464484
transform 1 0 3248 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_21
timestamp 1666464484
transform 1 0 3696 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_53
timestamp 1666464484
transform 1 0 7280 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_69
timestamp 1666464484
transform 1 0 9072 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_73
timestamp 1666464484
transform 1 0 9520 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_105
timestamp 1666464484
transform 1 0 13104 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_113
timestamp 1666464484
transform 1 0 14000 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_117
timestamp 1666464484
transform 1 0 14448 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_124
timestamp 1666464484
transform 1 0 15232 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_128
timestamp 1666464484
transform 1 0 15680 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_132
timestamp 1666464484
transform 1 0 16128 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_135
timestamp 1666464484
transform 1 0 16464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1666464484
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_144
timestamp 1666464484
transform 1 0 17472 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_148
timestamp 1666464484
transform 1 0 17920 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_152
timestamp 1666464484
transform 1 0 18368 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_162
timestamp 1666464484
transform 1 0 19488 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_194
timestamp 1666464484
transform 1 0 23072 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_210
timestamp 1666464484
transform 1 0 24864 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1666464484
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1666464484
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1666464484
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1666464484
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1666464484
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1666464484
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1666464484
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1666464484
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1666464484
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1666464484
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_428
timestamp 1666464484
transform 1 0 49280 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_460
timestamp 1666464484
transform 1 0 52864 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_476
timestamp 1666464484
transform 1 0 54656 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_478
timestamp 1666464484
transform 1 0 54880 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_481
timestamp 1666464484
transform 1 0 55216 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_489
timestamp 1666464484
transform 1 0 56112 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1666464484
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1666464484
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1666464484
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1666464484
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1666464484
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1666464484
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_641
timestamp 1666464484
transform 1 0 73136 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_649
timestamp 1666464484
transform 1 0 74032 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_655
timestamp 1666464484
transform 1 0 74704 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_671
timestamp 1666464484
transform 1 0 76496 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_687
timestamp 1666464484
transform 1 0 78288 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1666464484
transform 1 0 1568 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_17
timestamp 1666464484
transform 1 0 3248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_21
timestamp 1666464484
transform 1 0 3696 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_25
timestamp 1666464484
transform 1 0 4144 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_33
timestamp 1666464484
transform 1 0 5040 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1666464484
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1666464484
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1666464484
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_108
timestamp 1666464484
transform 1 0 13440 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_124
timestamp 1666464484
transform 1 0 15232 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_126
timestamp 1666464484
transform 1 0 15456 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_133
timestamp 1666464484
transform 1 0 16240 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_137
timestamp 1666464484
transform 1 0 16688 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_140
timestamp 1666464484
transform 1 0 17024 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_144
timestamp 1666464484
transform 1 0 17472 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_148
timestamp 1666464484
transform 1 0 17920 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_160
timestamp 1666464484
transform 1 0 19264 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_168
timestamp 1666464484
transform 1 0 20160 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1666464484
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_179
timestamp 1666464484
transform 1 0 21392 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_187
timestamp 1666464484
transform 1 0 22288 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_197
timestamp 1666464484
transform 1 0 23408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_203
timestamp 1666464484
transform 1 0 24080 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_235
timestamp 1666464484
transform 1 0 27664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1666464484
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1666464484
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1666464484
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1666464484
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1666464484
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1666464484
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1666464484
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1666464484
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1666464484
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1666464484
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1666464484
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1666464484
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1666464484
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1666464484
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1666464484
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_598
timestamp 1666464484
transform 1 0 68320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1666464484
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_605
timestamp 1666464484
transform 1 0 69104 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_637
timestamp 1666464484
transform 1 0 72688 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_653
timestamp 1666464484
transform 1 0 74480 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_657
timestamp 1666464484
transform 1 0 74928 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_673
timestamp 1666464484
transform 1 0 76720 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_676
timestamp 1666464484
transform 1 0 77056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_679
timestamp 1666464484
transform 1 0 77392 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_687
timestamp 1666464484
transform 1 0 78288 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_2
timestamp 1666464484
transform 1 0 1568 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_17
timestamp 1666464484
transform 1 0 3248 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_33
timestamp 1666464484
transform 1 0 5040 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_37
timestamp 1666464484
transform 1 0 5488 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_69
timestamp 1666464484
transform 1 0 9072 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_73
timestamp 1666464484
transform 1 0 9520 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_105
timestamp 1666464484
transform 1 0 13104 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_121
timestamp 1666464484
transform 1 0 14896 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_125
timestamp 1666464484
transform 1 0 15344 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_133
timestamp 1666464484
transform 1 0 16240 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1666464484
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_144
timestamp 1666464484
transform 1 0 17472 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_148
timestamp 1666464484
transform 1 0 17920 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_156
timestamp 1666464484
transform 1 0 18816 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_160
timestamp 1666464484
transform 1 0 19264 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_167
timestamp 1666464484
transform 1 0 20048 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_171
timestamp 1666464484
transform 1 0 20496 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_175
timestamp 1666464484
transform 1 0 20944 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_181
timestamp 1666464484
transform 1 0 21616 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_185
timestamp 1666464484
transform 1 0 22064 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_189
timestamp 1666464484
transform 1 0 22512 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_201
timestamp 1666464484
transform 1 0 23856 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_205
timestamp 1666464484
transform 1 0 24304 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_208
timestamp 1666464484
transform 1 0 24640 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1666464484
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_215
timestamp 1666464484
transform 1 0 25424 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_227
timestamp 1666464484
transform 1 0 26768 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_259
timestamp 1666464484
transform 1 0 30352 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_275
timestamp 1666464484
transform 1 0 32144 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1666464484
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1666464484
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1666464484
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1666464484
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1666464484
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1666464484
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1666464484
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_428
timestamp 1666464484
transform 1 0 49280 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_460
timestamp 1666464484
transform 1 0 52864 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_468
timestamp 1666464484
transform 1 0 53760 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_472
timestamp 1666464484
transform 1 0 54208 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_476
timestamp 1666464484
transform 1 0 54656 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1666464484
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1666464484
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1666464484
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_563
timestamp 1666464484
transform 1 0 64400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1666464484
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1666464484
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_634
timestamp 1666464484
transform 1 0 72352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1666464484
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_641
timestamp 1666464484
transform 1 0 73136 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_649
timestamp 1666464484
transform 1 0 74032 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_655
timestamp 1666464484
transform 1 0 74704 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_671
timestamp 1666464484
transform 1 0 76496 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_687
timestamp 1666464484
transform 1 0 78288 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_2
timestamp 1666464484
transform 1 0 1568 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_17
timestamp 1666464484
transform 1 0 3248 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_21
timestamp 1666464484
transform 1 0 3696 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_29
timestamp 1666464484
transform 1 0 4592 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_33
timestamp 1666464484
transform 1 0 5040 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1666464484
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1666464484
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1666464484
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_108
timestamp 1666464484
transform 1 0 13440 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_124
timestamp 1666464484
transform 1 0 15232 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_132
timestamp 1666464484
transform 1 0 16128 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_135
timestamp 1666464484
transform 1 0 16464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_139
timestamp 1666464484
transform 1 0 16912 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_143
timestamp 1666464484
transform 1 0 17360 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_151
timestamp 1666464484
transform 1 0 18256 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_159
timestamp 1666464484
transform 1 0 19152 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_163
timestamp 1666464484
transform 1 0 19600 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_165
timestamp 1666464484
transform 1 0 19824 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1666464484
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_179
timestamp 1666464484
transform 1 0 21392 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_182
timestamp 1666464484
transform 1 0 21728 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_186
timestamp 1666464484
transform 1 0 22176 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_202
timestamp 1666464484
transform 1 0 23968 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_210
timestamp 1666464484
transform 1 0 24864 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_214
timestamp 1666464484
transform 1 0 25312 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_216
timestamp 1666464484
transform 1 0 25536 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_223
timestamp 1666464484
transform 1 0 26320 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_227
timestamp 1666464484
transform 1 0 26768 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_231
timestamp 1666464484
transform 1 0 27216 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1666464484
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1666464484
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1666464484
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1666464484
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1666464484
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1666464484
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1666464484
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1666464484
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1666464484
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1666464484
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_463
timestamp 1666464484
transform 1 0 53200 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_465
timestamp 1666464484
transform 1 0 53424 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_468
timestamp 1666464484
transform 1 0 53760 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_472
timestamp 1666464484
transform 1 0 54208 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_485
timestamp 1666464484
transform 1 0 55664 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_491
timestamp 1666464484
transform 1 0 56336 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_495
timestamp 1666464484
transform 1 0 56784 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_527
timestamp 1666464484
transform 1 0 60368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1666464484
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1666464484
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_598
timestamp 1666464484
transform 1 0 68320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1666464484
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_605
timestamp 1666464484
transform 1 0 69104 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_669
timestamp 1666464484
transform 1 0 76272 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_673
timestamp 1666464484
transform 1 0 76720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_676
timestamp 1666464484
transform 1 0 77056 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_684
timestamp 1666464484
transform 1 0 77952 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_2
timestamp 1666464484
transform 1 0 1568 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_17
timestamp 1666464484
transform 1 0 3248 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_21
timestamp 1666464484
transform 1 0 3696 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_53
timestamp 1666464484
transform 1 0 7280 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_69
timestamp 1666464484
transform 1 0 9072 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1666464484
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1666464484
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1666464484
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_144
timestamp 1666464484
transform 1 0 17472 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_148
timestamp 1666464484
transform 1 0 17920 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_151
timestamp 1666464484
transform 1 0 18256 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_159
timestamp 1666464484
transform 1 0 19152 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_165
timestamp 1666464484
transform 1 0 19824 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_169
timestamp 1666464484
transform 1 0 20272 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_171
timestamp 1666464484
transform 1 0 20496 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_178
timestamp 1666464484
transform 1 0 21280 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_182
timestamp 1666464484
transform 1 0 21728 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_198
timestamp 1666464484
transform 1 0 23520 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_206
timestamp 1666464484
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_210
timestamp 1666464484
transform 1 0 24864 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1666464484
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1666464484
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1666464484
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1666464484
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1666464484
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1666464484
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1666464484
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1666464484
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1666464484
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1666464484
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_428
timestamp 1666464484
transform 1 0 49280 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_460
timestamp 1666464484
transform 1 0 52864 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_468
timestamp 1666464484
transform 1 0 53760 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_472
timestamp 1666464484
transform 1 0 54208 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_474
timestamp 1666464484
transform 1 0 54432 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_477
timestamp 1666464484
transform 1 0 54768 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_481
timestamp 1666464484
transform 1 0 55216 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1666464484
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1666464484
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1666464484
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_563
timestamp 1666464484
transform 1 0 64400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1666464484
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1666464484
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1666464484
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1666464484
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_641
timestamp 1666464484
transform 1 0 73136 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_649
timestamp 1666464484
transform 1 0 74032 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_655
timestamp 1666464484
transform 1 0 74704 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_671
timestamp 1666464484
transform 1 0 76496 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_687
timestamp 1666464484
transform 1 0 78288 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_2
timestamp 1666464484
transform 1 0 1568 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_17
timestamp 1666464484
transform 1 0 3248 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_21
timestamp 1666464484
transform 1 0 3696 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_29
timestamp 1666464484
transform 1 0 4592 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_33
timestamp 1666464484
transform 1 0 5040 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1666464484
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1666464484
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1666464484
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_108
timestamp 1666464484
transform 1 0 13440 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_140
timestamp 1666464484
transform 1 0 17024 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_148
timestamp 1666464484
transform 1 0 17920 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_151
timestamp 1666464484
transform 1 0 18256 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_159
timestamp 1666464484
transform 1 0 19152 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_167
timestamp 1666464484
transform 1 0 20048 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_175
timestamp 1666464484
transform 1 0 20944 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_179
timestamp 1666464484
transform 1 0 21392 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_186
timestamp 1666464484
transform 1 0 22176 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_218
timestamp 1666464484
transform 1 0 25760 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_234
timestamp 1666464484
transform 1 0 27552 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_242
timestamp 1666464484
transform 1 0 28448 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_246
timestamp 1666464484
transform 1 0 28896 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1666464484
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1666464484
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1666464484
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1666464484
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1666464484
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1666464484
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1666464484
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1666464484
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1666464484
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1666464484
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_527
timestamp 1666464484
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1666464484
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1666464484
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_598
timestamp 1666464484
transform 1 0 68320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1666464484
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_605
timestamp 1666464484
transform 1 0 69104 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_669
timestamp 1666464484
transform 1 0 76272 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_673
timestamp 1666464484
transform 1 0 76720 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_676
timestamp 1666464484
transform 1 0 77056 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_684
timestamp 1666464484
transform 1 0 77952 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_2
timestamp 1666464484
transform 1 0 1568 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_17
timestamp 1666464484
transform 1 0 3248 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_21
timestamp 1666464484
transform 1 0 3696 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_53
timestamp 1666464484
transform 1 0 7280 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_69
timestamp 1666464484
transform 1 0 9072 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1666464484
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1666464484
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1666464484
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_144
timestamp 1666464484
transform 1 0 17472 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_160
timestamp 1666464484
transform 1 0 19264 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_163
timestamp 1666464484
transform 1 0 19600 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_171
timestamp 1666464484
transform 1 0 20496 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_179
timestamp 1666464484
transform 1 0 21392 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_183
timestamp 1666464484
transform 1 0 21840 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_185
timestamp 1666464484
transform 1 0 22064 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_188
timestamp 1666464484
transform 1 0 22400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_194
timestamp 1666464484
transform 1 0 23072 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_210
timestamp 1666464484
transform 1 0 24864 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1666464484
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1666464484
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1666464484
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1666464484
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1666464484
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1666464484
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1666464484
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1666464484
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1666464484
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1666464484
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1666464484
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1666464484
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1666464484
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1666464484
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_563
timestamp 1666464484
transform 1 0 64400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1666464484
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1666464484
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_634
timestamp 1666464484
transform 1 0 72352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1666464484
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_641
timestamp 1666464484
transform 1 0 73136 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_649
timestamp 1666464484
transform 1 0 74032 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_655
timestamp 1666464484
transform 1 0 74704 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_671
timestamp 1666464484
transform 1 0 76496 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_687
timestamp 1666464484
transform 1 0 78288 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_2
timestamp 1666464484
transform 1 0 1568 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_17
timestamp 1666464484
transform 1 0 3248 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_21
timestamp 1666464484
transform 1 0 3696 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_25
timestamp 1666464484
transform 1 0 4144 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_33
timestamp 1666464484
transform 1 0 5040 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1666464484
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1666464484
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1666464484
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_108
timestamp 1666464484
transform 1 0 13440 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_140
timestamp 1666464484
transform 1 0 17024 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_156
timestamp 1666464484
transform 1 0 18816 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_164
timestamp 1666464484
transform 1 0 19712 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_168
timestamp 1666464484
transform 1 0 20160 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_170
timestamp 1666464484
transform 1 0 20384 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_173
timestamp 1666464484
transform 1 0 20720 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_179
timestamp 1666464484
transform 1 0 21392 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_186
timestamp 1666464484
transform 1 0 22176 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_190
timestamp 1666464484
transform 1 0 22624 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_200
timestamp 1666464484
transform 1 0 23744 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_232
timestamp 1666464484
transform 1 0 27328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1666464484
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1666464484
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1666464484
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1666464484
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1666464484
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1666464484
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1666464484
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1666464484
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1666464484
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1666464484
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_527
timestamp 1666464484
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1666464484
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1666464484
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_598
timestamp 1666464484
transform 1 0 68320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1666464484
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_605
timestamp 1666464484
transform 1 0 69104 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_637
timestamp 1666464484
transform 1 0 72688 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_653
timestamp 1666464484
transform 1 0 74480 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_657
timestamp 1666464484
transform 1 0 74928 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_673
timestamp 1666464484
transform 1 0 76720 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_676
timestamp 1666464484
transform 1 0 77056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_679
timestamp 1666464484
transform 1 0 77392 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_687
timestamp 1666464484
transform 1 0 78288 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1666464484
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_17
timestamp 1666464484
transform 1 0 3248 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_33
timestamp 1666464484
transform 1 0 5040 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_37
timestamp 1666464484
transform 1 0 5488 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_69
timestamp 1666464484
transform 1 0 9072 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1666464484
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1666464484
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1666464484
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_144
timestamp 1666464484
transform 1 0 17472 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_176
timestamp 1666464484
transform 1 0 21056 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_186
timestamp 1666464484
transform 1 0 22176 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_192
timestamp 1666464484
transform 1 0 22848 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_196
timestamp 1666464484
transform 1 0 23296 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_204
timestamp 1666464484
transform 1 0 24192 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1666464484
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1666464484
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1666464484
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1666464484
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1666464484
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1666464484
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1666464484
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1666464484
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1666464484
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1666464484
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1666464484
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1666464484
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1666464484
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1666464484
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_563
timestamp 1666464484
transform 1 0 64400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1666464484
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1666464484
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_634
timestamp 1666464484
transform 1 0 72352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1666464484
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_641
timestamp 1666464484
transform 1 0 73136 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_649
timestamp 1666464484
transform 1 0 74032 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_655
timestamp 1666464484
transform 1 0 74704 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_671
timestamp 1666464484
transform 1 0 76496 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_687
timestamp 1666464484
transform 1 0 78288 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1666464484
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_17
timestamp 1666464484
transform 1 0 3248 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_21
timestamp 1666464484
transform 1 0 3696 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_29
timestamp 1666464484
transform 1 0 4592 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_33
timestamp 1666464484
transform 1 0 5040 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1666464484
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1666464484
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1666464484
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1666464484
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1666464484
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1666464484
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_179
timestamp 1666464484
transform 1 0 21392 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_182
timestamp 1666464484
transform 1 0 21728 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_190
timestamp 1666464484
transform 1 0 22624 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_198
timestamp 1666464484
transform 1 0 23520 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_230
timestamp 1666464484
transform 1 0 27104 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_246
timestamp 1666464484
transform 1 0 28896 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1666464484
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1666464484
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1666464484
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1666464484
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1666464484
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1666464484
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1666464484
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1666464484
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1666464484
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1666464484
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_527
timestamp 1666464484
transform 1 0 60368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1666464484
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1666464484
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_598
timestamp 1666464484
transform 1 0 68320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1666464484
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_605
timestamp 1666464484
transform 1 0 69104 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_669
timestamp 1666464484
transform 1 0 76272 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1666464484
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_676
timestamp 1666464484
transform 1 0 77056 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_684
timestamp 1666464484
transform 1 0 77952 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_2
timestamp 1666464484
transform 1 0 1568 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_17
timestamp 1666464484
transform 1 0 3248 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_21
timestamp 1666464484
transform 1 0 3696 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_53
timestamp 1666464484
transform 1 0 7280 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_69
timestamp 1666464484
transform 1 0 9072 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1666464484
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1666464484
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1666464484
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_144
timestamp 1666464484
transform 1 0 17472 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_176
timestamp 1666464484
transform 1 0 21056 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_184
timestamp 1666464484
transform 1 0 21952 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_186
timestamp 1666464484
transform 1 0 22176 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_193
timestamp 1666464484
transform 1 0 22960 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_203
timestamp 1666464484
transform 1 0 24080 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_207
timestamp 1666464484
transform 1 0 24528 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_211
timestamp 1666464484
transform 1 0 24976 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_215
timestamp 1666464484
transform 1 0 25424 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_218
timestamp 1666464484
transform 1 0 25760 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_222
timestamp 1666464484
transform 1 0 26208 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_254
timestamp 1666464484
transform 1 0 29792 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_270
timestamp 1666464484
transform 1 0 31584 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_278
timestamp 1666464484
transform 1 0 32480 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_282
timestamp 1666464484
transform 1 0 32928 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1666464484
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1666464484
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1666464484
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1666464484
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1666464484
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1666464484
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1666464484
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1666464484
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1666464484
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1666464484
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_563
timestamp 1666464484
transform 1 0 64400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1666464484
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1666464484
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1666464484
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1666464484
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_641
timestamp 1666464484
transform 1 0 73136 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_649
timestamp 1666464484
transform 1 0 74032 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_655
timestamp 1666464484
transform 1 0 74704 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_671
timestamp 1666464484
transform 1 0 76496 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_687
timestamp 1666464484
transform 1 0 78288 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_2
timestamp 1666464484
transform 1 0 1568 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_17
timestamp 1666464484
transform 1 0 3248 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_21
timestamp 1666464484
transform 1 0 3696 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_29
timestamp 1666464484
transform 1 0 4592 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_33
timestamp 1666464484
transform 1 0 5040 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1666464484
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1666464484
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1666464484
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1666464484
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1666464484
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1666464484
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_179
timestamp 1666464484
transform 1 0 21392 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_187
timestamp 1666464484
transform 1 0 22288 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_191
timestamp 1666464484
transform 1 0 22736 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_195
timestamp 1666464484
transform 1 0 23184 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_197
timestamp 1666464484
transform 1 0 23408 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_204
timestamp 1666464484
transform 1 0 24192 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_210
timestamp 1666464484
transform 1 0 24864 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_220
timestamp 1666464484
transform 1 0 25984 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_228
timestamp 1666464484
transform 1 0 26880 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_244
timestamp 1666464484
transform 1 0 28672 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1666464484
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1666464484
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1666464484
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1666464484
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1666464484
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1666464484
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1666464484
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1666464484
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1666464484
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1666464484
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_527
timestamp 1666464484
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1666464484
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1666464484
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_598
timestamp 1666464484
transform 1 0 68320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1666464484
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605
timestamp 1666464484
transform 1 0 69104 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_669
timestamp 1666464484
transform 1 0 76272 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1666464484
transform 1 0 76720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_676
timestamp 1666464484
transform 1 0 77056 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_684
timestamp 1666464484
transform 1 0 77952 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_2
timestamp 1666464484
transform 1 0 1568 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_17
timestamp 1666464484
transform 1 0 3248 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_21
timestamp 1666464484
transform 1 0 3696 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_53
timestamp 1666464484
transform 1 0 7280 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_69
timestamp 1666464484
transform 1 0 9072 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1666464484
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1666464484
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1666464484
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_144
timestamp 1666464484
transform 1 0 17472 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_176
timestamp 1666464484
transform 1 0 21056 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_192
timestamp 1666464484
transform 1 0 22848 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_200
timestamp 1666464484
transform 1 0 23744 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_208
timestamp 1666464484
transform 1 0 24640 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1666464484
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_215
timestamp 1666464484
transform 1 0 25424 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_223
timestamp 1666464484
transform 1 0 26320 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_227
timestamp 1666464484
transform 1 0 26768 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_231
timestamp 1666464484
transform 1 0 27216 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_263
timestamp 1666464484
transform 1 0 30800 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1666464484
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1666464484
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1666464484
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1666464484
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1666464484
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1666464484
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1666464484
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1666464484
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1666464484
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1666464484
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1666464484
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1666464484
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_563
timestamp 1666464484
transform 1 0 64400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1666464484
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1666464484
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1666464484
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1666464484
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_641
timestamp 1666464484
transform 1 0 73136 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_649
timestamp 1666464484
transform 1 0 74032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_655
timestamp 1666464484
transform 1 0 74704 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_671
timestamp 1666464484
transform 1 0 76496 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_687
timestamp 1666464484
transform 1 0 78288 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_2
timestamp 1666464484
transform 1 0 1568 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_17
timestamp 1666464484
transform 1 0 3248 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_21
timestamp 1666464484
transform 1 0 3696 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_25
timestamp 1666464484
transform 1 0 4144 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_33
timestamp 1666464484
transform 1 0 5040 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1666464484
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1666464484
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1666464484
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1666464484
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1666464484
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1666464484
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_179
timestamp 1666464484
transform 1 0 21392 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_195
timestamp 1666464484
transform 1 0 23184 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_203
timestamp 1666464484
transform 1 0 24080 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_210
timestamp 1666464484
transform 1 0 24864 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_218
timestamp 1666464484
transform 1 0 25760 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_228
timestamp 1666464484
transform 1 0 26880 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_232
timestamp 1666464484
transform 1 0 27328 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_236
timestamp 1666464484
transform 1 0 27776 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_244
timestamp 1666464484
transform 1 0 28672 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1666464484
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1666464484
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1666464484
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1666464484
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1666464484
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1666464484
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1666464484
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1666464484
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1666464484
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1666464484
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_527
timestamp 1666464484
transform 1 0 60368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1666464484
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1666464484
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1666464484
transform 1 0 68320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1666464484
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_605
timestamp 1666464484
transform 1 0 69104 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_637
timestamp 1666464484
transform 1 0 72688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_653
timestamp 1666464484
transform 1 0 74480 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_657
timestamp 1666464484
transform 1 0 74928 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1666464484
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_676
timestamp 1666464484
transform 1 0 77056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_679
timestamp 1666464484
transform 1 0 77392 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_687
timestamp 1666464484
transform 1 0 78288 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_2
timestamp 1666464484
transform 1 0 1568 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_17
timestamp 1666464484
transform 1 0 3248 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_33
timestamp 1666464484
transform 1 0 5040 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_37
timestamp 1666464484
transform 1 0 5488 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_69
timestamp 1666464484
transform 1 0 9072 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1666464484
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1666464484
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1666464484
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1666464484
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1666464484
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1666464484
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_215
timestamp 1666464484
transform 1 0 25424 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_219
timestamp 1666464484
transform 1 0 25872 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_227
timestamp 1666464484
transform 1 0 26768 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_237
timestamp 1666464484
transform 1 0 27888 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_269
timestamp 1666464484
transform 1 0 31472 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_277
timestamp 1666464484
transform 1 0 32368 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_281
timestamp 1666464484
transform 1 0 32816 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1666464484
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1666464484
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1666464484
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1666464484
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1666464484
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1666464484
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1666464484
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1666464484
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1666464484
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1666464484
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1666464484
transform 1 0 57232 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_563
timestamp 1666464484
transform 1 0 64400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1666464484
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1666464484
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1666464484
transform 1 0 72352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1666464484
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_641
timestamp 1666464484
transform 1 0 73136 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_649
timestamp 1666464484
transform 1 0 74032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_655
timestamp 1666464484
transform 1 0 74704 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_671
timestamp 1666464484
transform 1 0 76496 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_687
timestamp 1666464484
transform 1 0 78288 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_2
timestamp 1666464484
transform 1 0 1568 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_17
timestamp 1666464484
transform 1 0 3248 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_21
timestamp 1666464484
transform 1 0 3696 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_29
timestamp 1666464484
transform 1 0 4592 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_33
timestamp 1666464484
transform 1 0 5040 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1666464484
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1666464484
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1666464484
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1666464484
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1666464484
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1666464484
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_179
timestamp 1666464484
transform 1 0 21392 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_211
timestamp 1666464484
transform 1 0 24976 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_219
timestamp 1666464484
transform 1 0 25872 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_225
timestamp 1666464484
transform 1 0 26544 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_233
timestamp 1666464484
transform 1 0 27440 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_243
timestamp 1666464484
transform 1 0 28560 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1666464484
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1666464484
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1666464484
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1666464484
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1666464484
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1666464484
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1666464484
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1666464484
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1666464484
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1666464484
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1666464484
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1666464484
transform 1 0 60368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1666464484
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1666464484
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1666464484
transform 1 0 68320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1666464484
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1666464484
transform 1 0 69104 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_669
timestamp 1666464484
transform 1 0 76272 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1666464484
transform 1 0 76720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_676
timestamp 1666464484
transform 1 0 77056 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_684
timestamp 1666464484
transform 1 0 77952 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_2
timestamp 1666464484
transform 1 0 1568 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_17
timestamp 1666464484
transform 1 0 3248 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_21
timestamp 1666464484
transform 1 0 3696 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_53
timestamp 1666464484
transform 1 0 7280 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_69
timestamp 1666464484
transform 1 0 9072 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1666464484
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1666464484
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1666464484
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1666464484
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1666464484
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1666464484
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_215
timestamp 1666464484
transform 1 0 25424 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_223
timestamp 1666464484
transform 1 0 26320 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_227
timestamp 1666464484
transform 1 0 26768 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_231
timestamp 1666464484
transform 1 0 27216 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_239
timestamp 1666464484
transform 1 0 28112 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_241
timestamp 1666464484
transform 1 0 28336 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_248
timestamp 1666464484
transform 1 0 29120 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_252
timestamp 1666464484
transform 1 0 29568 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_256
timestamp 1666464484
transform 1 0 30016 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_272
timestamp 1666464484
transform 1 0 31808 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_280
timestamp 1666464484
transform 1 0 32704 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1666464484
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1666464484
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1666464484
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1666464484
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1666464484
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1666464484
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1666464484
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1666464484
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1666464484
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1666464484
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1666464484
transform 1 0 64400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1666464484
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1666464484
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1666464484
transform 1 0 72352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1666464484
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_641
timestamp 1666464484
transform 1 0 73136 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_649
timestamp 1666464484
transform 1 0 74032 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_655
timestamp 1666464484
transform 1 0 74704 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_671
timestamp 1666464484
transform 1 0 76496 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_687
timestamp 1666464484
transform 1 0 78288 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_2
timestamp 1666464484
transform 1 0 1568 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_17
timestamp 1666464484
transform 1 0 3248 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_21
timestamp 1666464484
transform 1 0 3696 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_29
timestamp 1666464484
transform 1 0 4592 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_33
timestamp 1666464484
transform 1 0 5040 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1666464484
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1666464484
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1666464484
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1666464484
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1666464484
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1666464484
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_179
timestamp 1666464484
transform 1 0 21392 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_211
timestamp 1666464484
transform 1 0 24976 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_227
timestamp 1666464484
transform 1 0 26768 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_237
timestamp 1666464484
transform 1 0 27888 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_245
timestamp 1666464484
transform 1 0 28784 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1666464484
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_250
timestamp 1666464484
transform 1 0 29344 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_257
timestamp 1666464484
transform 1 0 30128 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_261
timestamp 1666464484
transform 1 0 30576 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_265
timestamp 1666464484
transform 1 0 31024 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_297
timestamp 1666464484
transform 1 0 34608 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_313
timestamp 1666464484
transform 1 0 36400 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_317
timestamp 1666464484
transform 1 0 36848 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1666464484
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1666464484
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1666464484
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1666464484
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1666464484
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1666464484
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1666464484
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1666464484
transform 1 0 60368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1666464484
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1666464484
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1666464484
transform 1 0 68320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1666464484
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1666464484
transform 1 0 69104 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_669
timestamp 1666464484
transform 1 0 76272 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1666464484
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_676
timestamp 1666464484
transform 1 0 77056 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_684
timestamp 1666464484
transform 1 0 77952 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_2
timestamp 1666464484
transform 1 0 1568 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_17
timestamp 1666464484
transform 1 0 3248 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_21
timestamp 1666464484
transform 1 0 3696 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_53
timestamp 1666464484
transform 1 0 7280 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_69
timestamp 1666464484
transform 1 0 9072 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1666464484
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1666464484
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1666464484
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1666464484
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1666464484
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1666464484
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_215
timestamp 1666464484
transform 1 0 25424 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_231
timestamp 1666464484
transform 1 0 27216 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_241
timestamp 1666464484
transform 1 0 28336 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_249
timestamp 1666464484
transform 1 0 29232 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_257
timestamp 1666464484
transform 1 0 30128 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_265
timestamp 1666464484
transform 1 0 31024 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_269
timestamp 1666464484
transform 1 0 31472 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_277
timestamp 1666464484
transform 1 0 32368 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_281
timestamp 1666464484
transform 1 0 32816 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1666464484
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1666464484
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1666464484
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1666464484
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1666464484
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1666464484
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1666464484
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1666464484
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1666464484
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1666464484
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1666464484
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1666464484
transform 1 0 64400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1666464484
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1666464484
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1666464484
transform 1 0 72352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1666464484
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_641
timestamp 1666464484
transform 1 0 73136 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_649
timestamp 1666464484
transform 1 0 74032 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_655
timestamp 1666464484
transform 1 0 74704 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_671
timestamp 1666464484
transform 1 0 76496 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_687
timestamp 1666464484
transform 1 0 78288 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_2
timestamp 1666464484
transform 1 0 1568 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_17
timestamp 1666464484
transform 1 0 3248 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_21
timestamp 1666464484
transform 1 0 3696 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_25
timestamp 1666464484
transform 1 0 4144 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_33
timestamp 1666464484
transform 1 0 5040 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1666464484
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1666464484
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1666464484
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1666464484
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1666464484
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1666464484
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1666464484
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1666464484
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1666464484
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_250
timestamp 1666464484
transform 1 0 29344 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_256
timestamp 1666464484
transform 1 0 30016 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_264
timestamp 1666464484
transform 1 0 30912 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_272
timestamp 1666464484
transform 1 0 31808 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_276
timestamp 1666464484
transform 1 0 32256 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_308
timestamp 1666464484
transform 1 0 35840 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_316
timestamp 1666464484
transform 1 0 36736 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1666464484
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1666464484
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1666464484
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1666464484
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1666464484
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1666464484
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1666464484
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1666464484
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1666464484
transform 1 0 60368 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1666464484
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1666464484
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1666464484
transform 1 0 68320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1666464484
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_605
timestamp 1666464484
transform 1 0 69104 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_637
timestamp 1666464484
transform 1 0 72688 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_653
timestamp 1666464484
transform 1 0 74480 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_657
timestamp 1666464484
transform 1 0 74928 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1666464484
transform 1 0 76720 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_676
timestamp 1666464484
transform 1 0 77056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_679
timestamp 1666464484
transform 1 0 77392 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_687
timestamp 1666464484
transform 1 0 78288 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_2
timestamp 1666464484
transform 1 0 1568 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_17
timestamp 1666464484
transform 1 0 3248 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_33
timestamp 1666464484
transform 1 0 5040 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_37
timestamp 1666464484
transform 1 0 5488 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_69
timestamp 1666464484
transform 1 0 9072 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1666464484
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1666464484
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1666464484
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1666464484
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1666464484
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1666464484
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_215
timestamp 1666464484
transform 1 0 25424 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_247
timestamp 1666464484
transform 1 0 29008 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_261
timestamp 1666464484
transform 1 0 30576 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_269
timestamp 1666464484
transform 1 0 31472 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_271
timestamp 1666464484
transform 1 0 31696 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_278
timestamp 1666464484
transform 1 0 32480 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_282
timestamp 1666464484
transform 1 0 32928 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1666464484
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1666464484
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1666464484
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1666464484
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1666464484
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1666464484
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1666464484
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1666464484
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1666464484
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1666464484
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1666464484
transform 1 0 64400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1666464484
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1666464484
transform 1 0 65184 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1666464484
transform 1 0 72352 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1666464484
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_641
timestamp 1666464484
transform 1 0 73136 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_649
timestamp 1666464484
transform 1 0 74032 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_655
timestamp 1666464484
transform 1 0 74704 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_671
timestamp 1666464484
transform 1 0 76496 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_687
timestamp 1666464484
transform 1 0 78288 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_2
timestamp 1666464484
transform 1 0 1568 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_17
timestamp 1666464484
transform 1 0 3248 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_21
timestamp 1666464484
transform 1 0 3696 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_29
timestamp 1666464484
transform 1 0 4592 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_33
timestamp 1666464484
transform 1 0 5040 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1666464484
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1666464484
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1666464484
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1666464484
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1666464484
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1666464484
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1666464484
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1666464484
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1666464484
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_250
timestamp 1666464484
transform 1 0 29344 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_258
timestamp 1666464484
transform 1 0 30240 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_260
timestamp 1666464484
transform 1 0 30464 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_263
timestamp 1666464484
transform 1 0 30800 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_267
timestamp 1666464484
transform 1 0 31248 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_275
timestamp 1666464484
transform 1 0 32144 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_277
timestamp 1666464484
transform 1 0 32368 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_284
timestamp 1666464484
transform 1 0 33152 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_288
timestamp 1666464484
transform 1 0 33600 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_292
timestamp 1666464484
transform 1 0 34048 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_308
timestamp 1666464484
transform 1 0 35840 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_316
timestamp 1666464484
transform 1 0 36736 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1666464484
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1666464484
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1666464484
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1666464484
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1666464484
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1666464484
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1666464484
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1666464484
transform 1 0 53200 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1666464484
transform 1 0 60368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1666464484
transform 1 0 60816 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1666464484
transform 1 0 61152 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_598
timestamp 1666464484
transform 1 0 68320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1666464484
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1666464484
transform 1 0 69104 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_669
timestamp 1666464484
transform 1 0 76272 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1666464484
transform 1 0 76720 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_676
timestamp 1666464484
transform 1 0 77056 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_684
timestamp 1666464484
transform 1 0 77952 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_2
timestamp 1666464484
transform 1 0 1568 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_17
timestamp 1666464484
transform 1 0 3248 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_21
timestamp 1666464484
transform 1 0 3696 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_53
timestamp 1666464484
transform 1 0 7280 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_69
timestamp 1666464484
transform 1 0 9072 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1666464484
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1666464484
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1666464484
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1666464484
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1666464484
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1666464484
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_215
timestamp 1666464484
transform 1 0 25424 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_247
timestamp 1666464484
transform 1 0 29008 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_263
timestamp 1666464484
transform 1 0 30800 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_267
timestamp 1666464484
transform 1 0 31248 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_269
timestamp 1666464484
transform 1 0 31472 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_272
timestamp 1666464484
transform 1 0 31808 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_280
timestamp 1666464484
transform 1 0 32704 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_286
timestamp 1666464484
transform 1 0 33376 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_293
timestamp 1666464484
transform 1 0 34160 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_297
timestamp 1666464484
transform 1 0 34608 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_329
timestamp 1666464484
transform 1 0 38192 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_345
timestamp 1666464484
transform 1 0 39984 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_353
timestamp 1666464484
transform 1 0 40880 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1666464484
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1666464484
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1666464484
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1666464484
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1666464484
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1666464484
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_499
timestamp 1666464484
transform 1 0 57232 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_563
timestamp 1666464484
transform 1 0 64400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1666464484
transform 1 0 64848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1666464484
transform 1 0 65184 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_634
timestamp 1666464484
transform 1 0 72352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1666464484
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_641
timestamp 1666464484
transform 1 0 73136 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_649
timestamp 1666464484
transform 1 0 74032 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_655
timestamp 1666464484
transform 1 0 74704 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_671
timestamp 1666464484
transform 1 0 76496 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_687
timestamp 1666464484
transform 1 0 78288 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_2
timestamp 1666464484
transform 1 0 1568 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_17
timestamp 1666464484
transform 1 0 3248 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_21
timestamp 1666464484
transform 1 0 3696 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_29
timestamp 1666464484
transform 1 0 4592 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_33
timestamp 1666464484
transform 1 0 5040 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1666464484
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1666464484
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1666464484
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1666464484
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1666464484
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1666464484
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1666464484
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1666464484
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1666464484
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_250
timestamp 1666464484
transform 1 0 29344 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_266
timestamp 1666464484
transform 1 0 31136 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_274
timestamp 1666464484
transform 1 0 32032 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_276
timestamp 1666464484
transform 1 0 32256 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_279
timestamp 1666464484
transform 1 0 32592 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_287
timestamp 1666464484
transform 1 0 33488 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_297
timestamp 1666464484
transform 1 0 34608 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_301
timestamp 1666464484
transform 1 0 35056 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_317
timestamp 1666464484
transform 1 0 36848 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1666464484
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1666464484
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1666464484
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1666464484
transform 1 0 45248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1666464484
transform 1 0 52416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1666464484
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_463
timestamp 1666464484
transform 1 0 53200 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_527
timestamp 1666464484
transform 1 0 60368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1666464484
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_534
timestamp 1666464484
transform 1 0 61152 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_598
timestamp 1666464484
transform 1 0 68320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1666464484
transform 1 0 68768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_605
timestamp 1666464484
transform 1 0 69104 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_669
timestamp 1666464484
transform 1 0 76272 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1666464484
transform 1 0 76720 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_676
timestamp 1666464484
transform 1 0 77056 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_684
timestamp 1666464484
transform 1 0 77952 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_2
timestamp 1666464484
transform 1 0 1568 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_17
timestamp 1666464484
transform 1 0 3248 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_21
timestamp 1666464484
transform 1 0 3696 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_53
timestamp 1666464484
transform 1 0 7280 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_69
timestamp 1666464484
transform 1 0 9072 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1666464484
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1666464484
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1666464484
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1666464484
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1666464484
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1666464484
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1666464484
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_279
timestamp 1666464484
transform 1 0 32592 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1666464484
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_286
timestamp 1666464484
transform 1 0 33376 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_293
timestamp 1666464484
transform 1 0 34160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_303
timestamp 1666464484
transform 1 0 35280 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_305
timestamp 1666464484
transform 1 0 35504 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_308
timestamp 1666464484
transform 1 0 35840 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_312
timestamp 1666464484
transform 1 0 36288 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_344
timestamp 1666464484
transform 1 0 39872 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_352
timestamp 1666464484
transform 1 0 40768 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1666464484
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1666464484
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1666464484
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1666464484
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1666464484
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1666464484
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1666464484
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_499
timestamp 1666464484
transform 1 0 57232 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_563
timestamp 1666464484
transform 1 0 64400 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1666464484
transform 1 0 64848 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_570
timestamp 1666464484
transform 1 0 65184 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_634
timestamp 1666464484
transform 1 0 72352 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1666464484
transform 1 0 72800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_641
timestamp 1666464484
transform 1 0 73136 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_649
timestamp 1666464484
transform 1 0 74032 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_655
timestamp 1666464484
transform 1 0 74704 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_671
timestamp 1666464484
transform 1 0 76496 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_687
timestamp 1666464484
transform 1 0 78288 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_2
timestamp 1666464484
transform 1 0 1568 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_17
timestamp 1666464484
transform 1 0 3248 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_21
timestamp 1666464484
transform 1 0 3696 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_25
timestamp 1666464484
transform 1 0 4144 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_33
timestamp 1666464484
transform 1 0 5040 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1666464484
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1666464484
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1666464484
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1666464484
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1666464484
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1666464484
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1666464484
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1666464484
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1666464484
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_250
timestamp 1666464484
transform 1 0 29344 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_282
timestamp 1666464484
transform 1 0 32928 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_286
timestamp 1666464484
transform 1 0 33376 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_290
timestamp 1666464484
transform 1 0 33824 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_298
timestamp 1666464484
transform 1 0 34720 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_306
timestamp 1666464484
transform 1 0 35616 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_314
timestamp 1666464484
transform 1 0 36512 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1666464484
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1666464484
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1666464484
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1666464484
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1666464484
transform 1 0 45248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1666464484
transform 1 0 52416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1666464484
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_463
timestamp 1666464484
transform 1 0 53200 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_527
timestamp 1666464484
transform 1 0 60368 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_534
timestamp 1666464484
transform 1 0 61152 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_598
timestamp 1666464484
transform 1 0 68320 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1666464484
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_605
timestamp 1666464484
transform 1 0 69104 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_637
timestamp 1666464484
transform 1 0 72688 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_653
timestamp 1666464484
transform 1 0 74480 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_657
timestamp 1666464484
transform 1 0 74928 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1666464484
transform 1 0 76720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_676
timestamp 1666464484
transform 1 0 77056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_679
timestamp 1666464484
transform 1 0 77392 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_687
timestamp 1666464484
transform 1 0 78288 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_2
timestamp 1666464484
transform 1 0 1568 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_17
timestamp 1666464484
transform 1 0 3248 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_33
timestamp 1666464484
transform 1 0 5040 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_37
timestamp 1666464484
transform 1 0 5488 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_69
timestamp 1666464484
transform 1 0 9072 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1666464484
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1666464484
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1666464484
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1666464484
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1666464484
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1666464484
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1666464484
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1666464484
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1666464484
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_286
timestamp 1666464484
transform 1 0 33376 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_294
timestamp 1666464484
transform 1 0 34272 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_302
timestamp 1666464484
transform 1 0 35168 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_310
timestamp 1666464484
transform 1 0 36064 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_320
timestamp 1666464484
transform 1 0 37184 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_324
timestamp 1666464484
transform 1 0 37632 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_340
timestamp 1666464484
transform 1 0 39424 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_348
timestamp 1666464484
transform 1 0 40320 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_352
timestamp 1666464484
transform 1 0 40768 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1666464484
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1666464484
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1666464484
transform 1 0 48496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1666464484
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1666464484
transform 1 0 49280 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1666464484
transform 1 0 56448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1666464484
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_499
timestamp 1666464484
transform 1 0 57232 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_563
timestamp 1666464484
transform 1 0 64400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1666464484
transform 1 0 64848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_570
timestamp 1666464484
transform 1 0 65184 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_634
timestamp 1666464484
transform 1 0 72352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1666464484
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_641
timestamp 1666464484
transform 1 0 73136 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_649
timestamp 1666464484
transform 1 0 74032 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_655
timestamp 1666464484
transform 1 0 74704 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_671
timestamp 1666464484
transform 1 0 76496 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_687
timestamp 1666464484
transform 1 0 78288 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_2
timestamp 1666464484
transform 1 0 1568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_17
timestamp 1666464484
transform 1 0 3248 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_21
timestamp 1666464484
transform 1 0 3696 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_29
timestamp 1666464484
transform 1 0 4592 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_33
timestamp 1666464484
transform 1 0 5040 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1666464484
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1666464484
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1666464484
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1666464484
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1666464484
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1666464484
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1666464484
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1666464484
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1666464484
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_250
timestamp 1666464484
transform 1 0 29344 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_282
timestamp 1666464484
transform 1 0 32928 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_298
timestamp 1666464484
transform 1 0 34720 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_304
timestamp 1666464484
transform 1 0 35392 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_306
timestamp 1666464484
transform 1 0 35616 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_309
timestamp 1666464484
transform 1 0 35952 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_317
timestamp 1666464484
transform 1 0 36848 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_321
timestamp 1666464484
transform 1 0 37296 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_328
timestamp 1666464484
transform 1 0 38080 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_332
timestamp 1666464484
transform 1 0 38528 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_336
timestamp 1666464484
transform 1 0 38976 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_368
timestamp 1666464484
transform 1 0 42560 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_384
timestamp 1666464484
transform 1 0 44352 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_388
timestamp 1666464484
transform 1 0 44800 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_392
timestamp 1666464484
transform 1 0 45248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_456
timestamp 1666464484
transform 1 0 52416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1666464484
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_463
timestamp 1666464484
transform 1 0 53200 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_527
timestamp 1666464484
transform 1 0 60368 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_531
timestamp 1666464484
transform 1 0 60816 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_534
timestamp 1666464484
transform 1 0 61152 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_598
timestamp 1666464484
transform 1 0 68320 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_602
timestamp 1666464484
transform 1 0 68768 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_605
timestamp 1666464484
transform 1 0 69104 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_669
timestamp 1666464484
transform 1 0 76272 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_673
timestamp 1666464484
transform 1 0 76720 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_676
timestamp 1666464484
transform 1 0 77056 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_684
timestamp 1666464484
transform 1 0 77952 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_2
timestamp 1666464484
transform 1 0 1568 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_17
timestamp 1666464484
transform 1 0 3248 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_21
timestamp 1666464484
transform 1 0 3696 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_53
timestamp 1666464484
transform 1 0 7280 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_69
timestamp 1666464484
transform 1 0 9072 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1666464484
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1666464484
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1666464484
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1666464484
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1666464484
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1666464484
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1666464484
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1666464484
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1666464484
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_286
timestamp 1666464484
transform 1 0 33376 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_302
timestamp 1666464484
transform 1 0 35168 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_310
timestamp 1666464484
transform 1 0 36064 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_312
timestamp 1666464484
transform 1 0 36288 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_315
timestamp 1666464484
transform 1 0 36624 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_323
timestamp 1666464484
transform 1 0 37520 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_325
timestamp 1666464484
transform 1 0 37744 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_332
timestamp 1666464484
transform 1 0 38528 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_336
timestamp 1666464484
transform 1 0 38976 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_352
timestamp 1666464484
transform 1 0 40768 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1666464484
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_357
timestamp 1666464484
transform 1 0 41328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_421
timestamp 1666464484
transform 1 0 48496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1666464484
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_428
timestamp 1666464484
transform 1 0 49280 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_492
timestamp 1666464484
transform 1 0 56448 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_496
timestamp 1666464484
transform 1 0 56896 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_499
timestamp 1666464484
transform 1 0 57232 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_563
timestamp 1666464484
transform 1 0 64400 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_567
timestamp 1666464484
transform 1 0 64848 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_570
timestamp 1666464484
transform 1 0 65184 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_634
timestamp 1666464484
transform 1 0 72352 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_638
timestamp 1666464484
transform 1 0 72800 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_641
timestamp 1666464484
transform 1 0 73136 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_649
timestamp 1666464484
transform 1 0 74032 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_655
timestamp 1666464484
transform 1 0 74704 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_671
timestamp 1666464484
transform 1 0 76496 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_687
timestamp 1666464484
transform 1 0 78288 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_2
timestamp 1666464484
transform 1 0 1568 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_17
timestamp 1666464484
transform 1 0 3248 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_21
timestamp 1666464484
transform 1 0 3696 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_29
timestamp 1666464484
transform 1 0 4592 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_33
timestamp 1666464484
transform 1 0 5040 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1666464484
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1666464484
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1666464484
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1666464484
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1666464484
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1666464484
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1666464484
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1666464484
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1666464484
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1666464484
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1666464484
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1666464484
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_321
timestamp 1666464484
transform 1 0 37296 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_329
timestamp 1666464484
transform 1 0 38192 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_331
timestamp 1666464484
transform 1 0 38416 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_338
timestamp 1666464484
transform 1 0 39200 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_342
timestamp 1666464484
transform 1 0 39648 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_374
timestamp 1666464484
transform 1 0 43232 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_392
timestamp 1666464484
transform 1 0 45248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_456
timestamp 1666464484
transform 1 0 52416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1666464484
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_463
timestamp 1666464484
transform 1 0 53200 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_527
timestamp 1666464484
transform 1 0 60368 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_531
timestamp 1666464484
transform 1 0 60816 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_534
timestamp 1666464484
transform 1 0 61152 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_598
timestamp 1666464484
transform 1 0 68320 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_602
timestamp 1666464484
transform 1 0 68768 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_605
timestamp 1666464484
transform 1 0 69104 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_669
timestamp 1666464484
transform 1 0 76272 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_673
timestamp 1666464484
transform 1 0 76720 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_676
timestamp 1666464484
transform 1 0 77056 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_684
timestamp 1666464484
transform 1 0 77952 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_2
timestamp 1666464484
transform 1 0 1568 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_17
timestamp 1666464484
transform 1 0 3248 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_21
timestamp 1666464484
transform 1 0 3696 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_53
timestamp 1666464484
transform 1 0 7280 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_69
timestamp 1666464484
transform 1 0 9072 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1666464484
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1666464484
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1666464484
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1666464484
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1666464484
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1666464484
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1666464484
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1666464484
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1666464484
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_286
timestamp 1666464484
transform 1 0 33376 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_318
timestamp 1666464484
transform 1 0 36960 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_322
timestamp 1666464484
transform 1 0 37408 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_324
timestamp 1666464484
transform 1 0 37632 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_327
timestamp 1666464484
transform 1 0 37968 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_335
timestamp 1666464484
transform 1 0 38864 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_345
timestamp 1666464484
transform 1 0 39984 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_349
timestamp 1666464484
transform 1 0 40432 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_353
timestamp 1666464484
transform 1 0 40880 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_357
timestamp 1666464484
transform 1 0 41328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_421
timestamp 1666464484
transform 1 0 48496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1666464484
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_428
timestamp 1666464484
transform 1 0 49280 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_492
timestamp 1666464484
transform 1 0 56448 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1666464484
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_499
timestamp 1666464484
transform 1 0 57232 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_563
timestamp 1666464484
transform 1 0 64400 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_567
timestamp 1666464484
transform 1 0 64848 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_570
timestamp 1666464484
transform 1 0 65184 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_634
timestamp 1666464484
transform 1 0 72352 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_638
timestamp 1666464484
transform 1 0 72800 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_641
timestamp 1666464484
transform 1 0 73136 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_649
timestamp 1666464484
transform 1 0 74032 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_655
timestamp 1666464484
transform 1 0 74704 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_671
timestamp 1666464484
transform 1 0 76496 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_687
timestamp 1666464484
transform 1 0 78288 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_2
timestamp 1666464484
transform 1 0 1568 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_17
timestamp 1666464484
transform 1 0 3248 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_21
timestamp 1666464484
transform 1 0 3696 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_29
timestamp 1666464484
transform 1 0 4592 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_33
timestamp 1666464484
transform 1 0 5040 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1666464484
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1666464484
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1666464484
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1666464484
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1666464484
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1666464484
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1666464484
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1666464484
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1666464484
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1666464484
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1666464484
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1666464484
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_321
timestamp 1666464484
transform 1 0 37296 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_331
timestamp 1666464484
transform 1 0 38416 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_339
timestamp 1666464484
transform 1 0 39312 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_347
timestamp 1666464484
transform 1 0 40208 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_355
timestamp 1666464484
transform 1 0 41104 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_359
timestamp 1666464484
transform 1 0 41552 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_375
timestamp 1666464484
transform 1 0 43344 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_383
timestamp 1666464484
transform 1 0 44240 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_387
timestamp 1666464484
transform 1 0 44688 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1666464484
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_392
timestamp 1666464484
transform 1 0 45248 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_456
timestamp 1666464484
transform 1 0 52416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_460
timestamp 1666464484
transform 1 0 52864 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_463
timestamp 1666464484
transform 1 0 53200 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_527
timestamp 1666464484
transform 1 0 60368 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_531
timestamp 1666464484
transform 1 0 60816 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_534
timestamp 1666464484
transform 1 0 61152 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_598
timestamp 1666464484
transform 1 0 68320 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_602
timestamp 1666464484
transform 1 0 68768 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_605
timestamp 1666464484
transform 1 0 69104 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_637
timestamp 1666464484
transform 1 0 72688 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_653
timestamp 1666464484
transform 1 0 74480 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_657
timestamp 1666464484
transform 1 0 74928 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_673
timestamp 1666464484
transform 1 0 76720 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_676
timestamp 1666464484
transform 1 0 77056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_679
timestamp 1666464484
transform 1 0 77392 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_687
timestamp 1666464484
transform 1 0 78288 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_2
timestamp 1666464484
transform 1 0 1568 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_17
timestamp 1666464484
transform 1 0 3248 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_21
timestamp 1666464484
transform 1 0 3696 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_53
timestamp 1666464484
transform 1 0 7280 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_69
timestamp 1666464484
transform 1 0 9072 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1666464484
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1666464484
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1666464484
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1666464484
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1666464484
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1666464484
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1666464484
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1666464484
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1666464484
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_286
timestamp 1666464484
transform 1 0 33376 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_318
timestamp 1666464484
transform 1 0 36960 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_336
timestamp 1666464484
transform 1 0 38976 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_344
timestamp 1666464484
transform 1 0 39872 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_352
timestamp 1666464484
transform 1 0 40768 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1666464484
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_357
timestamp 1666464484
transform 1 0 41328 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_364
timestamp 1666464484
transform 1 0 42112 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_368
timestamp 1666464484
transform 1 0 42560 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_400
timestamp 1666464484
transform 1 0 46144 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_416
timestamp 1666464484
transform 1 0 47936 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_424
timestamp 1666464484
transform 1 0 48832 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_428
timestamp 1666464484
transform 1 0 49280 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_492
timestamp 1666464484
transform 1 0 56448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1666464484
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_499
timestamp 1666464484
transform 1 0 57232 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_563
timestamp 1666464484
transform 1 0 64400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_567
timestamp 1666464484
transform 1 0 64848 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_570
timestamp 1666464484
transform 1 0 65184 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_634
timestamp 1666464484
transform 1 0 72352 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_638
timestamp 1666464484
transform 1 0 72800 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_641
timestamp 1666464484
transform 1 0 73136 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_649
timestamp 1666464484
transform 1 0 74032 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_655
timestamp 1666464484
transform 1 0 74704 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_671
timestamp 1666464484
transform 1 0 76496 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_687
timestamp 1666464484
transform 1 0 78288 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_2
timestamp 1666464484
transform 1 0 1568 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_17
timestamp 1666464484
transform 1 0 3248 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_21
timestamp 1666464484
transform 1 0 3696 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_29
timestamp 1666464484
transform 1 0 4592 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_33
timestamp 1666464484
transform 1 0 5040 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1666464484
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1666464484
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1666464484
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1666464484
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1666464484
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1666464484
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1666464484
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1666464484
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1666464484
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1666464484
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1666464484
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1666464484
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_321
timestamp 1666464484
transform 1 0 37296 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_337
timestamp 1666464484
transform 1 0 39088 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_341
timestamp 1666464484
transform 1 0 39536 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_343
timestamp 1666464484
transform 1 0 39760 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_346
timestamp 1666464484
transform 1 0 40096 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_348
timestamp 1666464484
transform 1 0 40320 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_351
timestamp 1666464484
transform 1 0 40656 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_359
timestamp 1666464484
transform 1 0 41552 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_361
timestamp 1666464484
transform 1 0 41776 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_368
timestamp 1666464484
transform 1 0 42560 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_372
timestamp 1666464484
transform 1 0 43008 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_388
timestamp 1666464484
transform 1 0 44800 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_392
timestamp 1666464484
transform 1 0 45248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_456
timestamp 1666464484
transform 1 0 52416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1666464484
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_463
timestamp 1666464484
transform 1 0 53200 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_527
timestamp 1666464484
transform 1 0 60368 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_531
timestamp 1666464484
transform 1 0 60816 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_534
timestamp 1666464484
transform 1 0 61152 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_598
timestamp 1666464484
transform 1 0 68320 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_602
timestamp 1666464484
transform 1 0 68768 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_605
timestamp 1666464484
transform 1 0 69104 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_669
timestamp 1666464484
transform 1 0 76272 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_673
timestamp 1666464484
transform 1 0 76720 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_676
timestamp 1666464484
transform 1 0 77056 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_684
timestamp 1666464484
transform 1 0 77952 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_2
timestamp 1666464484
transform 1 0 1568 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_17
timestamp 1666464484
transform 1 0 3248 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_21
timestamp 1666464484
transform 1 0 3696 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_53
timestamp 1666464484
transform 1 0 7280 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_69
timestamp 1666464484
transform 1 0 9072 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1666464484
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1666464484
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1666464484
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1666464484
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1666464484
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1666464484
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1666464484
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1666464484
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1666464484
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1666464484
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1666464484
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1666464484
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_357
timestamp 1666464484
transform 1 0 41328 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_365
timestamp 1666464484
transform 1 0 42224 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_367
timestamp 1666464484
transform 1 0 42448 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_374
timestamp 1666464484
transform 1 0 43232 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_378
timestamp 1666464484
transform 1 0 43680 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_382
timestamp 1666464484
transform 1 0 44128 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_414
timestamp 1666464484
transform 1 0 47712 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_422
timestamp 1666464484
transform 1 0 48608 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_428
timestamp 1666464484
transform 1 0 49280 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_492
timestamp 1666464484
transform 1 0 56448 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1666464484
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_499
timestamp 1666464484
transform 1 0 57232 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_563
timestamp 1666464484
transform 1 0 64400 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_567
timestamp 1666464484
transform 1 0 64848 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_570
timestamp 1666464484
transform 1 0 65184 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_634
timestamp 1666464484
transform 1 0 72352 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_638
timestamp 1666464484
transform 1 0 72800 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_641
timestamp 1666464484
transform 1 0 73136 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_649
timestamp 1666464484
transform 1 0 74032 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_655
timestamp 1666464484
transform 1 0 74704 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_671
timestamp 1666464484
transform 1 0 76496 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_687
timestamp 1666464484
transform 1 0 78288 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_2
timestamp 1666464484
transform 1 0 1568 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_17
timestamp 1666464484
transform 1 0 3248 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_21
timestamp 1666464484
transform 1 0 3696 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_29
timestamp 1666464484
transform 1 0 4592 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_33
timestamp 1666464484
transform 1 0 5040 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1666464484
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1666464484
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1666464484
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1666464484
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1666464484
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1666464484
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1666464484
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1666464484
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1666464484
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1666464484
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1666464484
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1666464484
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_321
timestamp 1666464484
transform 1 0 37296 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_353
timestamp 1666464484
transform 1 0 40880 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_363
timestamp 1666464484
transform 1 0 42000 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_371
timestamp 1666464484
transform 1 0 42896 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_373
timestamp 1666464484
transform 1 0 43120 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_380
timestamp 1666464484
transform 1 0 43904 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_384
timestamp 1666464484
transform 1 0 44352 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_388
timestamp 1666464484
transform 1 0 44800 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_392
timestamp 1666464484
transform 1 0 45248 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_456
timestamp 1666464484
transform 1 0 52416 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_460
timestamp 1666464484
transform 1 0 52864 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_463
timestamp 1666464484
transform 1 0 53200 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_527
timestamp 1666464484
transform 1 0 60368 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_531
timestamp 1666464484
transform 1 0 60816 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_534
timestamp 1666464484
transform 1 0 61152 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_598
timestamp 1666464484
transform 1 0 68320 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_602
timestamp 1666464484
transform 1 0 68768 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_605
timestamp 1666464484
transform 1 0 69104 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_669
timestamp 1666464484
transform 1 0 76272 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_673
timestamp 1666464484
transform 1 0 76720 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_676
timestamp 1666464484
transform 1 0 77056 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_684
timestamp 1666464484
transform 1 0 77952 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_2
timestamp 1666464484
transform 1 0 1568 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_17
timestamp 1666464484
transform 1 0 3248 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_21
timestamp 1666464484
transform 1 0 3696 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_53
timestamp 1666464484
transform 1 0 7280 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_69
timestamp 1666464484
transform 1 0 9072 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1666464484
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1666464484
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1666464484
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1666464484
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1666464484
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1666464484
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1666464484
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1666464484
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1666464484
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1666464484
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1666464484
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1666464484
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_357
timestamp 1666464484
transform 1 0 41328 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_365
timestamp 1666464484
transform 1 0 42224 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_368
timestamp 1666464484
transform 1 0 42560 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_376
timestamp 1666464484
transform 1 0 43456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_386
timestamp 1666464484
transform 1 0 44576 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_390
timestamp 1666464484
transform 1 0 45024 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_394
timestamp 1666464484
transform 1 0 45472 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_398
timestamp 1666464484
transform 1 0 45920 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_401
timestamp 1666464484
transform 1 0 46256 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_417
timestamp 1666464484
transform 1 0 48048 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1666464484
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_428
timestamp 1666464484
transform 1 0 49280 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_492
timestamp 1666464484
transform 1 0 56448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1666464484
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_499
timestamp 1666464484
transform 1 0 57232 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_563
timestamp 1666464484
transform 1 0 64400 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_567
timestamp 1666464484
transform 1 0 64848 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_570
timestamp 1666464484
transform 1 0 65184 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_634
timestamp 1666464484
transform 1 0 72352 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_638
timestamp 1666464484
transform 1 0 72800 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_641
timestamp 1666464484
transform 1 0 73136 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_657
timestamp 1666464484
transform 1 0 74928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_665
timestamp 1666464484
transform 1 0 75824 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_671
timestamp 1666464484
transform 1 0 76496 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_687
timestamp 1666464484
transform 1 0 78288 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_2
timestamp 1666464484
transform 1 0 1568 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_17
timestamp 1666464484
transform 1 0 3248 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_21
timestamp 1666464484
transform 1 0 3696 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_29
timestamp 1666464484
transform 1 0 4592 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_33
timestamp 1666464484
transform 1 0 5040 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1666464484
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1666464484
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1666464484
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1666464484
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1666464484
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1666464484
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1666464484
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1666464484
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1666464484
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1666464484
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1666464484
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1666464484
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_321
timestamp 1666464484
transform 1 0 37296 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_353
timestamp 1666464484
transform 1 0 40880 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_369
timestamp 1666464484
transform 1 0 42672 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_383
timestamp 1666464484
transform 1 0 44240 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_387
timestamp 1666464484
transform 1 0 44688 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1666464484
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_392
timestamp 1666464484
transform 1 0 45248 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_399
timestamp 1666464484
transform 1 0 46032 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_407
timestamp 1666464484
transform 1 0 46928 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_439
timestamp 1666464484
transform 1 0 50512 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_455
timestamp 1666464484
transform 1 0 52304 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_459
timestamp 1666464484
transform 1 0 52752 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_463
timestamp 1666464484
transform 1 0 53200 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_527
timestamp 1666464484
transform 1 0 60368 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_531
timestamp 1666464484
transform 1 0 60816 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_534
timestamp 1666464484
transform 1 0 61152 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_598
timestamp 1666464484
transform 1 0 68320 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_602
timestamp 1666464484
transform 1 0 68768 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_605
timestamp 1666464484
transform 1 0 69104 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_669
timestamp 1666464484
transform 1 0 76272 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_673
timestamp 1666464484
transform 1 0 76720 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_676
timestamp 1666464484
transform 1 0 77056 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_684
timestamp 1666464484
transform 1 0 77952 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_2
timestamp 1666464484
transform 1 0 1568 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_17
timestamp 1666464484
transform 1 0 3248 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_21
timestamp 1666464484
transform 1 0 3696 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_53
timestamp 1666464484
transform 1 0 7280 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_69
timestamp 1666464484
transform 1 0 9072 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1666464484
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1666464484
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1666464484
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1666464484
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1666464484
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1666464484
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1666464484
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1666464484
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1666464484
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1666464484
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1666464484
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1666464484
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_357
timestamp 1666464484
transform 1 0 41328 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_373
timestamp 1666464484
transform 1 0 43120 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_377
timestamp 1666464484
transform 1 0 43568 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_381
timestamp 1666464484
transform 1 0 44016 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_389
timestamp 1666464484
transform 1 0 44912 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_397
timestamp 1666464484
transform 1 0 45808 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_405
timestamp 1666464484
transform 1 0 46704 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_409
timestamp 1666464484
transform 1 0 47152 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_413
timestamp 1666464484
transform 1 0 47600 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_421
timestamp 1666464484
transform 1 0 48496 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1666464484
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_428
timestamp 1666464484
transform 1 0 49280 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_492
timestamp 1666464484
transform 1 0 56448 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_496
timestamp 1666464484
transform 1 0 56896 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_499
timestamp 1666464484
transform 1 0 57232 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_563
timestamp 1666464484
transform 1 0 64400 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_567
timestamp 1666464484
transform 1 0 64848 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_570
timestamp 1666464484
transform 1 0 65184 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_634
timestamp 1666464484
transform 1 0 72352 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_638
timestamp 1666464484
transform 1 0 72800 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_641
timestamp 1666464484
transform 1 0 73136 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_649
timestamp 1666464484
transform 1 0 74032 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_655
timestamp 1666464484
transform 1 0 74704 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_671
timestamp 1666464484
transform 1 0 76496 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_687
timestamp 1666464484
transform 1 0 78288 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_2
timestamp 1666464484
transform 1 0 1568 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_17
timestamp 1666464484
transform 1 0 3248 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_21
timestamp 1666464484
transform 1 0 3696 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_29
timestamp 1666464484
transform 1 0 4592 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_33
timestamp 1666464484
transform 1 0 5040 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1666464484
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1666464484
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1666464484
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_108
timestamp 1666464484
transform 1 0 13440 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_172
timestamp 1666464484
transform 1 0 20608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1666464484
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_179
timestamp 1666464484
transform 1 0 21392 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_243
timestamp 1666464484
transform 1 0 28560 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1666464484
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_250
timestamp 1666464484
transform 1 0 29344 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_314
timestamp 1666464484
transform 1 0 36512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1666464484
transform 1 0 36960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_321
timestamp 1666464484
transform 1 0 37296 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_385
timestamp 1666464484
transform 1 0 44464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_389
timestamp 1666464484
transform 1 0 44912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_392
timestamp 1666464484
transform 1 0 45248 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_402
timestamp 1666464484
transform 1 0 46368 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_404
timestamp 1666464484
transform 1 0 46592 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_411
timestamp 1666464484
transform 1 0 47376 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_415
timestamp 1666464484
transform 1 0 47824 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_419
timestamp 1666464484
transform 1 0 48272 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_451
timestamp 1666464484
transform 1 0 51856 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_459
timestamp 1666464484
transform 1 0 52752 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_463
timestamp 1666464484
transform 1 0 53200 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_527
timestamp 1666464484
transform 1 0 60368 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_531
timestamp 1666464484
transform 1 0 60816 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_534
timestamp 1666464484
transform 1 0 61152 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_598
timestamp 1666464484
transform 1 0 68320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_602
timestamp 1666464484
transform 1 0 68768 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_605
timestamp 1666464484
transform 1 0 69104 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_637
timestamp 1666464484
transform 1 0 72688 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_653
timestamp 1666464484
transform 1 0 74480 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_657
timestamp 1666464484
transform 1 0 74928 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_673
timestamp 1666464484
transform 1 0 76720 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_676
timestamp 1666464484
transform 1 0 77056 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_684
timestamp 1666464484
transform 1 0 77952 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_2
timestamp 1666464484
transform 1 0 1568 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_17
timestamp 1666464484
transform 1 0 3248 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_21
timestamp 1666464484
transform 1 0 3696 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_53
timestamp 1666464484
transform 1 0 7280 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_69
timestamp 1666464484
transform 1 0 9072 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_73
timestamp 1666464484
transform 1 0 9520 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_137
timestamp 1666464484
transform 1 0 16688 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1666464484
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_144
timestamp 1666464484
transform 1 0 17472 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_208
timestamp 1666464484
transform 1 0 24640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1666464484
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_215
timestamp 1666464484
transform 1 0 25424 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_279
timestamp 1666464484
transform 1 0 32592 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1666464484
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_286
timestamp 1666464484
transform 1 0 33376 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_350
timestamp 1666464484
transform 1 0 40544 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1666464484
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_357
timestamp 1666464484
transform 1 0 41328 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_389
timestamp 1666464484
transform 1 0 44912 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_397
timestamp 1666464484
transform 1 0 45808 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_400
timestamp 1666464484
transform 1 0 46144 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_408
timestamp 1666464484
transform 1 0 47040 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_410
timestamp 1666464484
transform 1 0 47264 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_417
timestamp 1666464484
transform 1 0 48048 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_421
timestamp 1666464484
transform 1 0 48496 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1666464484
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_428
timestamp 1666464484
transform 1 0 49280 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_492
timestamp 1666464484
transform 1 0 56448 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1666464484
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_499
timestamp 1666464484
transform 1 0 57232 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_563
timestamp 1666464484
transform 1 0 64400 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_567
timestamp 1666464484
transform 1 0 64848 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_570
timestamp 1666464484
transform 1 0 65184 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_634
timestamp 1666464484
transform 1 0 72352 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_638
timestamp 1666464484
transform 1 0 72800 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_641
timestamp 1666464484
transform 1 0 73136 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_649
timestamp 1666464484
transform 1 0 74032 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_655
timestamp 1666464484
transform 1 0 74704 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_671
timestamp 1666464484
transform 1 0 76496 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_687
timestamp 1666464484
transform 1 0 78288 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_2
timestamp 1666464484
transform 1 0 1568 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_17
timestamp 1666464484
transform 1 0 3248 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_21
timestamp 1666464484
transform 1 0 3696 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_29
timestamp 1666464484
transform 1 0 4592 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_33
timestamp 1666464484
transform 1 0 5040 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1666464484
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1666464484
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1666464484
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_108
timestamp 1666464484
transform 1 0 13440 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_172
timestamp 1666464484
transform 1 0 20608 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1666464484
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_179
timestamp 1666464484
transform 1 0 21392 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_243
timestamp 1666464484
transform 1 0 28560 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1666464484
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_250
timestamp 1666464484
transform 1 0 29344 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_314
timestamp 1666464484
transform 1 0 36512 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1666464484
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_321
timestamp 1666464484
transform 1 0 37296 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_385
timestamp 1666464484
transform 1 0 44464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1666464484
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_392
timestamp 1666464484
transform 1 0 45248 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_414
timestamp 1666464484
transform 1 0 47712 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_416
timestamp 1666464484
transform 1 0 47936 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_423
timestamp 1666464484
transform 1 0 48720 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_427
timestamp 1666464484
transform 1 0 49168 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_459
timestamp 1666464484
transform 1 0 52752 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_463
timestamp 1666464484
transform 1 0 53200 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_527
timestamp 1666464484
transform 1 0 60368 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_531
timestamp 1666464484
transform 1 0 60816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_534
timestamp 1666464484
transform 1 0 61152 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_598
timestamp 1666464484
transform 1 0 68320 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_602
timestamp 1666464484
transform 1 0 68768 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_605
timestamp 1666464484
transform 1 0 69104 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_669
timestamp 1666464484
transform 1 0 76272 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_673
timestamp 1666464484
transform 1 0 76720 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_676
timestamp 1666464484
transform 1 0 77056 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_684
timestamp 1666464484
transform 1 0 77952 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_2
timestamp 1666464484
transform 1 0 1568 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_17
timestamp 1666464484
transform 1 0 3248 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_21
timestamp 1666464484
transform 1 0 3696 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_53
timestamp 1666464484
transform 1 0 7280 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_69
timestamp 1666464484
transform 1 0 9072 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_73
timestamp 1666464484
transform 1 0 9520 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_137
timestamp 1666464484
transform 1 0 16688 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1666464484
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_144
timestamp 1666464484
transform 1 0 17472 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_208
timestamp 1666464484
transform 1 0 24640 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1666464484
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_215
timestamp 1666464484
transform 1 0 25424 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_279
timestamp 1666464484
transform 1 0 32592 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1666464484
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_286
timestamp 1666464484
transform 1 0 33376 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_350
timestamp 1666464484
transform 1 0 40544 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1666464484
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_357
timestamp 1666464484
transform 1 0 41328 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_389
timestamp 1666464484
transform 1 0 44912 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_405
timestamp 1666464484
transform 1 0 46704 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_409
timestamp 1666464484
transform 1 0 47152 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_412
timestamp 1666464484
transform 1 0 47488 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_416
timestamp 1666464484
transform 1 0 47936 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_418
timestamp 1666464484
transform 1 0 48160 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_423
timestamp 1666464484
transform 1 0 48720 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_425
timestamp 1666464484
transform 1 0 48944 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_428
timestamp 1666464484
transform 1 0 49280 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_430
timestamp 1666464484
transform 1 0 49504 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_435
timestamp 1666464484
transform 1 0 50064 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_439
timestamp 1666464484
transform 1 0 50512 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_471
timestamp 1666464484
transform 1 0 54096 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_487
timestamp 1666464484
transform 1 0 55888 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_495
timestamp 1666464484
transform 1 0 56784 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_499
timestamp 1666464484
transform 1 0 57232 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_563
timestamp 1666464484
transform 1 0 64400 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_567
timestamp 1666464484
transform 1 0 64848 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_570
timestamp 1666464484
transform 1 0 65184 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_586
timestamp 1666464484
transform 1 0 66976 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_594
timestamp 1666464484
transform 1 0 67872 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_598
timestamp 1666464484
transform 1 0 68320 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_600
timestamp 1666464484
transform 1 0 68544 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_605
timestamp 1666464484
transform 1 0 69104 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_609
timestamp 1666464484
transform 1 0 69552 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_613
timestamp 1666464484
transform 1 0 70000 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_629
timestamp 1666464484
transform 1 0 71792 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_637
timestamp 1666464484
transform 1 0 72688 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_641
timestamp 1666464484
transform 1 0 73136 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_649
timestamp 1666464484
transform 1 0 74032 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_655
timestamp 1666464484
transform 1 0 74704 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_671
timestamp 1666464484
transform 1 0 76496 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_687
timestamp 1666464484
transform 1 0 78288 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_2
timestamp 1666464484
transform 1 0 1568 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_17
timestamp 1666464484
transform 1 0 3248 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_21
timestamp 1666464484
transform 1 0 3696 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_29
timestamp 1666464484
transform 1 0 4592 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_33
timestamp 1666464484
transform 1 0 5040 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1666464484
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1666464484
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1666464484
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_108
timestamp 1666464484
transform 1 0 13440 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_172
timestamp 1666464484
transform 1 0 20608 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1666464484
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_179
timestamp 1666464484
transform 1 0 21392 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_243
timestamp 1666464484
transform 1 0 28560 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1666464484
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_250
timestamp 1666464484
transform 1 0 29344 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_314
timestamp 1666464484
transform 1 0 36512 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1666464484
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_321
timestamp 1666464484
transform 1 0 37296 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_385
timestamp 1666464484
transform 1 0 44464 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1666464484
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_392
timestamp 1666464484
transform 1 0 45248 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_408
timestamp 1666464484
transform 1 0 47040 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_412
timestamp 1666464484
transform 1 0 47488 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_414
timestamp 1666464484
transform 1 0 47712 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_419
timestamp 1666464484
transform 1 0 48272 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_423
timestamp 1666464484
transform 1 0 48720 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_435
timestamp 1666464484
transform 1 0 50064 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_441
timestamp 1666464484
transform 1 0 50736 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_445
timestamp 1666464484
transform 1 0 51184 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_463
timestamp 1666464484
transform 1 0 53200 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_527
timestamp 1666464484
transform 1 0 60368 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_531
timestamp 1666464484
transform 1 0 60816 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_534
timestamp 1666464484
transform 1 0 61152 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_566
timestamp 1666464484
transform 1 0 64736 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_582
timestamp 1666464484
transform 1 0 66528 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_590
timestamp 1666464484
transform 1 0 67424 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_598
timestamp 1666464484
transform 1 0 68320 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_602
timestamp 1666464484
transform 1 0 68768 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_605
timestamp 1666464484
transform 1 0 69104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_616
timestamp 1666464484
transform 1 0 70336 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_620
timestamp 1666464484
transform 1 0 70784 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_652
timestamp 1666464484
transform 1 0 74368 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_668
timestamp 1666464484
transform 1 0 76160 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_670
timestamp 1666464484
transform 1 0 76384 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_673
timestamp 1666464484
transform 1 0 76720 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_676
timestamp 1666464484
transform 1 0 77056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_679
timestamp 1666464484
transform 1 0 77392 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_687
timestamp 1666464484
transform 1 0 78288 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_2
timestamp 1666464484
transform 1 0 1568 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_9
timestamp 1666464484
transform 1 0 2352 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_17
timestamp 1666464484
transform 1 0 3248 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_21
timestamp 1666464484
transform 1 0 3696 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_53
timestamp 1666464484
transform 1 0 7280 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_69
timestamp 1666464484
transform 1 0 9072 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_73
timestamp 1666464484
transform 1 0 9520 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_137
timestamp 1666464484
transform 1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1666464484
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_144
timestamp 1666464484
transform 1 0 17472 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_208
timestamp 1666464484
transform 1 0 24640 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1666464484
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_215
timestamp 1666464484
transform 1 0 25424 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_279
timestamp 1666464484
transform 1 0 32592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1666464484
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_286
timestamp 1666464484
transform 1 0 33376 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_350
timestamp 1666464484
transform 1 0 40544 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1666464484
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_357
timestamp 1666464484
transform 1 0 41328 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_389
timestamp 1666464484
transform 1 0 44912 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_397
timestamp 1666464484
transform 1 0 45808 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_401
timestamp 1666464484
transform 1 0 46256 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_406
timestamp 1666464484
transform 1 0 46816 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_410
timestamp 1666464484
transform 1 0 47264 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_428
timestamp 1666464484
transform 1 0 49280 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_439
timestamp 1666464484
transform 1 0 50512 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_451
timestamp 1666464484
transform 1 0 51856 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_457
timestamp 1666464484
transform 1 0 52528 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_461
timestamp 1666464484
transform 1 0 52976 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_493
timestamp 1666464484
transform 1 0 56560 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_499
timestamp 1666464484
transform 1 0 57232 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_563
timestamp 1666464484
transform 1 0 64400 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_567
timestamp 1666464484
transform 1 0 64848 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_570
timestamp 1666464484
transform 1 0 65184 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_602
timestamp 1666464484
transform 1 0 68768 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_605
timestamp 1666464484
transform 1 0 69104 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_617
timestamp 1666464484
transform 1 0 70448 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_621
timestamp 1666464484
transform 1 0 70896 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_637
timestamp 1666464484
transform 1 0 72688 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_641
timestamp 1666464484
transform 1 0 73136 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_673
timestamp 1666464484
transform 1 0 76720 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_679
timestamp 1666464484
transform 1 0 77392 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_687
timestamp 1666464484
transform 1 0 78288 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_2
timestamp 1666464484
transform 1 0 1568 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_9
timestamp 1666464484
transform 1 0 2352 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_13
timestamp 1666464484
transform 1 0 2800 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_17
timestamp 1666464484
transform 1 0 3248 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_33
timestamp 1666464484
transform 1 0 5040 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1666464484
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1666464484
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1666464484
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_108
timestamp 1666464484
transform 1 0 13440 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_172
timestamp 1666464484
transform 1 0 20608 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1666464484
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1666464484
transform 1 0 21392 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1666464484
transform 1 0 28560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1666464484
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_250
timestamp 1666464484
transform 1 0 29344 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_314
timestamp 1666464484
transform 1 0 36512 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1666464484
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_321
timestamp 1666464484
transform 1 0 37296 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_385
timestamp 1666464484
transform 1 0 44464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1666464484
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_392
timestamp 1666464484
transform 1 0 45248 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_424
timestamp 1666464484
transform 1 0 48832 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_428
timestamp 1666464484
transform 1 0 49280 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_434
timestamp 1666464484
transform 1 0 49952 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_446
timestamp 1666464484
transform 1 0 51296 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_452
timestamp 1666464484
transform 1 0 51968 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_456
timestamp 1666464484
transform 1 0 52416 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1666464484
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_463
timestamp 1666464484
transform 1 0 53200 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_470
timestamp 1666464484
transform 1 0 53984 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_486
timestamp 1666464484
transform 1 0 55776 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_494
timestamp 1666464484
transform 1 0 56672 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_500
timestamp 1666464484
transform 1 0 57344 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_534
timestamp 1666464484
transform 1 0 61152 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_598
timestamp 1666464484
transform 1 0 68320 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_602
timestamp 1666464484
transform 1 0 68768 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_605
timestamp 1666464484
transform 1 0 69104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_610
timestamp 1666464484
transform 1 0 69664 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_616
timestamp 1666464484
transform 1 0 70336 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_620
timestamp 1666464484
transform 1 0 70784 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_652
timestamp 1666464484
transform 1 0 74368 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_668
timestamp 1666464484
transform 1 0 76160 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_672
timestamp 1666464484
transform 1 0 76608 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_676
timestamp 1666464484
transform 1 0 77056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_679
timestamp 1666464484
transform 1 0 77392 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_687
timestamp 1666464484
transform 1 0 78288 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_2
timestamp 1666464484
transform 1 0 1568 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_9
timestamp 1666464484
transform 1 0 2352 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_13
timestamp 1666464484
transform 1 0 2800 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_45
timestamp 1666464484
transform 1 0 6384 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_61
timestamp 1666464484
transform 1 0 8176 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_69
timestamp 1666464484
transform 1 0 9072 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_73
timestamp 1666464484
transform 1 0 9520 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_137
timestamp 1666464484
transform 1 0 16688 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1666464484
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_144
timestamp 1666464484
transform 1 0 17472 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_208
timestamp 1666464484
transform 1 0 24640 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1666464484
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1666464484
transform 1 0 25424 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1666464484
transform 1 0 32592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1666464484
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_286
timestamp 1666464484
transform 1 0 33376 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_350
timestamp 1666464484
transform 1 0 40544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1666464484
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_357
timestamp 1666464484
transform 1 0 41328 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_421
timestamp 1666464484
transform 1 0 48496 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1666464484
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_428
timestamp 1666464484
transform 1 0 49280 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_444
timestamp 1666464484
transform 1 0 51072 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_448
timestamp 1666464484
transform 1 0 51520 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_459
timestamp 1666464484
transform 1 0 52752 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_469
timestamp 1666464484
transform 1 0 53872 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_477
timestamp 1666464484
transform 1 0 54768 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_481
timestamp 1666464484
transform 1 0 55216 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_483
timestamp 1666464484
transform 1 0 55440 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_486
timestamp 1666464484
transform 1 0 55776 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_494
timestamp 1666464484
transform 1 0 56672 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1666464484
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_499
timestamp 1666464484
transform 1 0 57232 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_506
timestamp 1666464484
transform 1 0 58016 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_538
timestamp 1666464484
transform 1 0 61600 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_554
timestamp 1666464484
transform 1 0 63392 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_562
timestamp 1666464484
transform 1 0 64288 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_566
timestamp 1666464484
transform 1 0 64736 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_570
timestamp 1666464484
transform 1 0 65184 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_634
timestamp 1666464484
transform 1 0 72352 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_638
timestamp 1666464484
transform 1 0 72800 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_641
timestamp 1666464484
transform 1 0 73136 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_673
timestamp 1666464484
transform 1 0 76720 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_679
timestamp 1666464484
transform 1 0 77392 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_687
timestamp 1666464484
transform 1 0 78288 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_2
timestamp 1666464484
transform 1 0 1568 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_9
timestamp 1666464484
transform 1 0 2352 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_13
timestamp 1666464484
transform 1 0 2800 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_29
timestamp 1666464484
transform 1 0 4592 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_33
timestamp 1666464484
transform 1 0 5040 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1666464484
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1666464484
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1666464484
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1666464484
transform 1 0 13440 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_172
timestamp 1666464484
transform 1 0 20608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1666464484
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1666464484
transform 1 0 21392 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_243
timestamp 1666464484
transform 1 0 28560 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1666464484
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1666464484
transform 1 0 29344 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1666464484
transform 1 0 36512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1666464484
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_321
timestamp 1666464484
transform 1 0 37296 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_385
timestamp 1666464484
transform 1 0 44464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1666464484
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_392
timestamp 1666464484
transform 1 0 45248 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_400
timestamp 1666464484
transform 1 0 46144 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_404
timestamp 1666464484
transform 1 0 46592 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_410
timestamp 1666464484
transform 1 0 47264 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_414
timestamp 1666464484
transform 1 0 47712 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_426
timestamp 1666464484
transform 1 0 49056 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_430
timestamp 1666464484
transform 1 0 49504 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_444
timestamp 1666464484
transform 1 0 51072 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_448
timestamp 1666464484
transform 1 0 51520 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_460
timestamp 1666464484
transform 1 0 52864 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_463
timestamp 1666464484
transform 1 0 53200 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_479
timestamp 1666464484
transform 1 0 54992 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_493
timestamp 1666464484
transform 1 0 56560 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_497
timestamp 1666464484
transform 1 0 57008 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_501
timestamp 1666464484
transform 1 0 57456 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_509
timestamp 1666464484
transform 1 0 58352 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_513
timestamp 1666464484
transform 1 0 58800 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_519
timestamp 1666464484
transform 1 0 59472 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_523
timestamp 1666464484
transform 1 0 59920 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_529
timestamp 1666464484
transform 1 0 60592 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_531
timestamp 1666464484
transform 1 0 60816 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_534
timestamp 1666464484
transform 1 0 61152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_537
timestamp 1666464484
transform 1 0 61488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_601
timestamp 1666464484
transform 1 0 68656 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_605
timestamp 1666464484
transform 1 0 69104 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_669
timestamp 1666464484
transform 1 0 76272 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_673
timestamp 1666464484
transform 1 0 76720 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_676
timestamp 1666464484
transform 1 0 77056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_679
timestamp 1666464484
transform 1 0 77392 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_687
timestamp 1666464484
transform 1 0 78288 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_2
timestamp 1666464484
transform 1 0 1568 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_9
timestamp 1666464484
transform 1 0 2352 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_13
timestamp 1666464484
transform 1 0 2800 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_45
timestamp 1666464484
transform 1 0 6384 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_61
timestamp 1666464484
transform 1 0 8176 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_69
timestamp 1666464484
transform 1 0 9072 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1666464484
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_137
timestamp 1666464484
transform 1 0 16688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1666464484
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1666464484
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1666464484
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1666464484
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1666464484
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1666464484
transform 1 0 32592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1666464484
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_286
timestamp 1666464484
transform 1 0 33376 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_350
timestamp 1666464484
transform 1 0 40544 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1666464484
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_357
timestamp 1666464484
transform 1 0 41328 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_389
timestamp 1666464484
transform 1 0 44912 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_405
timestamp 1666464484
transform 1 0 46704 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_413
timestamp 1666464484
transform 1 0 47600 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_416
timestamp 1666464484
transform 1 0 47936 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_422
timestamp 1666464484
transform 1 0 48608 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_428
timestamp 1666464484
transform 1 0 49280 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_432
timestamp 1666464484
transform 1 0 49728 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_434
timestamp 1666464484
transform 1 0 49952 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_439
timestamp 1666464484
transform 1 0 50512 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_443
timestamp 1666464484
transform 1 0 50960 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_453
timestamp 1666464484
transform 1 0 52080 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_455
timestamp 1666464484
transform 1 0 52304 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_466
timestamp 1666464484
transform 1 0 53536 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_478
timestamp 1666464484
transform 1 0 54880 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_486
timestamp 1666464484
transform 1 0 55776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_490
timestamp 1666464484
transform 1 0 56224 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1666464484
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_499
timestamp 1666464484
transform 1 0 57232 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_506
timestamp 1666464484
transform 1 0 58016 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_538
timestamp 1666464484
transform 1 0 61600 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_554
timestamp 1666464484
transform 1 0 63392 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_562
timestamp 1666464484
transform 1 0 64288 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_566
timestamp 1666464484
transform 1 0 64736 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_570
timestamp 1666464484
transform 1 0 65184 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_634
timestamp 1666464484
transform 1 0 72352 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_638
timestamp 1666464484
transform 1 0 72800 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_641
timestamp 1666464484
transform 1 0 73136 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_673
timestamp 1666464484
transform 1 0 76720 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_679
timestamp 1666464484
transform 1 0 77392 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_687
timestamp 1666464484
transform 1 0 78288 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_2
timestamp 1666464484
transform 1 0 1568 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_9
timestamp 1666464484
transform 1 0 2352 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_13
timestamp 1666464484
transform 1 0 2800 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_17
timestamp 1666464484
transform 1 0 3248 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_33
timestamp 1666464484
transform 1 0 5040 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1666464484
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1666464484
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1666464484
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1666464484
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1666464484
transform 1 0 20608 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1666464484
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1666464484
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1666464484
transform 1 0 28560 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1666464484
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1666464484
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1666464484
transform 1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1666464484
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_321
timestamp 1666464484
transform 1 0 37296 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_385
timestamp 1666464484
transform 1 0 44464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1666464484
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_392
timestamp 1666464484
transform 1 0 45248 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_424
timestamp 1666464484
transform 1 0 48832 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_440
timestamp 1666464484
transform 1 0 50624 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_448
timestamp 1666464484
transform 1 0 51520 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_452
timestamp 1666464484
transform 1 0 51968 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_455
timestamp 1666464484
transform 1 0 52304 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_457
timestamp 1666464484
transform 1 0 52528 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_460
timestamp 1666464484
transform 1 0 52864 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_463
timestamp 1666464484
transform 1 0 53200 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_468
timestamp 1666464484
transform 1 0 53760 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_470
timestamp 1666464484
transform 1 0 53984 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_481
timestamp 1666464484
transform 1 0 55216 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_489
timestamp 1666464484
transform 1 0 56112 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_493
timestamp 1666464484
transform 1 0 56560 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_495
timestamp 1666464484
transform 1 0 56784 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_498
timestamp 1666464484
transform 1 0 57120 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_502
timestamp 1666464484
transform 1 0 57568 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_518
timestamp 1666464484
transform 1 0 59360 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_526
timestamp 1666464484
transform 1 0 60256 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_530
timestamp 1666464484
transform 1 0 60704 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_534
timestamp 1666464484
transform 1 0 61152 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_598
timestamp 1666464484
transform 1 0 68320 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_602
timestamp 1666464484
transform 1 0 68768 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_605
timestamp 1666464484
transform 1 0 69104 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_669
timestamp 1666464484
transform 1 0 76272 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_673
timestamp 1666464484
transform 1 0 76720 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_676
timestamp 1666464484
transform 1 0 77056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_679
timestamp 1666464484
transform 1 0 77392 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_687
timestamp 1666464484
transform 1 0 78288 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_2
timestamp 1666464484
transform 1 0 1568 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_9
timestamp 1666464484
transform 1 0 2352 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_17
timestamp 1666464484
transform 1 0 3248 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_21
timestamp 1666464484
transform 1 0 3696 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_53
timestamp 1666464484
transform 1 0 7280 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_69
timestamp 1666464484
transform 1 0 9072 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1666464484
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1666464484
transform 1 0 16688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1666464484
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1666464484
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1666464484
transform 1 0 24640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1666464484
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1666464484
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1666464484
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1666464484
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1666464484
transform 1 0 33376 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_350
timestamp 1666464484
transform 1 0 40544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1666464484
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_357
timestamp 1666464484
transform 1 0 41328 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_421
timestamp 1666464484
transform 1 0 48496 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1666464484
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_428
timestamp 1666464484
transform 1 0 49280 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_444
timestamp 1666464484
transform 1 0 51072 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_450
timestamp 1666464484
transform 1 0 51744 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_456
timestamp 1666464484
transform 1 0 52416 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_462
timestamp 1666464484
transform 1 0 53088 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_466
timestamp 1666464484
transform 1 0 53536 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_471
timestamp 1666464484
transform 1 0 54096 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_483
timestamp 1666464484
transform 1 0 55440 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_489
timestamp 1666464484
transform 1 0 56112 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_495
timestamp 1666464484
transform 1 0 56784 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_499
timestamp 1666464484
transform 1 0 57232 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_506
timestamp 1666464484
transform 1 0 58016 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_538
timestamp 1666464484
transform 1 0 61600 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_554
timestamp 1666464484
transform 1 0 63392 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_562
timestamp 1666464484
transform 1 0 64288 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_566
timestamp 1666464484
transform 1 0 64736 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_570
timestamp 1666464484
transform 1 0 65184 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_634
timestamp 1666464484
transform 1 0 72352 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_638
timestamp 1666464484
transform 1 0 72800 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_641
timestamp 1666464484
transform 1 0 73136 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_657
timestamp 1666464484
transform 1 0 74928 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_665
timestamp 1666464484
transform 1 0 75824 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_671
timestamp 1666464484
transform 1 0 76496 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_679
timestamp 1666464484
transform 1 0 77392 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_687
timestamp 1666464484
transform 1 0 78288 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_2
timestamp 1666464484
transform 1 0 1568 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_9
timestamp 1666464484
transform 1 0 2352 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_13
timestamp 1666464484
transform 1 0 2800 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_29
timestamp 1666464484
transform 1 0 4592 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_33
timestamp 1666464484
transform 1 0 5040 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1666464484
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1666464484
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1666464484
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_108
timestamp 1666464484
transform 1 0 13440 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_172
timestamp 1666464484
transform 1 0 20608 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1666464484
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1666464484
transform 1 0 21392 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_243
timestamp 1666464484
transform 1 0 28560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1666464484
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1666464484
transform 1 0 29344 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1666464484
transform 1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1666464484
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_321
timestamp 1666464484
transform 1 0 37296 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_385
timestamp 1666464484
transform 1 0 44464 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1666464484
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_392
timestamp 1666464484
transform 1 0 45248 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_424
timestamp 1666464484
transform 1 0 48832 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_432
timestamp 1666464484
transform 1 0 49728 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_440
timestamp 1666464484
transform 1 0 50624 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_444
timestamp 1666464484
transform 1 0 51072 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_452
timestamp 1666464484
transform 1 0 51968 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_458
timestamp 1666464484
transform 1 0 52640 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_460
timestamp 1666464484
transform 1 0 52864 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_463
timestamp 1666464484
transform 1 0 53200 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_467
timestamp 1666464484
transform 1 0 53648 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_475
timestamp 1666464484
transform 1 0 54544 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_477
timestamp 1666464484
transform 1 0 54768 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_488
timestamp 1666464484
transform 1 0 56000 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_492
timestamp 1666464484
transform 1 0 56448 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_494
timestamp 1666464484
transform 1 0 56672 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_501
timestamp 1666464484
transform 1 0 57456 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_505
timestamp 1666464484
transform 1 0 57904 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_521
timestamp 1666464484
transform 1 0 59696 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_529
timestamp 1666464484
transform 1 0 60592 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_531
timestamp 1666464484
transform 1 0 60816 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_534
timestamp 1666464484
transform 1 0 61152 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_598
timestamp 1666464484
transform 1 0 68320 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_602
timestamp 1666464484
transform 1 0 68768 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_605
timestamp 1666464484
transform 1 0 69104 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_669
timestamp 1666464484
transform 1 0 76272 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_673
timestamp 1666464484
transform 1 0 76720 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_676
timestamp 1666464484
transform 1 0 77056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_679
timestamp 1666464484
transform 1 0 77392 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_687
timestamp 1666464484
transform 1 0 78288 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_2
timestamp 1666464484
transform 1 0 1568 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_9
timestamp 1666464484
transform 1 0 2352 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_13
timestamp 1666464484
transform 1 0 2800 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_45
timestamp 1666464484
transform 1 0 6384 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_61
timestamp 1666464484
transform 1 0 8176 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_69
timestamp 1666464484
transform 1 0 9072 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_73
timestamp 1666464484
transform 1 0 9520 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_137
timestamp 1666464484
transform 1 0 16688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_141
timestamp 1666464484
transform 1 0 17136 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_144
timestamp 1666464484
transform 1 0 17472 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_208
timestamp 1666464484
transform 1 0 24640 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1666464484
transform 1 0 25088 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_215
timestamp 1666464484
transform 1 0 25424 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_279
timestamp 1666464484
transform 1 0 32592 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_283
timestamp 1666464484
transform 1 0 33040 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_286
timestamp 1666464484
transform 1 0 33376 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_350
timestamp 1666464484
transform 1 0 40544 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1666464484
transform 1 0 40992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_357
timestamp 1666464484
transform 1 0 41328 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_421
timestamp 1666464484
transform 1 0 48496 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_425
timestamp 1666464484
transform 1 0 48944 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_428
timestamp 1666464484
transform 1 0 49280 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_444
timestamp 1666464484
transform 1 0 51072 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_456
timestamp 1666464484
transform 1 0 52416 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_460
timestamp 1666464484
transform 1 0 52864 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_468
timestamp 1666464484
transform 1 0 53760 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_472
timestamp 1666464484
transform 1 0 54208 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_474
timestamp 1666464484
transform 1 0 54432 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_477
timestamp 1666464484
transform 1 0 54768 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_479
timestamp 1666464484
transform 1 0 54992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_490
timestamp 1666464484
transform 1 0 56224 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_496
timestamp 1666464484
transform 1 0 56896 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_499
timestamp 1666464484
transform 1 0 57232 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_510
timestamp 1666464484
transform 1 0 58464 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_514
timestamp 1666464484
transform 1 0 58912 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_546
timestamp 1666464484
transform 1 0 62496 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_562
timestamp 1666464484
transform 1 0 64288 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_566
timestamp 1666464484
transform 1 0 64736 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_570
timestamp 1666464484
transform 1 0 65184 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_634
timestamp 1666464484
transform 1 0 72352 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_638
timestamp 1666464484
transform 1 0 72800 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_641
timestamp 1666464484
transform 1 0 73136 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_673
timestamp 1666464484
transform 1 0 76720 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_679
timestamp 1666464484
transform 1 0 77392 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_687
timestamp 1666464484
transform 1 0 78288 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_2
timestamp 1666464484
transform 1 0 1568 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_9
timestamp 1666464484
transform 1 0 2352 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_13
timestamp 1666464484
transform 1 0 2800 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_29
timestamp 1666464484
transform 1 0 4592 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_33
timestamp 1666464484
transform 1 0 5040 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_37
timestamp 1666464484
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_101
timestamp 1666464484
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_105
timestamp 1666464484
transform 1 0 13104 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_108
timestamp 1666464484
transform 1 0 13440 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_172
timestamp 1666464484
transform 1 0 20608 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_176
timestamp 1666464484
transform 1 0 21056 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_179
timestamp 1666464484
transform 1 0 21392 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_243
timestamp 1666464484
transform 1 0 28560 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_247
timestamp 1666464484
transform 1 0 29008 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_250
timestamp 1666464484
transform 1 0 29344 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_314
timestamp 1666464484
transform 1 0 36512 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_318
timestamp 1666464484
transform 1 0 36960 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_321
timestamp 1666464484
transform 1 0 37296 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_385
timestamp 1666464484
transform 1 0 44464 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_389
timestamp 1666464484
transform 1 0 44912 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_392
timestamp 1666464484
transform 1 0 45248 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_456
timestamp 1666464484
transform 1 0 52416 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_460
timestamp 1666464484
transform 1 0 52864 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_463
timestamp 1666464484
transform 1 0 53200 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_479
timestamp 1666464484
transform 1 0 54992 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_487
timestamp 1666464484
transform 1 0 55888 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_491
timestamp 1666464484
transform 1 0 56336 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_497
timestamp 1666464484
transform 1 0 57008 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_501
timestamp 1666464484
transform 1 0 57456 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_512
timestamp 1666464484
transform 1 0 58688 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_518
timestamp 1666464484
transform 1 0 59360 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_522
timestamp 1666464484
transform 1 0 59808 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_530
timestamp 1666464484
transform 1 0 60704 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_534
timestamp 1666464484
transform 1 0 61152 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_598
timestamp 1666464484
transform 1 0 68320 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_602
timestamp 1666464484
transform 1 0 68768 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_605
timestamp 1666464484
transform 1 0 69104 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_669
timestamp 1666464484
transform 1 0 76272 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_673
timestamp 1666464484
transform 1 0 76720 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_676
timestamp 1666464484
transform 1 0 77056 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_679
timestamp 1666464484
transform 1 0 77392 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_687
timestamp 1666464484
transform 1 0 78288 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_2
timestamp 1666464484
transform 1 0 1568 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_9
timestamp 1666464484
transform 1 0 2352 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_13
timestamp 1666464484
transform 1 0 2800 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_45
timestamp 1666464484
transform 1 0 6384 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_61
timestamp 1666464484
transform 1 0 8176 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_69
timestamp 1666464484
transform 1 0 9072 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_73
timestamp 1666464484
transform 1 0 9520 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_137
timestamp 1666464484
transform 1 0 16688 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_141
timestamp 1666464484
transform 1 0 17136 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_144
timestamp 1666464484
transform 1 0 17472 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_208
timestamp 1666464484
transform 1 0 24640 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1666464484
transform 1 0 25088 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_215
timestamp 1666464484
transform 1 0 25424 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_279
timestamp 1666464484
transform 1 0 32592 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_283
timestamp 1666464484
transform 1 0 33040 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_286
timestamp 1666464484
transform 1 0 33376 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_350
timestamp 1666464484
transform 1 0 40544 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_354
timestamp 1666464484
transform 1 0 40992 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_357
timestamp 1666464484
transform 1 0 41328 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_421
timestamp 1666464484
transform 1 0 48496 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_425
timestamp 1666464484
transform 1 0 48944 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_428
timestamp 1666464484
transform 1 0 49280 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_460
timestamp 1666464484
transform 1 0 52864 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_476
timestamp 1666464484
transform 1 0 54656 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_482
timestamp 1666464484
transform 1 0 55328 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_486
timestamp 1666464484
transform 1 0 55776 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_494
timestamp 1666464484
transform 1 0 56672 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_496
timestamp 1666464484
transform 1 0 56896 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_499
timestamp 1666464484
transform 1 0 57232 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_510
timestamp 1666464484
transform 1 0 58464 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_522
timestamp 1666464484
transform 1 0 59808 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_538
timestamp 1666464484
transform 1 0 61600 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_550
timestamp 1666464484
transform 1 0 62944 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_554
timestamp 1666464484
transform 1 0 63392 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_562
timestamp 1666464484
transform 1 0 64288 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_566
timestamp 1666464484
transform 1 0 64736 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_570
timestamp 1666464484
transform 1 0 65184 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_634
timestamp 1666464484
transform 1 0 72352 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_638
timestamp 1666464484
transform 1 0 72800 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_641
timestamp 1666464484
transform 1 0 73136 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_673
timestamp 1666464484
transform 1 0 76720 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_679
timestamp 1666464484
transform 1 0 77392 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_687
timestamp 1666464484
transform 1 0 78288 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_2
timestamp 1666464484
transform 1 0 1568 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_9
timestamp 1666464484
transform 1 0 2352 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_13
timestamp 1666464484
transform 1 0 2800 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_17
timestamp 1666464484
transform 1 0 3248 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_33
timestamp 1666464484
transform 1 0 5040 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_37
timestamp 1666464484
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_101
timestamp 1666464484
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_105
timestamp 1666464484
transform 1 0 13104 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_108
timestamp 1666464484
transform 1 0 13440 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_172
timestamp 1666464484
transform 1 0 20608 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_176
timestamp 1666464484
transform 1 0 21056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_179
timestamp 1666464484
transform 1 0 21392 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_243
timestamp 1666464484
transform 1 0 28560 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_247
timestamp 1666464484
transform 1 0 29008 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_250
timestamp 1666464484
transform 1 0 29344 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_314
timestamp 1666464484
transform 1 0 36512 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_318
timestamp 1666464484
transform 1 0 36960 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_321
timestamp 1666464484
transform 1 0 37296 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_385
timestamp 1666464484
transform 1 0 44464 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_389
timestamp 1666464484
transform 1 0 44912 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_392
timestamp 1666464484
transform 1 0 45248 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_456
timestamp 1666464484
transform 1 0 52416 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_460
timestamp 1666464484
transform 1 0 52864 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_463
timestamp 1666464484
transform 1 0 53200 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_479
timestamp 1666464484
transform 1 0 54992 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_487
timestamp 1666464484
transform 1 0 55888 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_492
timestamp 1666464484
transform 1 0 56448 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_496
timestamp 1666464484
transform 1 0 56896 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_502
timestamp 1666464484
transform 1 0 57568 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_506
timestamp 1666464484
transform 1 0 58016 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_508
timestamp 1666464484
transform 1 0 58240 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_513
timestamp 1666464484
transform 1 0 58800 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_515
timestamp 1666464484
transform 1 0 59024 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_520
timestamp 1666464484
transform 1 0 59584 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_524
timestamp 1666464484
transform 1 0 60032 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_528
timestamp 1666464484
transform 1 0 60480 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_534
timestamp 1666464484
transform 1 0 61152 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_598
timestamp 1666464484
transform 1 0 68320 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_602
timestamp 1666464484
transform 1 0 68768 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_605
timestamp 1666464484
transform 1 0 69104 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_669
timestamp 1666464484
transform 1 0 76272 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_673
timestamp 1666464484
transform 1 0 76720 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_676
timestamp 1666464484
transform 1 0 77056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_679
timestamp 1666464484
transform 1 0 77392 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_687
timestamp 1666464484
transform 1 0 78288 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_2
timestamp 1666464484
transform 1 0 1568 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_9
timestamp 1666464484
transform 1 0 2352 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_17
timestamp 1666464484
transform 1 0 3248 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_21
timestamp 1666464484
transform 1 0 3696 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_53
timestamp 1666464484
transform 1 0 7280 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_69
timestamp 1666464484
transform 1 0 9072 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_73
timestamp 1666464484
transform 1 0 9520 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_137
timestamp 1666464484
transform 1 0 16688 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_141
timestamp 1666464484
transform 1 0 17136 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_144
timestamp 1666464484
transform 1 0 17472 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_208
timestamp 1666464484
transform 1 0 24640 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_212
timestamp 1666464484
transform 1 0 25088 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_215
timestamp 1666464484
transform 1 0 25424 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_279
timestamp 1666464484
transform 1 0 32592 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_283
timestamp 1666464484
transform 1 0 33040 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_286
timestamp 1666464484
transform 1 0 33376 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_350
timestamp 1666464484
transform 1 0 40544 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_354
timestamp 1666464484
transform 1 0 40992 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_357
timestamp 1666464484
transform 1 0 41328 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_421
timestamp 1666464484
transform 1 0 48496 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_425
timestamp 1666464484
transform 1 0 48944 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_428
timestamp 1666464484
transform 1 0 49280 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_492
timestamp 1666464484
transform 1 0 56448 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_496
timestamp 1666464484
transform 1 0 56896 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_499
timestamp 1666464484
transform 1 0 57232 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_515
timestamp 1666464484
transform 1 0 59024 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_517
timestamp 1666464484
transform 1 0 59248 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_528
timestamp 1666464484
transform 1 0 60480 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_538
timestamp 1666464484
transform 1 0 61600 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_542
timestamp 1666464484
transform 1 0 62048 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_558
timestamp 1666464484
transform 1 0 63840 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_566
timestamp 1666464484
transform 1 0 64736 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_570
timestamp 1666464484
transform 1 0 65184 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_634
timestamp 1666464484
transform 1 0 72352 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_638
timestamp 1666464484
transform 1 0 72800 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_641
timestamp 1666464484
transform 1 0 73136 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_657
timestamp 1666464484
transform 1 0 74928 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_665
timestamp 1666464484
transform 1 0 75824 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_671
timestamp 1666464484
transform 1 0 76496 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_679
timestamp 1666464484
transform 1 0 77392 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_687
timestamp 1666464484
transform 1 0 78288 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_2
timestamp 1666464484
transform 1 0 1568 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_9
timestamp 1666464484
transform 1 0 2352 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_13
timestamp 1666464484
transform 1 0 2800 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_29
timestamp 1666464484
transform 1 0 4592 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_33
timestamp 1666464484
transform 1 0 5040 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_37
timestamp 1666464484
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_101
timestamp 1666464484
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_105
timestamp 1666464484
transform 1 0 13104 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_108
timestamp 1666464484
transform 1 0 13440 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_172
timestamp 1666464484
transform 1 0 20608 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_176
timestamp 1666464484
transform 1 0 21056 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_179
timestamp 1666464484
transform 1 0 21392 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_243
timestamp 1666464484
transform 1 0 28560 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_247
timestamp 1666464484
transform 1 0 29008 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_250
timestamp 1666464484
transform 1 0 29344 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_314
timestamp 1666464484
transform 1 0 36512 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_318
timestamp 1666464484
transform 1 0 36960 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_321
timestamp 1666464484
transform 1 0 37296 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_385
timestamp 1666464484
transform 1 0 44464 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_389
timestamp 1666464484
transform 1 0 44912 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_392
timestamp 1666464484
transform 1 0 45248 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_456
timestamp 1666464484
transform 1 0 52416 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_460
timestamp 1666464484
transform 1 0 52864 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_463
timestamp 1666464484
transform 1 0 53200 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_495
timestamp 1666464484
transform 1 0 56784 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_503
timestamp 1666464484
transform 1 0 57680 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_507
timestamp 1666464484
transform 1 0 58128 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_515
timestamp 1666464484
transform 1 0 59024 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_519
timestamp 1666464484
transform 1 0 59472 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_531
timestamp 1666464484
transform 1 0 60816 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_534
timestamp 1666464484
transform 1 0 61152 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_539
timestamp 1666464484
transform 1 0 61712 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_543
timestamp 1666464484
transform 1 0 62160 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_575
timestamp 1666464484
transform 1 0 65744 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_579
timestamp 1666464484
transform 1 0 66192 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_585
timestamp 1666464484
transform 1 0 66864 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_589
timestamp 1666464484
transform 1 0 67312 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_597
timestamp 1666464484
transform 1 0 68208 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_601
timestamp 1666464484
transform 1 0 68656 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_605
timestamp 1666464484
transform 1 0 69104 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_669
timestamp 1666464484
transform 1 0 76272 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_673
timestamp 1666464484
transform 1 0 76720 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_676
timestamp 1666464484
transform 1 0 77056 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_679
timestamp 1666464484
transform 1 0 77392 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_687
timestamp 1666464484
transform 1 0 78288 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_2
timestamp 1666464484
transform 1 0 1568 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_9
timestamp 1666464484
transform 1 0 2352 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_13
timestamp 1666464484
transform 1 0 2800 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_45
timestamp 1666464484
transform 1 0 6384 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_61
timestamp 1666464484
transform 1 0 8176 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_69
timestamp 1666464484
transform 1 0 9072 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_73
timestamp 1666464484
transform 1 0 9520 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_137
timestamp 1666464484
transform 1 0 16688 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_141
timestamp 1666464484
transform 1 0 17136 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_144
timestamp 1666464484
transform 1 0 17472 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_208
timestamp 1666464484
transform 1 0 24640 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_212
timestamp 1666464484
transform 1 0 25088 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_215
timestamp 1666464484
transform 1 0 25424 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_279
timestamp 1666464484
transform 1 0 32592 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_283
timestamp 1666464484
transform 1 0 33040 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_286
timestamp 1666464484
transform 1 0 33376 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_350
timestamp 1666464484
transform 1 0 40544 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_354
timestamp 1666464484
transform 1 0 40992 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_357
timestamp 1666464484
transform 1 0 41328 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_421
timestamp 1666464484
transform 1 0 48496 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_425
timestamp 1666464484
transform 1 0 48944 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_428
timestamp 1666464484
transform 1 0 49280 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_492
timestamp 1666464484
transform 1 0 56448 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_496
timestamp 1666464484
transform 1 0 56896 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_499
timestamp 1666464484
transform 1 0 57232 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_504
timestamp 1666464484
transform 1 0 57792 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_508
timestamp 1666464484
transform 1 0 58240 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_512
timestamp 1666464484
transform 1 0 58688 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_515
timestamp 1666464484
transform 1 0 59024 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_523
timestamp 1666464484
transform 1 0 59920 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_537
timestamp 1666464484
transform 1 0 61488 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_549
timestamp 1666464484
transform 1 0 62832 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_553
timestamp 1666464484
transform 1 0 63280 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_561
timestamp 1666464484
transform 1 0 64176 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_567
timestamp 1666464484
transform 1 0 64848 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_570
timestamp 1666464484
transform 1 0 65184 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_573
timestamp 1666464484
transform 1 0 65520 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_637
timestamp 1666464484
transform 1 0 72688 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_641
timestamp 1666464484
transform 1 0 73136 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_673
timestamp 1666464484
transform 1 0 76720 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_679
timestamp 1666464484
transform 1 0 77392 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_687
timestamp 1666464484
transform 1 0 78288 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_2
timestamp 1666464484
transform 1 0 1568 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_9
timestamp 1666464484
transform 1 0 2352 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_13
timestamp 1666464484
transform 1 0 2800 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_29
timestamp 1666464484
transform 1 0 4592 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_33
timestamp 1666464484
transform 1 0 5040 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_37
timestamp 1666464484
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_101
timestamp 1666464484
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_105
timestamp 1666464484
transform 1 0 13104 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_108
timestamp 1666464484
transform 1 0 13440 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_172
timestamp 1666464484
transform 1 0 20608 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_176
timestamp 1666464484
transform 1 0 21056 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_179
timestamp 1666464484
transform 1 0 21392 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_243
timestamp 1666464484
transform 1 0 28560 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_247
timestamp 1666464484
transform 1 0 29008 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_250
timestamp 1666464484
transform 1 0 29344 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_314
timestamp 1666464484
transform 1 0 36512 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_318
timestamp 1666464484
transform 1 0 36960 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_321
timestamp 1666464484
transform 1 0 37296 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_385
timestamp 1666464484
transform 1 0 44464 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_389
timestamp 1666464484
transform 1 0 44912 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_392
timestamp 1666464484
transform 1 0 45248 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_456
timestamp 1666464484
transform 1 0 52416 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_460
timestamp 1666464484
transform 1 0 52864 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_463
timestamp 1666464484
transform 1 0 53200 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_495
timestamp 1666464484
transform 1 0 56784 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_511
timestamp 1666464484
transform 1 0 58576 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_519
timestamp 1666464484
transform 1 0 59472 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_522
timestamp 1666464484
transform 1 0 59808 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_528
timestamp 1666464484
transform 1 0 60480 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_534
timestamp 1666464484
transform 1 0 61152 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_539
timestamp 1666464484
transform 1 0 61712 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_543
timestamp 1666464484
transform 1 0 62160 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_545
timestamp 1666464484
transform 1 0 62384 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_550
timestamp 1666464484
transform 1 0 62944 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_558
timestamp 1666464484
transform 1 0 63840 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_562
timestamp 1666464484
transform 1 0 64288 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_594
timestamp 1666464484
transform 1 0 67872 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_602
timestamp 1666464484
transform 1 0 68768 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_605
timestamp 1666464484
transform 1 0 69104 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_669
timestamp 1666464484
transform 1 0 76272 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_673
timestamp 1666464484
transform 1 0 76720 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_676
timestamp 1666464484
transform 1 0 77056 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_679
timestamp 1666464484
transform 1 0 77392 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_687
timestamp 1666464484
transform 1 0 78288 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_2
timestamp 1666464484
transform 1 0 1568 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_9
timestamp 1666464484
transform 1 0 2352 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_13
timestamp 1666464484
transform 1 0 2800 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_45
timestamp 1666464484
transform 1 0 6384 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_61
timestamp 1666464484
transform 1 0 8176 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_69
timestamp 1666464484
transform 1 0 9072 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_73
timestamp 1666464484
transform 1 0 9520 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_137
timestamp 1666464484
transform 1 0 16688 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_141
timestamp 1666464484
transform 1 0 17136 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_144
timestamp 1666464484
transform 1 0 17472 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_208
timestamp 1666464484
transform 1 0 24640 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_212
timestamp 1666464484
transform 1 0 25088 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_215
timestamp 1666464484
transform 1 0 25424 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_279
timestamp 1666464484
transform 1 0 32592 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_283
timestamp 1666464484
transform 1 0 33040 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_286
timestamp 1666464484
transform 1 0 33376 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_350
timestamp 1666464484
transform 1 0 40544 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_354
timestamp 1666464484
transform 1 0 40992 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_357
timestamp 1666464484
transform 1 0 41328 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_421
timestamp 1666464484
transform 1 0 48496 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_425
timestamp 1666464484
transform 1 0 48944 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_428
timestamp 1666464484
transform 1 0 49280 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_492
timestamp 1666464484
transform 1 0 56448 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_496
timestamp 1666464484
transform 1 0 56896 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_499
timestamp 1666464484
transform 1 0 57232 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_515
timestamp 1666464484
transform 1 0 59024 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_519
timestamp 1666464484
transform 1 0 59472 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_524
timestamp 1666464484
transform 1 0 60032 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_528
timestamp 1666464484
transform 1 0 60480 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_536
timestamp 1666464484
transform 1 0 61376 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_540
timestamp 1666464484
transform 1 0 61824 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_552
timestamp 1666464484
transform 1 0 63168 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_564
timestamp 1666464484
transform 1 0 64512 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_570
timestamp 1666464484
transform 1 0 65184 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_586
timestamp 1666464484
transform 1 0 66976 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_594
timestamp 1666464484
transform 1 0 67872 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_600
timestamp 1666464484
transform 1 0 68544 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_604
timestamp 1666464484
transform 1 0 68992 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_636
timestamp 1666464484
transform 1 0 72576 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_638
timestamp 1666464484
transform 1 0 72800 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_641
timestamp 1666464484
transform 1 0 73136 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_673
timestamp 1666464484
transform 1 0 76720 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_679
timestamp 1666464484
transform 1 0 77392 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_687
timestamp 1666464484
transform 1 0 78288 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_2
timestamp 1666464484
transform 1 0 1568 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_9
timestamp 1666464484
transform 1 0 2352 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_13
timestamp 1666464484
transform 1 0 2800 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_17
timestamp 1666464484
transform 1 0 3248 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_33
timestamp 1666464484
transform 1 0 5040 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_37
timestamp 1666464484
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_101
timestamp 1666464484
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_105
timestamp 1666464484
transform 1 0 13104 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_108
timestamp 1666464484
transform 1 0 13440 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_172
timestamp 1666464484
transform 1 0 20608 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_176
timestamp 1666464484
transform 1 0 21056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_179
timestamp 1666464484
transform 1 0 21392 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_243
timestamp 1666464484
transform 1 0 28560 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_247
timestamp 1666464484
transform 1 0 29008 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_250
timestamp 1666464484
transform 1 0 29344 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_314
timestamp 1666464484
transform 1 0 36512 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_318
timestamp 1666464484
transform 1 0 36960 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_321
timestamp 1666464484
transform 1 0 37296 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_385
timestamp 1666464484
transform 1 0 44464 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_389
timestamp 1666464484
transform 1 0 44912 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_392
timestamp 1666464484
transform 1 0 45248 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_456
timestamp 1666464484
transform 1 0 52416 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_460
timestamp 1666464484
transform 1 0 52864 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_463
timestamp 1666464484
transform 1 0 53200 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_495
timestamp 1666464484
transform 1 0 56784 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_511
timestamp 1666464484
transform 1 0 58576 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_515
timestamp 1666464484
transform 1 0 59024 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_520
timestamp 1666464484
transform 1 0 59584 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_524
timestamp 1666464484
transform 1 0 60032 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_534
timestamp 1666464484
transform 1 0 61152 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_539
timestamp 1666464484
transform 1 0 61712 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_543
timestamp 1666464484
transform 1 0 62160 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_547
timestamp 1666464484
transform 1 0 62608 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_559
timestamp 1666464484
transform 1 0 63952 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_563
timestamp 1666464484
transform 1 0 64400 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_565
timestamp 1666464484
transform 1 0 64624 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_568
timestamp 1666464484
transform 1 0 64960 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_572
timestamp 1666464484
transform 1 0 65408 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_576
timestamp 1666464484
transform 1 0 65856 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_580
timestamp 1666464484
transform 1 0 66304 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_584
timestamp 1666464484
transform 1 0 66752 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_588
timestamp 1666464484
transform 1 0 67200 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_596
timestamp 1666464484
transform 1 0 68096 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_600
timestamp 1666464484
transform 1 0 68544 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_602
timestamp 1666464484
transform 1 0 68768 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_605
timestamp 1666464484
transform 1 0 69104 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_669
timestamp 1666464484
transform 1 0 76272 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_673
timestamp 1666464484
transform 1 0 76720 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_676
timestamp 1666464484
transform 1 0 77056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_679
timestamp 1666464484
transform 1 0 77392 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_687
timestamp 1666464484
transform 1 0 78288 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_2
timestamp 1666464484
transform 1 0 1568 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_9
timestamp 1666464484
transform 1 0 2352 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_17
timestamp 1666464484
transform 1 0 3248 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_21
timestamp 1666464484
transform 1 0 3696 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_77_53
timestamp 1666464484
transform 1 0 7280 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_69
timestamp 1666464484
transform 1 0 9072 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_73
timestamp 1666464484
transform 1 0 9520 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_137
timestamp 1666464484
transform 1 0 16688 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_141
timestamp 1666464484
transform 1 0 17136 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_144
timestamp 1666464484
transform 1 0 17472 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_208
timestamp 1666464484
transform 1 0 24640 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_212
timestamp 1666464484
transform 1 0 25088 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_215
timestamp 1666464484
transform 1 0 25424 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_279
timestamp 1666464484
transform 1 0 32592 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_283
timestamp 1666464484
transform 1 0 33040 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_286
timestamp 1666464484
transform 1 0 33376 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_350
timestamp 1666464484
transform 1 0 40544 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_354
timestamp 1666464484
transform 1 0 40992 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_357
timestamp 1666464484
transform 1 0 41328 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_421
timestamp 1666464484
transform 1 0 48496 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_425
timestamp 1666464484
transform 1 0 48944 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_428
timestamp 1666464484
transform 1 0 49280 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_492
timestamp 1666464484
transform 1 0 56448 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_496
timestamp 1666464484
transform 1 0 56896 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_499
timestamp 1666464484
transform 1 0 57232 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_531
timestamp 1666464484
transform 1 0 60816 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_536
timestamp 1666464484
transform 1 0 61376 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_540
timestamp 1666464484
transform 1 0 61824 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_548
timestamp 1666464484
transform 1 0 62720 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_560
timestamp 1666464484
transform 1 0 64064 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_566
timestamp 1666464484
transform 1 0 64736 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_570
timestamp 1666464484
transform 1 0 65184 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_578
timestamp 1666464484
transform 1 0 66080 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_586
timestamp 1666464484
transform 1 0 66976 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_594
timestamp 1666464484
transform 1 0 67872 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_598
timestamp 1666464484
transform 1 0 68320 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_606
timestamp 1666464484
transform 1 0 69216 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_638
timestamp 1666464484
transform 1 0 72800 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_77_641
timestamp 1666464484
transform 1 0 73136 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_657
timestamp 1666464484
transform 1 0 74928 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_665
timestamp 1666464484
transform 1 0 75824 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_671
timestamp 1666464484
transform 1 0 76496 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_679
timestamp 1666464484
transform 1 0 77392 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_687
timestamp 1666464484
transform 1 0 78288 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_2
timestamp 1666464484
transform 1 0 1568 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_9
timestamp 1666464484
transform 1 0 2352 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_13
timestamp 1666464484
transform 1 0 2800 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_29
timestamp 1666464484
transform 1 0 4592 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_33
timestamp 1666464484
transform 1 0 5040 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_37
timestamp 1666464484
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_101
timestamp 1666464484
transform 1 0 12656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_105
timestamp 1666464484
transform 1 0 13104 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_108
timestamp 1666464484
transform 1 0 13440 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_172
timestamp 1666464484
transform 1 0 20608 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_176
timestamp 1666464484
transform 1 0 21056 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_179
timestamp 1666464484
transform 1 0 21392 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_243
timestamp 1666464484
transform 1 0 28560 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_247
timestamp 1666464484
transform 1 0 29008 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_250
timestamp 1666464484
transform 1 0 29344 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_314
timestamp 1666464484
transform 1 0 36512 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_318
timestamp 1666464484
transform 1 0 36960 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_321
timestamp 1666464484
transform 1 0 37296 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_385
timestamp 1666464484
transform 1 0 44464 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_389
timestamp 1666464484
transform 1 0 44912 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_392
timestamp 1666464484
transform 1 0 45248 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_456
timestamp 1666464484
transform 1 0 52416 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_460
timestamp 1666464484
transform 1 0 52864 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_463
timestamp 1666464484
transform 1 0 53200 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_527
timestamp 1666464484
transform 1 0 60368 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_531
timestamp 1666464484
transform 1 0 60816 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_534
timestamp 1666464484
transform 1 0 61152 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_539
timestamp 1666464484
transform 1 0 61712 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_543
timestamp 1666464484
transform 1 0 62160 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_551
timestamp 1666464484
transform 1 0 63056 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_553
timestamp 1666464484
transform 1 0 63280 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_558
timestamp 1666464484
transform 1 0 63840 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_562
timestamp 1666464484
transform 1 0 64288 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_566
timestamp 1666464484
transform 1 0 64736 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_577
timestamp 1666464484
transform 1 0 65968 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_583
timestamp 1666464484
transform 1 0 66640 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_587
timestamp 1666464484
transform 1 0 67088 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_595
timestamp 1666464484
transform 1 0 67984 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_605
timestamp 1666464484
transform 1 0 69104 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_78_612
timestamp 1666464484
transform 1 0 69888 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_644
timestamp 1666464484
transform 1 0 73472 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_660
timestamp 1666464484
transform 1 0 75264 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_668
timestamp 1666464484
transform 1 0 76160 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_670
timestamp 1666464484
transform 1 0 76384 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_673
timestamp 1666464484
transform 1 0 76720 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_676
timestamp 1666464484
transform 1 0 77056 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_679
timestamp 1666464484
transform 1 0 77392 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_687
timestamp 1666464484
transform 1 0 78288 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_2
timestamp 1666464484
transform 1 0 1568 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_9
timestamp 1666464484
transform 1 0 2352 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_13
timestamp 1666464484
transform 1 0 2800 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_45
timestamp 1666464484
transform 1 0 6384 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_61
timestamp 1666464484
transform 1 0 8176 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_69
timestamp 1666464484
transform 1 0 9072 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_73
timestamp 1666464484
transform 1 0 9520 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_137
timestamp 1666464484
transform 1 0 16688 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_141
timestamp 1666464484
transform 1 0 17136 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_144
timestamp 1666464484
transform 1 0 17472 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_208
timestamp 1666464484
transform 1 0 24640 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_212
timestamp 1666464484
transform 1 0 25088 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_215
timestamp 1666464484
transform 1 0 25424 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_279
timestamp 1666464484
transform 1 0 32592 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_283
timestamp 1666464484
transform 1 0 33040 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_286
timestamp 1666464484
transform 1 0 33376 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_350
timestamp 1666464484
transform 1 0 40544 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_354
timestamp 1666464484
transform 1 0 40992 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_357
timestamp 1666464484
transform 1 0 41328 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_421
timestamp 1666464484
transform 1 0 48496 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_425
timestamp 1666464484
transform 1 0 48944 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_428
timestamp 1666464484
transform 1 0 49280 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_492
timestamp 1666464484
transform 1 0 56448 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_496
timestamp 1666464484
transform 1 0 56896 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_499
timestamp 1666464484
transform 1 0 57232 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_531
timestamp 1666464484
transform 1 0 60816 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_535
timestamp 1666464484
transform 1 0 61264 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_537
timestamp 1666464484
transform 1 0 61488 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_542
timestamp 1666464484
transform 1 0 62048 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_546
timestamp 1666464484
transform 1 0 62496 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_562
timestamp 1666464484
transform 1 0 64288 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_567
timestamp 1666464484
transform 1 0 64848 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_570
timestamp 1666464484
transform 1 0 65184 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_581
timestamp 1666464484
transform 1 0 66416 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_585
timestamp 1666464484
transform 1 0 66864 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_589
timestamp 1666464484
transform 1 0 67312 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_603
timestamp 1666464484
transform 1 0 68880 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_635
timestamp 1666464484
transform 1 0 72464 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_641
timestamp 1666464484
transform 1 0 73136 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_673
timestamp 1666464484
transform 1 0 76720 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_679
timestamp 1666464484
transform 1 0 77392 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_687
timestamp 1666464484
transform 1 0 78288 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_2
timestamp 1666464484
transform 1 0 1568 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_9
timestamp 1666464484
transform 1 0 2352 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_80_13
timestamp 1666464484
transform 1 0 2800 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_29
timestamp 1666464484
transform 1 0 4592 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_33
timestamp 1666464484
transform 1 0 5040 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_37
timestamp 1666464484
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_101
timestamp 1666464484
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_105
timestamp 1666464484
transform 1 0 13104 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_108
timestamp 1666464484
transform 1 0 13440 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_172
timestamp 1666464484
transform 1 0 20608 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_176
timestamp 1666464484
transform 1 0 21056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_179
timestamp 1666464484
transform 1 0 21392 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_243
timestamp 1666464484
transform 1 0 28560 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_247
timestamp 1666464484
transform 1 0 29008 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_250
timestamp 1666464484
transform 1 0 29344 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_314
timestamp 1666464484
transform 1 0 36512 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_318
timestamp 1666464484
transform 1 0 36960 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_321
timestamp 1666464484
transform 1 0 37296 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_385
timestamp 1666464484
transform 1 0 44464 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_389
timestamp 1666464484
transform 1 0 44912 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_392
timestamp 1666464484
transform 1 0 45248 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_456
timestamp 1666464484
transform 1 0 52416 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_460
timestamp 1666464484
transform 1 0 52864 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_463
timestamp 1666464484
transform 1 0 53200 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_527
timestamp 1666464484
transform 1 0 60368 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_531
timestamp 1666464484
transform 1 0 60816 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_534
timestamp 1666464484
transform 1 0 61152 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_538
timestamp 1666464484
transform 1 0 61600 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_542
timestamp 1666464484
transform 1 0 62048 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_548
timestamp 1666464484
transform 1 0 62720 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_556
timestamp 1666464484
transform 1 0 63616 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_560
timestamp 1666464484
transform 1 0 64064 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_564
timestamp 1666464484
transform 1 0 64512 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_566
timestamp 1666464484
transform 1 0 64736 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_569
timestamp 1666464484
transform 1 0 65072 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_571
timestamp 1666464484
transform 1 0 65296 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_582
timestamp 1666464484
transform 1 0 66528 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_588
timestamp 1666464484
transform 1 0 67200 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_600
timestamp 1666464484
transform 1 0 68544 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_602
timestamp 1666464484
transform 1 0 68768 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_605
timestamp 1666464484
transform 1 0 69104 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_669
timestamp 1666464484
transform 1 0 76272 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_673
timestamp 1666464484
transform 1 0 76720 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_676
timestamp 1666464484
transform 1 0 77056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_679
timestamp 1666464484
transform 1 0 77392 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_687
timestamp 1666464484
transform 1 0 78288 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_2
timestamp 1666464484
transform 1 0 1568 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_9
timestamp 1666464484
transform 1 0 2352 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_13
timestamp 1666464484
transform 1 0 2800 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_45
timestamp 1666464484
transform 1 0 6384 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_61
timestamp 1666464484
transform 1 0 8176 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_69
timestamp 1666464484
transform 1 0 9072 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_73
timestamp 1666464484
transform 1 0 9520 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_137
timestamp 1666464484
transform 1 0 16688 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_141
timestamp 1666464484
transform 1 0 17136 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_144
timestamp 1666464484
transform 1 0 17472 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_208
timestamp 1666464484
transform 1 0 24640 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_212
timestamp 1666464484
transform 1 0 25088 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_215
timestamp 1666464484
transform 1 0 25424 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_279
timestamp 1666464484
transform 1 0 32592 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_283
timestamp 1666464484
transform 1 0 33040 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_286
timestamp 1666464484
transform 1 0 33376 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_350
timestamp 1666464484
transform 1 0 40544 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_354
timestamp 1666464484
transform 1 0 40992 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_357
timestamp 1666464484
transform 1 0 41328 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_421
timestamp 1666464484
transform 1 0 48496 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_425
timestamp 1666464484
transform 1 0 48944 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_428
timestamp 1666464484
transform 1 0 49280 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_492
timestamp 1666464484
transform 1 0 56448 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_496
timestamp 1666464484
transform 1 0 56896 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_499
timestamp 1666464484
transform 1 0 57232 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_563
timestamp 1666464484
transform 1 0 64400 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_567
timestamp 1666464484
transform 1 0 64848 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_570
timestamp 1666464484
transform 1 0 65184 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_572
timestamp 1666464484
transform 1 0 65408 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_583
timestamp 1666464484
transform 1 0 66640 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_589
timestamp 1666464484
transform 1 0 67312 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_593
timestamp 1666464484
transform 1 0 67760 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_605
timestamp 1666464484
transform 1 0 69104 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_609
timestamp 1666464484
transform 1 0 69552 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_625
timestamp 1666464484
transform 1 0 71344 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_633
timestamp 1666464484
transform 1 0 72240 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_637
timestamp 1666464484
transform 1 0 72688 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_641
timestamp 1666464484
transform 1 0 73136 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_673
timestamp 1666464484
transform 1 0 76720 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_679
timestamp 1666464484
transform 1 0 77392 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_687
timestamp 1666464484
transform 1 0 78288 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_2
timestamp 1666464484
transform 1 0 1568 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_9
timestamp 1666464484
transform 1 0 2352 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_13
timestamp 1666464484
transform 1 0 2800 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_17
timestamp 1666464484
transform 1 0 3248 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_33
timestamp 1666464484
transform 1 0 5040 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_37
timestamp 1666464484
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_101
timestamp 1666464484
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_105
timestamp 1666464484
transform 1 0 13104 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_108
timestamp 1666464484
transform 1 0 13440 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_172
timestamp 1666464484
transform 1 0 20608 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_176
timestamp 1666464484
transform 1 0 21056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_179
timestamp 1666464484
transform 1 0 21392 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_243
timestamp 1666464484
transform 1 0 28560 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_247
timestamp 1666464484
transform 1 0 29008 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_250
timestamp 1666464484
transform 1 0 29344 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_314
timestamp 1666464484
transform 1 0 36512 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_318
timestamp 1666464484
transform 1 0 36960 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_321
timestamp 1666464484
transform 1 0 37296 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_385
timestamp 1666464484
transform 1 0 44464 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_389
timestamp 1666464484
transform 1 0 44912 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_392
timestamp 1666464484
transform 1 0 45248 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_456
timestamp 1666464484
transform 1 0 52416 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_460
timestamp 1666464484
transform 1 0 52864 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_463
timestamp 1666464484
transform 1 0 53200 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_527
timestamp 1666464484
transform 1 0 60368 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_531
timestamp 1666464484
transform 1 0 60816 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_534
timestamp 1666464484
transform 1 0 61152 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_566
timestamp 1666464484
transform 1 0 64736 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_584
timestamp 1666464484
transform 1 0 66752 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_590
timestamp 1666464484
transform 1 0 67424 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_596
timestamp 1666464484
transform 1 0 68096 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_602
timestamp 1666464484
transform 1 0 68768 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_605
timestamp 1666464484
transform 1 0 69104 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_610
timestamp 1666464484
transform 1 0 69664 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_614
timestamp 1666464484
transform 1 0 70112 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_646
timestamp 1666464484
transform 1 0 73696 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_662
timestamp 1666464484
transform 1 0 75488 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_670
timestamp 1666464484
transform 1 0 76384 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_676
timestamp 1666464484
transform 1 0 77056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_679
timestamp 1666464484
transform 1 0 77392 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_687
timestamp 1666464484
transform 1 0 78288 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_2
timestamp 1666464484
transform 1 0 1568 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_9
timestamp 1666464484
transform 1 0 2352 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_17
timestamp 1666464484
transform 1 0 3248 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_21
timestamp 1666464484
transform 1 0 3696 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_53
timestamp 1666464484
transform 1 0 7280 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_69
timestamp 1666464484
transform 1 0 9072 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_73
timestamp 1666464484
transform 1 0 9520 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_137
timestamp 1666464484
transform 1 0 16688 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_141
timestamp 1666464484
transform 1 0 17136 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_144
timestamp 1666464484
transform 1 0 17472 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_208
timestamp 1666464484
transform 1 0 24640 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_212
timestamp 1666464484
transform 1 0 25088 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_215
timestamp 1666464484
transform 1 0 25424 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_279
timestamp 1666464484
transform 1 0 32592 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_283
timestamp 1666464484
transform 1 0 33040 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_286
timestamp 1666464484
transform 1 0 33376 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_350
timestamp 1666464484
transform 1 0 40544 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_354
timestamp 1666464484
transform 1 0 40992 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_357
timestamp 1666464484
transform 1 0 41328 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_421
timestamp 1666464484
transform 1 0 48496 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_425
timestamp 1666464484
transform 1 0 48944 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_428
timestamp 1666464484
transform 1 0 49280 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_492
timestamp 1666464484
transform 1 0 56448 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_496
timestamp 1666464484
transform 1 0 56896 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_499
timestamp 1666464484
transform 1 0 57232 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_563
timestamp 1666464484
transform 1 0 64400 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_567
timestamp 1666464484
transform 1 0 64848 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_570
timestamp 1666464484
transform 1 0 65184 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_578
timestamp 1666464484
transform 1 0 66080 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_582
timestamp 1666464484
transform 1 0 66528 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_586
timestamp 1666464484
transform 1 0 66976 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_590
timestamp 1666464484
transform 1 0 67424 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_596
timestamp 1666464484
transform 1 0 68096 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_604
timestamp 1666464484
transform 1 0 68992 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_614
timestamp 1666464484
transform 1 0 70112 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_630
timestamp 1666464484
transform 1 0 71904 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_638
timestamp 1666464484
transform 1 0 72800 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_641
timestamp 1666464484
transform 1 0 73136 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_657
timestamp 1666464484
transform 1 0 74928 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_667
timestamp 1666464484
transform 1 0 76048 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_671
timestamp 1666464484
transform 1 0 76496 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_679
timestamp 1666464484
transform 1 0 77392 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_687
timestamp 1666464484
transform 1 0 78288 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_2
timestamp 1666464484
transform 1 0 1568 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_9
timestamp 1666464484
transform 1 0 2352 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_17
timestamp 1666464484
transform 1 0 3248 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_21
timestamp 1666464484
transform 1 0 3696 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_25
timestamp 1666464484
transform 1 0 4144 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_33
timestamp 1666464484
transform 1 0 5040 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_37
timestamp 1666464484
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_101
timestamp 1666464484
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_105
timestamp 1666464484
transform 1 0 13104 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_108
timestamp 1666464484
transform 1 0 13440 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_172
timestamp 1666464484
transform 1 0 20608 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_176
timestamp 1666464484
transform 1 0 21056 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_179
timestamp 1666464484
transform 1 0 21392 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_243
timestamp 1666464484
transform 1 0 28560 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_247
timestamp 1666464484
transform 1 0 29008 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_250
timestamp 1666464484
transform 1 0 29344 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_314
timestamp 1666464484
transform 1 0 36512 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_318
timestamp 1666464484
transform 1 0 36960 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_321
timestamp 1666464484
transform 1 0 37296 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_385
timestamp 1666464484
transform 1 0 44464 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_389
timestamp 1666464484
transform 1 0 44912 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_392
timestamp 1666464484
transform 1 0 45248 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_456
timestamp 1666464484
transform 1 0 52416 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_460
timestamp 1666464484
transform 1 0 52864 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_463
timestamp 1666464484
transform 1 0 53200 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_527
timestamp 1666464484
transform 1 0 60368 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_531
timestamp 1666464484
transform 1 0 60816 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_534
timestamp 1666464484
transform 1 0 61152 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_598
timestamp 1666464484
transform 1 0 68320 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_602
timestamp 1666464484
transform 1 0 68768 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_605
timestamp 1666464484
transform 1 0 69104 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_612
timestamp 1666464484
transform 1 0 69888 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_620
timestamp 1666464484
transform 1 0 70784 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_84_624
timestamp 1666464484
transform 1 0 71232 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_656
timestamp 1666464484
transform 1 0 74816 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_664
timestamp 1666464484
transform 1 0 75712 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_666
timestamp 1666464484
transform 1 0 75936 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_673
timestamp 1666464484
transform 1 0 76720 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_676
timestamp 1666464484
transform 1 0 77056 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_679
timestamp 1666464484
transform 1 0 77392 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_687
timestamp 1666464484
transform 1 0 78288 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_2
timestamp 1666464484
transform 1 0 1568 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_17
timestamp 1666464484
transform 1 0 3248 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_21
timestamp 1666464484
transform 1 0 3696 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_85_53
timestamp 1666464484
transform 1 0 7280 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_69
timestamp 1666464484
transform 1 0 9072 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_73
timestamp 1666464484
transform 1 0 9520 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_137
timestamp 1666464484
transform 1 0 16688 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_141
timestamp 1666464484
transform 1 0 17136 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_144
timestamp 1666464484
transform 1 0 17472 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_208
timestamp 1666464484
transform 1 0 24640 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_212
timestamp 1666464484
transform 1 0 25088 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_215
timestamp 1666464484
transform 1 0 25424 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_279
timestamp 1666464484
transform 1 0 32592 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_283
timestamp 1666464484
transform 1 0 33040 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_286
timestamp 1666464484
transform 1 0 33376 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_350
timestamp 1666464484
transform 1 0 40544 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_354
timestamp 1666464484
transform 1 0 40992 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_357
timestamp 1666464484
transform 1 0 41328 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_421
timestamp 1666464484
transform 1 0 48496 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_425
timestamp 1666464484
transform 1 0 48944 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_428
timestamp 1666464484
transform 1 0 49280 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_492
timestamp 1666464484
transform 1 0 56448 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_496
timestamp 1666464484
transform 1 0 56896 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_499
timestamp 1666464484
transform 1 0 57232 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_563
timestamp 1666464484
transform 1 0 64400 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_567
timestamp 1666464484
transform 1 0 64848 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_570
timestamp 1666464484
transform 1 0 65184 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_602
timestamp 1666464484
transform 1 0 68768 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_606
timestamp 1666464484
transform 1 0 69216 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_609
timestamp 1666464484
transform 1 0 69552 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_617
timestamp 1666464484
transform 1 0 70448 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_619
timestamp 1666464484
transform 1 0 70672 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_626
timestamp 1666464484
transform 1 0 71456 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_630
timestamp 1666464484
transform 1 0 71904 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_638
timestamp 1666464484
transform 1 0 72800 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_641
timestamp 1666464484
transform 1 0 73136 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_687
timestamp 1666464484
transform 1 0 78288 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_2
timestamp 1666464484
transform 1 0 1568 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_17
timestamp 1666464484
transform 1 0 3248 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_21
timestamp 1666464484
transform 1 0 3696 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_29
timestamp 1666464484
transform 1 0 4592 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_33
timestamp 1666464484
transform 1 0 5040 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_37
timestamp 1666464484
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_101
timestamp 1666464484
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_105
timestamp 1666464484
transform 1 0 13104 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_108
timestamp 1666464484
transform 1 0 13440 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_172
timestamp 1666464484
transform 1 0 20608 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_176
timestamp 1666464484
transform 1 0 21056 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_179
timestamp 1666464484
transform 1 0 21392 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_243
timestamp 1666464484
transform 1 0 28560 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_247
timestamp 1666464484
transform 1 0 29008 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_250
timestamp 1666464484
transform 1 0 29344 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_314
timestamp 1666464484
transform 1 0 36512 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_318
timestamp 1666464484
transform 1 0 36960 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_321
timestamp 1666464484
transform 1 0 37296 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_385
timestamp 1666464484
transform 1 0 44464 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_389
timestamp 1666464484
transform 1 0 44912 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_392
timestamp 1666464484
transform 1 0 45248 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_456
timestamp 1666464484
transform 1 0 52416 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_460
timestamp 1666464484
transform 1 0 52864 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_463
timestamp 1666464484
transform 1 0 53200 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_527
timestamp 1666464484
transform 1 0 60368 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_531
timestamp 1666464484
transform 1 0 60816 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_534
timestamp 1666464484
transform 1 0 61152 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_598
timestamp 1666464484
transform 1 0 68320 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_602
timestamp 1666464484
transform 1 0 68768 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_605
timestamp 1666464484
transform 1 0 69104 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_615
timestamp 1666464484
transform 1 0 70224 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_623
timestamp 1666464484
transform 1 0 71120 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_625
timestamp 1666464484
transform 1 0 71344 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_632
timestamp 1666464484
transform 1 0 72128 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_636
timestamp 1666464484
transform 1 0 72576 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_640
timestamp 1666464484
transform 1 0 73024 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_644
timestamp 1666464484
transform 1 0 73472 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_648
timestamp 1666464484
transform 1 0 73920 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_86_654
timestamp 1666464484
transform 1 0 74592 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_670
timestamp 1666464484
transform 1 0 76384 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_676
timestamp 1666464484
transform 1 0 77056 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_684
timestamp 1666464484
transform 1 0 77952 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_687
timestamp 1666464484
transform 1 0 78288 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_2
timestamp 1666464484
transform 1 0 1568 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_17
timestamp 1666464484
transform 1 0 3248 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_21
timestamp 1666464484
transform 1 0 3696 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_87_53
timestamp 1666464484
transform 1 0 7280 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_69
timestamp 1666464484
transform 1 0 9072 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_73
timestamp 1666464484
transform 1 0 9520 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_137
timestamp 1666464484
transform 1 0 16688 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_141
timestamp 1666464484
transform 1 0 17136 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_144
timestamp 1666464484
transform 1 0 17472 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_208
timestamp 1666464484
transform 1 0 24640 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_212
timestamp 1666464484
transform 1 0 25088 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_215
timestamp 1666464484
transform 1 0 25424 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_279
timestamp 1666464484
transform 1 0 32592 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_283
timestamp 1666464484
transform 1 0 33040 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_286
timestamp 1666464484
transform 1 0 33376 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_350
timestamp 1666464484
transform 1 0 40544 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_354
timestamp 1666464484
transform 1 0 40992 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_357
timestamp 1666464484
transform 1 0 41328 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_421
timestamp 1666464484
transform 1 0 48496 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_425
timestamp 1666464484
transform 1 0 48944 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_428
timestamp 1666464484
transform 1 0 49280 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_492
timestamp 1666464484
transform 1 0 56448 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_496
timestamp 1666464484
transform 1 0 56896 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_499
timestamp 1666464484
transform 1 0 57232 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_563
timestamp 1666464484
transform 1 0 64400 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_567
timestamp 1666464484
transform 1 0 64848 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_570
timestamp 1666464484
transform 1 0 65184 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_87_602
timestamp 1666464484
transform 1 0 68768 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_620
timestamp 1666464484
transform 1 0 70784 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_628
timestamp 1666464484
transform 1 0 71680 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_630
timestamp 1666464484
transform 1 0 71904 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_637
timestamp 1666464484
transform 1 0 72688 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_641
timestamp 1666464484
transform 1 0 73136 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_646
timestamp 1666464484
transform 1 0 73696 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_652
timestamp 1666464484
transform 1 0 74368 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_656
timestamp 1666464484
transform 1 0 74816 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_671
timestamp 1666464484
transform 1 0 76496 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_687
timestamp 1666464484
transform 1 0 78288 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_2
timestamp 1666464484
transform 1 0 1568 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_17
timestamp 1666464484
transform 1 0 3248 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_21
timestamp 1666464484
transform 1 0 3696 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_29
timestamp 1666464484
transform 1 0 4592 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_33
timestamp 1666464484
transform 1 0 5040 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_37
timestamp 1666464484
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_101
timestamp 1666464484
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_105
timestamp 1666464484
transform 1 0 13104 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_108
timestamp 1666464484
transform 1 0 13440 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_172
timestamp 1666464484
transform 1 0 20608 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_176
timestamp 1666464484
transform 1 0 21056 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_179
timestamp 1666464484
transform 1 0 21392 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_243
timestamp 1666464484
transform 1 0 28560 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_247
timestamp 1666464484
transform 1 0 29008 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_250
timestamp 1666464484
transform 1 0 29344 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_314
timestamp 1666464484
transform 1 0 36512 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_318
timestamp 1666464484
transform 1 0 36960 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_321
timestamp 1666464484
transform 1 0 37296 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_385
timestamp 1666464484
transform 1 0 44464 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_389
timestamp 1666464484
transform 1 0 44912 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_392
timestamp 1666464484
transform 1 0 45248 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_456
timestamp 1666464484
transform 1 0 52416 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_460
timestamp 1666464484
transform 1 0 52864 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_463
timestamp 1666464484
transform 1 0 53200 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_527
timestamp 1666464484
transform 1 0 60368 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_531
timestamp 1666464484
transform 1 0 60816 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_534
timestamp 1666464484
transform 1 0 61152 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_598
timestamp 1666464484
transform 1 0 68320 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_602
timestamp 1666464484
transform 1 0 68768 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_605
timestamp 1666464484
transform 1 0 69104 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_88_612
timestamp 1666464484
transform 1 0 69888 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_634
timestamp 1666464484
transform 1 0 72352 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_644
timestamp 1666464484
transform 1 0 73472 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_652
timestamp 1666464484
transform 1 0 74368 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_656
timestamp 1666464484
transform 1 0 74816 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_660
timestamp 1666464484
transform 1 0 75264 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_668
timestamp 1666464484
transform 1 0 76160 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_672
timestamp 1666464484
transform 1 0 76608 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_676
timestamp 1666464484
transform 1 0 77056 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_684
timestamp 1666464484
transform 1 0 77952 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_2
timestamp 1666464484
transform 1 0 1568 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_17
timestamp 1666464484
transform 1 0 3248 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_89_21
timestamp 1666464484
transform 1 0 3696 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_53
timestamp 1666464484
transform 1 0 7280 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_69
timestamp 1666464484
transform 1 0 9072 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_73
timestamp 1666464484
transform 1 0 9520 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_137
timestamp 1666464484
transform 1 0 16688 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_141
timestamp 1666464484
transform 1 0 17136 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_144
timestamp 1666464484
transform 1 0 17472 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_208
timestamp 1666464484
transform 1 0 24640 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_212
timestamp 1666464484
transform 1 0 25088 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_215
timestamp 1666464484
transform 1 0 25424 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_279
timestamp 1666464484
transform 1 0 32592 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_283
timestamp 1666464484
transform 1 0 33040 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_286
timestamp 1666464484
transform 1 0 33376 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_350
timestamp 1666464484
transform 1 0 40544 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_354
timestamp 1666464484
transform 1 0 40992 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_357
timestamp 1666464484
transform 1 0 41328 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_421
timestamp 1666464484
transform 1 0 48496 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_425
timestamp 1666464484
transform 1 0 48944 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_428
timestamp 1666464484
transform 1 0 49280 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_492
timestamp 1666464484
transform 1 0 56448 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_496
timestamp 1666464484
transform 1 0 56896 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_499
timestamp 1666464484
transform 1 0 57232 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_563
timestamp 1666464484
transform 1 0 64400 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_567
timestamp 1666464484
transform 1 0 64848 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_89_570
timestamp 1666464484
transform 1 0 65184 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_602
timestamp 1666464484
transform 1 0 68768 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_610
timestamp 1666464484
transform 1 0 69664 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_614
timestamp 1666464484
transform 1 0 70112 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_630
timestamp 1666464484
transform 1 0 71904 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_636
timestamp 1666464484
transform 1 0 72576 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_638
timestamp 1666464484
transform 1 0 72800 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_641
timestamp 1666464484
transform 1 0 73136 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_643
timestamp 1666464484
transform 1 0 73360 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_650
timestamp 1666464484
transform 1 0 74144 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_654
timestamp 1666464484
transform 1 0 74592 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_656
timestamp 1666464484
transform 1 0 74816 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_671
timestamp 1666464484
transform 1 0 76496 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_687
timestamp 1666464484
transform 1 0 78288 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_2
timestamp 1666464484
transform 1 0 1568 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_17
timestamp 1666464484
transform 1 0 3248 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_25
timestamp 1666464484
transform 1 0 4144 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_29
timestamp 1666464484
transform 1 0 4592 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_33
timestamp 1666464484
transform 1 0 5040 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_37
timestamp 1666464484
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_101
timestamp 1666464484
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_105
timestamp 1666464484
transform 1 0 13104 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_108
timestamp 1666464484
transform 1 0 13440 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_172
timestamp 1666464484
transform 1 0 20608 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_176
timestamp 1666464484
transform 1 0 21056 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_179
timestamp 1666464484
transform 1 0 21392 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_243
timestamp 1666464484
transform 1 0 28560 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_247
timestamp 1666464484
transform 1 0 29008 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_250
timestamp 1666464484
transform 1 0 29344 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_314
timestamp 1666464484
transform 1 0 36512 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_318
timestamp 1666464484
transform 1 0 36960 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_321
timestamp 1666464484
transform 1 0 37296 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_385
timestamp 1666464484
transform 1 0 44464 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_389
timestamp 1666464484
transform 1 0 44912 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_392
timestamp 1666464484
transform 1 0 45248 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_456
timestamp 1666464484
transform 1 0 52416 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_460
timestamp 1666464484
transform 1 0 52864 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_463
timestamp 1666464484
transform 1 0 53200 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_527
timestamp 1666464484
transform 1 0 60368 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_531
timestamp 1666464484
transform 1 0 60816 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_534
timestamp 1666464484
transform 1 0 61152 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_598
timestamp 1666464484
transform 1 0 68320 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_602
timestamp 1666464484
transform 1 0 68768 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_605
timestamp 1666464484
transform 1 0 69104 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_637
timestamp 1666464484
transform 1 0 72688 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_641
timestamp 1666464484
transform 1 0 73136 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_90_644
timestamp 1666464484
transform 1 0 73472 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_660
timestamp 1666464484
transform 1 0 75264 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_668
timestamp 1666464484
transform 1 0 76160 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_672
timestamp 1666464484
transform 1 0 76608 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_676
timestamp 1666464484
transform 1 0 77056 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_679
timestamp 1666464484
transform 1 0 77392 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_687
timestamp 1666464484
transform 1 0 78288 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_2
timestamp 1666464484
transform 1 0 1568 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_17
timestamp 1666464484
transform 1 0 3248 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_21
timestamp 1666464484
transform 1 0 3696 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_91_25
timestamp 1666464484
transform 1 0 4144 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_91_57
timestamp 1666464484
transform 1 0 7728 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_65
timestamp 1666464484
transform 1 0 8624 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_69
timestamp 1666464484
transform 1 0 9072 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_73
timestamp 1666464484
transform 1 0 9520 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_137
timestamp 1666464484
transform 1 0 16688 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_141
timestamp 1666464484
transform 1 0 17136 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_144
timestamp 1666464484
transform 1 0 17472 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_208
timestamp 1666464484
transform 1 0 24640 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_212
timestamp 1666464484
transform 1 0 25088 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_215
timestamp 1666464484
transform 1 0 25424 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_279
timestamp 1666464484
transform 1 0 32592 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_283
timestamp 1666464484
transform 1 0 33040 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_286
timestamp 1666464484
transform 1 0 33376 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_350
timestamp 1666464484
transform 1 0 40544 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_354
timestamp 1666464484
transform 1 0 40992 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_357
timestamp 1666464484
transform 1 0 41328 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_421
timestamp 1666464484
transform 1 0 48496 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_425
timestamp 1666464484
transform 1 0 48944 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_428
timestamp 1666464484
transform 1 0 49280 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_492
timestamp 1666464484
transform 1 0 56448 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_496
timestamp 1666464484
transform 1 0 56896 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_499
timestamp 1666464484
transform 1 0 57232 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_563
timestamp 1666464484
transform 1 0 64400 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_567
timestamp 1666464484
transform 1 0 64848 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_570
timestamp 1666464484
transform 1 0 65184 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_634
timestamp 1666464484
transform 1 0 72352 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_638
timestamp 1666464484
transform 1 0 72800 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_641
timestamp 1666464484
transform 1 0 73136 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_671
timestamp 1666464484
transform 1 0 76496 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_687
timestamp 1666464484
transform 1 0 78288 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_92_2
timestamp 1666464484
transform 1 0 1568 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_34
timestamp 1666464484
transform 1 0 5152 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_37
timestamp 1666464484
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_101
timestamp 1666464484
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_105
timestamp 1666464484
transform 1 0 13104 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_108
timestamp 1666464484
transform 1 0 13440 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_172
timestamp 1666464484
transform 1 0 20608 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_176
timestamp 1666464484
transform 1 0 21056 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_179
timestamp 1666464484
transform 1 0 21392 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_243
timestamp 1666464484
transform 1 0 28560 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_247
timestamp 1666464484
transform 1 0 29008 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_250
timestamp 1666464484
transform 1 0 29344 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_314
timestamp 1666464484
transform 1 0 36512 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_318
timestamp 1666464484
transform 1 0 36960 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_321
timestamp 1666464484
transform 1 0 37296 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_385
timestamp 1666464484
transform 1 0 44464 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_389
timestamp 1666464484
transform 1 0 44912 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_392
timestamp 1666464484
transform 1 0 45248 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_456
timestamp 1666464484
transform 1 0 52416 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_460
timestamp 1666464484
transform 1 0 52864 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_463
timestamp 1666464484
transform 1 0 53200 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_527
timestamp 1666464484
transform 1 0 60368 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_531
timestamp 1666464484
transform 1 0 60816 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_534
timestamp 1666464484
transform 1 0 61152 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_598
timestamp 1666464484
transform 1 0 68320 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_602
timestamp 1666464484
transform 1 0 68768 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_605
timestamp 1666464484
transform 1 0 69104 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_669
timestamp 1666464484
transform 1 0 76272 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_673
timestamp 1666464484
transform 1 0 76720 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_676
timestamp 1666464484
transform 1 0 77056 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_684
timestamp 1666464484
transform 1 0 77952 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_2
timestamp 1666464484
transform 1 0 1568 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_34
timestamp 1666464484
transform 1 0 5152 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_37
timestamp 1666464484
transform 1 0 5488 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_69
timestamp 1666464484
transform 1 0 9072 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_72
timestamp 1666464484
transform 1 0 9408 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_104
timestamp 1666464484
transform 1 0 12992 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_107
timestamp 1666464484
transform 1 0 13328 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_139
timestamp 1666464484
transform 1 0 16912 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_142
timestamp 1666464484
transform 1 0 17248 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_174
timestamp 1666464484
transform 1 0 20832 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_177
timestamp 1666464484
transform 1 0 21168 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_209
timestamp 1666464484
transform 1 0 24752 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_212
timestamp 1666464484
transform 1 0 25088 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_244
timestamp 1666464484
transform 1 0 28672 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_247
timestamp 1666464484
transform 1 0 29008 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_279
timestamp 1666464484
transform 1 0 32592 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_282
timestamp 1666464484
transform 1 0 32928 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_314
timestamp 1666464484
transform 1 0 36512 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_317
timestamp 1666464484
transform 1 0 36848 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_349
timestamp 1666464484
transform 1 0 40432 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_352
timestamp 1666464484
transform 1 0 40768 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_384
timestamp 1666464484
transform 1 0 44352 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_387
timestamp 1666464484
transform 1 0 44688 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_419
timestamp 1666464484
transform 1 0 48272 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_422
timestamp 1666464484
transform 1 0 48608 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_454
timestamp 1666464484
transform 1 0 52192 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_457
timestamp 1666464484
transform 1 0 52528 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_489
timestamp 1666464484
transform 1 0 56112 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_492
timestamp 1666464484
transform 1 0 56448 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_524
timestamp 1666464484
transform 1 0 60032 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_527
timestamp 1666464484
transform 1 0 60368 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_559
timestamp 1666464484
transform 1 0 63952 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_562
timestamp 1666464484
transform 1 0 64288 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_594
timestamp 1666464484
transform 1 0 67872 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_597
timestamp 1666464484
transform 1 0 68208 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_629
timestamp 1666464484
transform 1 0 71792 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_632
timestamp 1666464484
transform 1 0 72128 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_664
timestamp 1666464484
transform 1 0 75712 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_93_667
timestamp 1666464484
transform 1 0 76048 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_683
timestamp 1666464484
transform 1 0 77840 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_687
timestamp 1666464484
transform 1 0 78288 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1666464484
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1666464484
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1666464484
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1666464484
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1666464484
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1666464484
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1666464484
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1666464484
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1666464484
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1666464484
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1666464484
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1666464484
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1666464484
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1666464484
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1666464484
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1666464484
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1666464484
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1666464484
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1666464484
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1666464484
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1666464484
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1666464484
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1666464484
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1666464484
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1666464484
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1666464484
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1666464484
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1666464484
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1666464484
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1666464484
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1666464484
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1666464484
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1666464484
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1666464484
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1666464484
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1666464484
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1666464484
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1666464484
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1666464484
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1666464484
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1666464484
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1666464484
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1666464484
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1666464484
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1666464484
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1666464484
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1666464484
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1666464484
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1666464484
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1666464484
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1666464484
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1666464484
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1666464484
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1666464484
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1666464484
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1666464484
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1666464484
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1666464484
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1666464484
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1666464484
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1666464484
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1666464484
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1666464484
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1666464484
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1666464484
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1666464484
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1666464484
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1666464484
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1666464484
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1666464484
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1666464484
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1666464484
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1666464484
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1666464484
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1666464484
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1666464484
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1666464484
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1666464484
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1666464484
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1666464484
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1666464484
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1666464484
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1666464484
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1666464484
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1666464484
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1666464484
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1666464484
transform -1 0 78624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1666464484
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1666464484
transform -1 0 78624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1666464484
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1666464484
transform -1 0 78624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1666464484
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1666464484
transform -1 0 78624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1666464484
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1666464484
transform -1 0 78624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1666464484
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1666464484
transform -1 0 78624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1666464484
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1666464484
transform -1 0 78624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1666464484
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1666464484
transform -1 0 78624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1666464484
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1666464484
transform -1 0 78624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1666464484
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1666464484
transform -1 0 78624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1666464484
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1666464484
transform -1 0 78624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1666464484
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1666464484
transform -1 0 78624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1666464484
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1666464484
transform -1 0 78624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1666464484
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1666464484
transform -1 0 78624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1666464484
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1666464484
transform -1 0 78624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1666464484
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1666464484
transform -1 0 78624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1666464484
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1666464484
transform -1 0 78624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1666464484
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1666464484
transform -1 0 78624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1666464484
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1666464484
transform -1 0 78624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1666464484
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1666464484
transform -1 0 78624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1666464484
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1666464484
transform -1 0 78624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1666464484
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1666464484
transform -1 0 78624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1666464484
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1666464484
transform -1 0 78624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1666464484
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1666464484
transform -1 0 78624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1666464484
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1666464484
transform -1 0 78624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_136
timestamp 1666464484
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_137
timestamp 1666464484
transform -1 0 78624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_138
timestamp 1666464484
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_139
timestamp 1666464484
transform -1 0 78624 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_140
timestamp 1666464484
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_141
timestamp 1666464484
transform -1 0 78624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_142
timestamp 1666464484
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_143
timestamp 1666464484
transform -1 0 78624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_144
timestamp 1666464484
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_145
timestamp 1666464484
transform -1 0 78624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_146
timestamp 1666464484
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_147
timestamp 1666464484
transform -1 0 78624 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_148
timestamp 1666464484
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_149
timestamp 1666464484
transform -1 0 78624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_150
timestamp 1666464484
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_151
timestamp 1666464484
transform -1 0 78624 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_152
timestamp 1666464484
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_153
timestamp 1666464484
transform -1 0 78624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_154
timestamp 1666464484
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_155
timestamp 1666464484
transform -1 0 78624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_156
timestamp 1666464484
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_157
timestamp 1666464484
transform -1 0 78624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_158
timestamp 1666464484
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_159
timestamp 1666464484
transform -1 0 78624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_160
timestamp 1666464484
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_161
timestamp 1666464484
transform -1 0 78624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_162
timestamp 1666464484
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_163
timestamp 1666464484
transform -1 0 78624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_164
timestamp 1666464484
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_165
timestamp 1666464484
transform -1 0 78624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_166
timestamp 1666464484
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_167
timestamp 1666464484
transform -1 0 78624 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_168
timestamp 1666464484
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_169
timestamp 1666464484
transform -1 0 78624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_170
timestamp 1666464484
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_171
timestamp 1666464484
transform -1 0 78624 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_172
timestamp 1666464484
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_173
timestamp 1666464484
transform -1 0 78624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_174
timestamp 1666464484
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_175
timestamp 1666464484
transform -1 0 78624 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_176
timestamp 1666464484
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_177
timestamp 1666464484
transform -1 0 78624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_178
timestamp 1666464484
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_179
timestamp 1666464484
transform -1 0 78624 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_180
timestamp 1666464484
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_181
timestamp 1666464484
transform -1 0 78624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_182
timestamp 1666464484
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_183
timestamp 1666464484
transform -1 0 78624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_184
timestamp 1666464484
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_185
timestamp 1666464484
transform -1 0 78624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_186
timestamp 1666464484
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_187
timestamp 1666464484
transform -1 0 78624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1666464484
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1666464484
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1666464484
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1666464484
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1666464484
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1666464484
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1666464484
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1666464484
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1666464484
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1666464484
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1666464484
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1666464484
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1666464484
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1666464484
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1666464484
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1666464484
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1666464484
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1666464484
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1666464484
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1666464484
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1666464484
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1666464484
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1666464484
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1666464484
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1666464484
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1666464484
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1666464484
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1666464484
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1666464484
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1666464484
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1666464484
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1666464484
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1666464484
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1666464484
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1666464484
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1666464484
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1666464484
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1666464484
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1666464484
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1666464484
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1666464484
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1666464484
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1666464484
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1666464484
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1666464484
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1666464484
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1666464484
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1666464484
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1666464484
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1666464484
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1666464484
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1666464484
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1666464484
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1666464484
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1666464484
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1666464484
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1666464484
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1666464484
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1666464484
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1666464484
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1666464484
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1666464484
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1666464484
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1666464484
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1666464484
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1666464484
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1666464484
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1666464484
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1666464484
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1666464484
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1666464484
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1666464484
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1666464484
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1666464484
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1666464484
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1666464484
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1666464484
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1666464484
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1666464484
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1666464484
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1666464484
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1666464484
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1666464484
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1666464484
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1666464484
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1666464484
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1666464484
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1666464484
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1666464484
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1666464484
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1666464484
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1666464484
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1666464484
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1666464484
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1666464484
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1666464484
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1666464484
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1666464484
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1666464484
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1666464484
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1666464484
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1666464484
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1666464484
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1666464484
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1666464484
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1666464484
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1666464484
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1666464484
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1666464484
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1666464484
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1666464484
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1666464484
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1666464484
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1666464484
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1666464484
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1666464484
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1666464484
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1666464484
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1666464484
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1666464484
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1666464484
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1666464484
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1666464484
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1666464484
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1666464484
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1666464484
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1666464484
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1666464484
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1666464484
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1666464484
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1666464484
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1666464484
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1666464484
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1666464484
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1666464484
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1666464484
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1666464484
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1666464484
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1666464484
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1666464484
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1666464484
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1666464484
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1666464484
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1666464484
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1666464484
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1666464484
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1666464484
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1666464484
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1666464484
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1666464484
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1666464484
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1666464484
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1666464484
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1666464484
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1666464484
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1666464484
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1666464484
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1666464484
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1666464484
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1666464484
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1666464484
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1666464484
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1666464484
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1666464484
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1666464484
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1666464484
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1666464484
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1666464484
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1666464484
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1666464484
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1666464484
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1666464484
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1666464484
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1666464484
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1666464484
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1666464484
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1666464484
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1666464484
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1666464484
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1666464484
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1666464484
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1666464484
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1666464484
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1666464484
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1666464484
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1666464484
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1666464484
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1666464484
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1666464484
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1666464484
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1666464484
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1666464484
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1666464484
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1666464484
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1666464484
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1666464484
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1666464484
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1666464484
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1666464484
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1666464484
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1666464484
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1666464484
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1666464484
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1666464484
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1666464484
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1666464484
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1666464484
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1666464484
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1666464484
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1666464484
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1666464484
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1666464484
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1666464484
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1666464484
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1666464484
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1666464484
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1666464484
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1666464484
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1666464484
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1666464484
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1666464484
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1666464484
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1666464484
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1666464484
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1666464484
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1666464484
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1666464484
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1666464484
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1666464484
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1666464484
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1666464484
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1666464484
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1666464484
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1666464484
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1666464484
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1666464484
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1666464484
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1666464484
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1666464484
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1666464484
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1666464484
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1666464484
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1666464484
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1666464484
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1666464484
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1666464484
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1666464484
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1666464484
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1666464484
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1666464484
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1666464484
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1666464484
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1666464484
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1666464484
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1666464484
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1666464484
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1666464484
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1666464484
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1666464484
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1666464484
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1666464484
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1666464484
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1666464484
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1666464484
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1666464484
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1666464484
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1666464484
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1666464484
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1666464484
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1666464484
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1666464484
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1666464484
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1666464484
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1666464484
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1666464484
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1666464484
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1666464484
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1666464484
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1666464484
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1666464484
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1666464484
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1666464484
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1666464484
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1666464484
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1666464484
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1666464484
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1666464484
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1666464484
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1666464484
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1666464484
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1666464484
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1666464484
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1666464484
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1666464484
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1666464484
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1666464484
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1666464484
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1666464484
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1666464484
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1666464484
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1666464484
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1666464484
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1666464484
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1666464484
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1666464484
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1666464484
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1666464484
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1666464484
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1666464484
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1666464484
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1666464484
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1666464484
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1666464484
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1666464484
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1666464484
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1666464484
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1666464484
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1666464484
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1666464484
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1666464484
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1666464484
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1666464484
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1666464484
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1666464484
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1666464484
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1666464484
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1666464484
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1666464484
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1666464484
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1666464484
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1666464484
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1666464484
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1666464484
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1666464484
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1666464484
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1666464484
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1666464484
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1666464484
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1666464484
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1666464484
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1666464484
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1666464484
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1666464484
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1666464484
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1666464484
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1666464484
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1666464484
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1666464484
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1666464484
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1666464484
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1666464484
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1666464484
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1666464484
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1666464484
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1666464484
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1666464484
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1666464484
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1666464484
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1666464484
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1666464484
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1666464484
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1666464484
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1666464484
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1666464484
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1666464484
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1666464484
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1666464484
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1666464484
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1666464484
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1666464484
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1666464484
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1666464484
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1666464484
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1666464484
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1666464484
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1666464484
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1666464484
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1666464484
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1666464484
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1666464484
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1666464484
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1666464484
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1666464484
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1666464484
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1666464484
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1666464484
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1666464484
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1666464484
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1666464484
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1666464484
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1666464484
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1666464484
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1666464484
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1666464484
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1666464484
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1666464484
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1666464484
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1666464484
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1666464484
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1666464484
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1666464484
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1666464484
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1666464484
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1666464484
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1666464484
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1666464484
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1666464484
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1666464484
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1666464484
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1666464484
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1666464484
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1666464484
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1666464484
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1666464484
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1666464484
transform 1 0 60928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1666464484
transform 1 0 68880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1666464484
transform 1 0 76832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1666464484
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1666464484
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1666464484
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1666464484
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1666464484
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1666464484
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1666464484
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1666464484
transform 1 0 64960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1666464484
transform 1 0 72912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1666464484
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1666464484
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1666464484
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1666464484
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1666464484
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1666464484
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1666464484
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1666464484
transform 1 0 60928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1666464484
transform 1 0 68880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1666464484
transform 1 0 76832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1666464484
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1666464484
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1666464484
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1666464484
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1666464484
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1666464484
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1666464484
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1666464484
transform 1 0 64960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1666464484
transform 1 0 72912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1666464484
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1666464484
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1666464484
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1666464484
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1666464484
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1666464484
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1666464484
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1666464484
transform 1 0 60928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1666464484
transform 1 0 68880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1666464484
transform 1 0 76832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1666464484
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1666464484
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1666464484
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1666464484
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1666464484
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1666464484
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1666464484
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1666464484
transform 1 0 64960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1666464484
transform 1 0 72912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1666464484
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1666464484
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1666464484
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1666464484
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1666464484
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1666464484
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1666464484
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1666464484
transform 1 0 60928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1666464484
transform 1 0 68880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1666464484
transform 1 0 76832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1666464484
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1666464484
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1666464484
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1666464484
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1666464484
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1666464484
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1666464484
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1666464484
transform 1 0 64960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1666464484
transform 1 0 72912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1666464484
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1666464484
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1666464484
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1666464484
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1666464484
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1666464484
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1666464484
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1666464484
transform 1 0 60928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1666464484
transform 1 0 68880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1666464484
transform 1 0 76832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1666464484
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1666464484
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1666464484
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1666464484
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1666464484
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1666464484
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1666464484
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1666464484
transform 1 0 64960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1666464484
transform 1 0 72912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1666464484
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1666464484
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1666464484
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1666464484
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1666464484
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1666464484
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1666464484
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1666464484
transform 1 0 60928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1666464484
transform 1 0 68880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1666464484
transform 1 0 76832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1666464484
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1666464484
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1666464484
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1666464484
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1666464484
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1666464484
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1666464484
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1666464484
transform 1 0 64960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1666464484
transform 1 0 72912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1666464484
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1666464484
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1666464484
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1666464484
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1666464484
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1666464484
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1666464484
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1666464484
transform 1 0 60928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1666464484
transform 1 0 68880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1666464484
transform 1 0 76832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1666464484
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1666464484
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1666464484
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1666464484
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1666464484
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1666464484
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1666464484
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1666464484
transform 1 0 64960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1666464484
transform 1 0 72912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1666464484
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1666464484
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1666464484
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1666464484
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1666464484
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1666464484
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1666464484
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1666464484
transform 1 0 60928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1666464484
transform 1 0 68880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1666464484
transform 1 0 76832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1666464484
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1666464484
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1666464484
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1666464484
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1666464484
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1666464484
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1666464484
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1666464484
transform 1 0 64960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1666464484
transform 1 0 72912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1666464484
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1666464484
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1666464484
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1666464484
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1666464484
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1666464484
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1666464484
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1666464484
transform 1 0 60928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1666464484
transform 1 0 68880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1666464484
transform 1 0 76832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1666464484
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1666464484
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1666464484
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1666464484
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1666464484
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1666464484
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1666464484
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1666464484
transform 1 0 64960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1666464484
transform 1 0 72912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1666464484
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1666464484
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1666464484
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1666464484
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1666464484
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1666464484
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1666464484
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1666464484
transform 1 0 60928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1666464484
transform 1 0 68880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1666464484
transform 1 0 76832 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1666464484
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1666464484
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1666464484
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1666464484
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1666464484
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1666464484
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1666464484
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1666464484
transform 1 0 64960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1666464484
transform 1 0 72912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1666464484
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1666464484
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1666464484
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1666464484
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1666464484
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1666464484
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1666464484
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1666464484
transform 1 0 60928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1666464484
transform 1 0 68880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1666464484
transform 1 0 76832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1666464484
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1666464484
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1666464484
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1666464484
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1666464484
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1666464484
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1666464484
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1666464484
transform 1 0 64960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1666464484
transform 1 0 72912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1666464484
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1666464484
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1666464484
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1666464484
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1666464484
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1666464484
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1666464484
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1666464484
transform 1 0 60928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1666464484
transform 1 0 68880 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1666464484
transform 1 0 76832 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1666464484
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1666464484
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1666464484
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1666464484
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1666464484
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1666464484
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1666464484
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1666464484
transform 1 0 64960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1666464484
transform 1 0 72912 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1666464484
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1666464484
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1666464484
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1666464484
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1666464484
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1666464484
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1666464484
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1666464484
transform 1 0 60928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1666464484
transform 1 0 68880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1666464484
transform 1 0 76832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1666464484
transform 1 0 9296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1666464484
transform 1 0 17248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1666464484
transform 1 0 25200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1666464484
transform 1 0 33152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1666464484
transform 1 0 41104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1666464484
transform 1 0 49056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1666464484
transform 1 0 57008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1666464484
transform 1 0 64960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1666464484
transform 1 0 72912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1666464484
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1666464484
transform 1 0 13216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1666464484
transform 1 0 21168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1666464484
transform 1 0 29120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1666464484
transform 1 0 37072 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1666464484
transform 1 0 45024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1666464484
transform 1 0 52976 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1666464484
transform 1 0 60928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1666464484
transform 1 0 68880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1666464484
transform 1 0 76832 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1666464484
transform 1 0 9296 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1666464484
transform 1 0 17248 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1666464484
transform 1 0 25200 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1666464484
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1666464484
transform 1 0 41104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1666464484
transform 1 0 49056 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1666464484
transform 1 0 57008 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1666464484
transform 1 0 64960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1666464484
transform 1 0 72912 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1666464484
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1666464484
transform 1 0 13216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1666464484
transform 1 0 21168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1666464484
transform 1 0 29120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1666464484
transform 1 0 37072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1666464484
transform 1 0 45024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1666464484
transform 1 0 52976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1666464484
transform 1 0 60928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1666464484
transform 1 0 68880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1666464484
transform 1 0 76832 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1666464484
transform 1 0 9296 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1666464484
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1666464484
transform 1 0 25200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1666464484
transform 1 0 33152 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1666464484
transform 1 0 41104 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1666464484
transform 1 0 49056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1666464484
transform 1 0 57008 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1666464484
transform 1 0 64960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1666464484
transform 1 0 72912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1666464484
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1666464484
transform 1 0 13216 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1666464484
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1666464484
transform 1 0 29120 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1666464484
transform 1 0 37072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1666464484
transform 1 0 45024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1666464484
transform 1 0 52976 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1666464484
transform 1 0 60928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1666464484
transform 1 0 68880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1666464484
transform 1 0 76832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1666464484
transform 1 0 9296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1666464484
transform 1 0 17248 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1666464484
transform 1 0 25200 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1666464484
transform 1 0 33152 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1666464484
transform 1 0 41104 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1666464484
transform 1 0 49056 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1666464484
transform 1 0 57008 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_898
timestamp 1666464484
transform 1 0 64960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_899
timestamp 1666464484
transform 1 0 72912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_900
timestamp 1666464484
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_901
timestamp 1666464484
transform 1 0 13216 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_902
timestamp 1666464484
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_903
timestamp 1666464484
transform 1 0 29120 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_904
timestamp 1666464484
transform 1 0 37072 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_905
timestamp 1666464484
transform 1 0 45024 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_906
timestamp 1666464484
transform 1 0 52976 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_907
timestamp 1666464484
transform 1 0 60928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_908
timestamp 1666464484
transform 1 0 68880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_909
timestamp 1666464484
transform 1 0 76832 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_910
timestamp 1666464484
transform 1 0 9296 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_911
timestamp 1666464484
transform 1 0 17248 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_912
timestamp 1666464484
transform 1 0 25200 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_913
timestamp 1666464484
transform 1 0 33152 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_914
timestamp 1666464484
transform 1 0 41104 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_915
timestamp 1666464484
transform 1 0 49056 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_916
timestamp 1666464484
transform 1 0 57008 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_917
timestamp 1666464484
transform 1 0 64960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_918
timestamp 1666464484
transform 1 0 72912 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_919
timestamp 1666464484
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_920
timestamp 1666464484
transform 1 0 13216 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_921
timestamp 1666464484
transform 1 0 21168 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_922
timestamp 1666464484
transform 1 0 29120 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_923
timestamp 1666464484
transform 1 0 37072 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_924
timestamp 1666464484
transform 1 0 45024 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_925
timestamp 1666464484
transform 1 0 52976 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_926
timestamp 1666464484
transform 1 0 60928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_927
timestamp 1666464484
transform 1 0 68880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_928
timestamp 1666464484
transform 1 0 76832 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_929
timestamp 1666464484
transform 1 0 9296 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_930
timestamp 1666464484
transform 1 0 17248 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_931
timestamp 1666464484
transform 1 0 25200 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_932
timestamp 1666464484
transform 1 0 33152 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_933
timestamp 1666464484
transform 1 0 41104 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_934
timestamp 1666464484
transform 1 0 49056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_935
timestamp 1666464484
transform 1 0 57008 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_936
timestamp 1666464484
transform 1 0 64960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_937
timestamp 1666464484
transform 1 0 72912 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_938
timestamp 1666464484
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_939
timestamp 1666464484
transform 1 0 13216 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_940
timestamp 1666464484
transform 1 0 21168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_941
timestamp 1666464484
transform 1 0 29120 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_942
timestamp 1666464484
transform 1 0 37072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_943
timestamp 1666464484
transform 1 0 45024 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_944
timestamp 1666464484
transform 1 0 52976 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_945
timestamp 1666464484
transform 1 0 60928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_946
timestamp 1666464484
transform 1 0 68880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_947
timestamp 1666464484
transform 1 0 76832 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_948
timestamp 1666464484
transform 1 0 9296 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_949
timestamp 1666464484
transform 1 0 17248 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_950
timestamp 1666464484
transform 1 0 25200 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_951
timestamp 1666464484
transform 1 0 33152 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_952
timestamp 1666464484
transform 1 0 41104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_953
timestamp 1666464484
transform 1 0 49056 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_954
timestamp 1666464484
transform 1 0 57008 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_955
timestamp 1666464484
transform 1 0 64960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_956
timestamp 1666464484
transform 1 0 72912 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_957
timestamp 1666464484
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_958
timestamp 1666464484
transform 1 0 13216 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_959
timestamp 1666464484
transform 1 0 21168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_960
timestamp 1666464484
transform 1 0 29120 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_961
timestamp 1666464484
transform 1 0 37072 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_962
timestamp 1666464484
transform 1 0 45024 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_963
timestamp 1666464484
transform 1 0 52976 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_964
timestamp 1666464484
transform 1 0 60928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_965
timestamp 1666464484
transform 1 0 68880 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_966
timestamp 1666464484
transform 1 0 76832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_967
timestamp 1666464484
transform 1 0 9296 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_968
timestamp 1666464484
transform 1 0 17248 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_969
timestamp 1666464484
transform 1 0 25200 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_970
timestamp 1666464484
transform 1 0 33152 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_971
timestamp 1666464484
transform 1 0 41104 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_972
timestamp 1666464484
transform 1 0 49056 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_973
timestamp 1666464484
transform 1 0 57008 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_974
timestamp 1666464484
transform 1 0 64960 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_975
timestamp 1666464484
transform 1 0 72912 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_976
timestamp 1666464484
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_977
timestamp 1666464484
transform 1 0 13216 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_978
timestamp 1666464484
transform 1 0 21168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_979
timestamp 1666464484
transform 1 0 29120 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_980
timestamp 1666464484
transform 1 0 37072 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_981
timestamp 1666464484
transform 1 0 45024 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_982
timestamp 1666464484
transform 1 0 52976 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_983
timestamp 1666464484
transform 1 0 60928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_984
timestamp 1666464484
transform 1 0 68880 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_985
timestamp 1666464484
transform 1 0 76832 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_986
timestamp 1666464484
transform 1 0 9296 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_987
timestamp 1666464484
transform 1 0 17248 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_988
timestamp 1666464484
transform 1 0 25200 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_989
timestamp 1666464484
transform 1 0 33152 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_990
timestamp 1666464484
transform 1 0 41104 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_991
timestamp 1666464484
transform 1 0 49056 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_992
timestamp 1666464484
transform 1 0 57008 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_993
timestamp 1666464484
transform 1 0 64960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_994
timestamp 1666464484
transform 1 0 72912 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_995
timestamp 1666464484
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_996
timestamp 1666464484
transform 1 0 13216 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_997
timestamp 1666464484
transform 1 0 21168 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_998
timestamp 1666464484
transform 1 0 29120 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_999
timestamp 1666464484
transform 1 0 37072 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1000
timestamp 1666464484
transform 1 0 45024 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1001
timestamp 1666464484
transform 1 0 52976 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1002
timestamp 1666464484
transform 1 0 60928 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1003
timestamp 1666464484
transform 1 0 68880 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1004
timestamp 1666464484
transform 1 0 76832 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1005
timestamp 1666464484
transform 1 0 9296 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1006
timestamp 1666464484
transform 1 0 17248 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1007
timestamp 1666464484
transform 1 0 25200 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1008
timestamp 1666464484
transform 1 0 33152 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1009
timestamp 1666464484
transform 1 0 41104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1010
timestamp 1666464484
transform 1 0 49056 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1011
timestamp 1666464484
transform 1 0 57008 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1012
timestamp 1666464484
transform 1 0 64960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1013
timestamp 1666464484
transform 1 0 72912 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1014
timestamp 1666464484
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1015
timestamp 1666464484
transform 1 0 13216 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1016
timestamp 1666464484
transform 1 0 21168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1017
timestamp 1666464484
transform 1 0 29120 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1018
timestamp 1666464484
transform 1 0 37072 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1019
timestamp 1666464484
transform 1 0 45024 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1020
timestamp 1666464484
transform 1 0 52976 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1021
timestamp 1666464484
transform 1 0 60928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1022
timestamp 1666464484
transform 1 0 68880 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1023
timestamp 1666464484
transform 1 0 76832 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1024
timestamp 1666464484
transform 1 0 9296 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1025
timestamp 1666464484
transform 1 0 17248 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1026
timestamp 1666464484
transform 1 0 25200 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1027
timestamp 1666464484
transform 1 0 33152 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1028
timestamp 1666464484
transform 1 0 41104 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1029
timestamp 1666464484
transform 1 0 49056 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1030
timestamp 1666464484
transform 1 0 57008 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1031
timestamp 1666464484
transform 1 0 64960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1032
timestamp 1666464484
transform 1 0 72912 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1033
timestamp 1666464484
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1034
timestamp 1666464484
transform 1 0 13216 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1035
timestamp 1666464484
transform 1 0 21168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1036
timestamp 1666464484
transform 1 0 29120 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1037
timestamp 1666464484
transform 1 0 37072 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1038
timestamp 1666464484
transform 1 0 45024 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1039
timestamp 1666464484
transform 1 0 52976 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1040
timestamp 1666464484
transform 1 0 60928 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1041
timestamp 1666464484
transform 1 0 68880 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1042
timestamp 1666464484
transform 1 0 76832 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1043
timestamp 1666464484
transform 1 0 9296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1044
timestamp 1666464484
transform 1 0 17248 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1045
timestamp 1666464484
transform 1 0 25200 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1046
timestamp 1666464484
transform 1 0 33152 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1047
timestamp 1666464484
transform 1 0 41104 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1048
timestamp 1666464484
transform 1 0 49056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1049
timestamp 1666464484
transform 1 0 57008 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1050
timestamp 1666464484
transform 1 0 64960 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1051
timestamp 1666464484
transform 1 0 72912 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1052
timestamp 1666464484
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1053
timestamp 1666464484
transform 1 0 13216 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1054
timestamp 1666464484
transform 1 0 21168 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1055
timestamp 1666464484
transform 1 0 29120 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1056
timestamp 1666464484
transform 1 0 37072 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1057
timestamp 1666464484
transform 1 0 45024 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1058
timestamp 1666464484
transform 1 0 52976 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1059
timestamp 1666464484
transform 1 0 60928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1060
timestamp 1666464484
transform 1 0 68880 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1061
timestamp 1666464484
transform 1 0 76832 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1062
timestamp 1666464484
transform 1 0 9296 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1063
timestamp 1666464484
transform 1 0 17248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1064
timestamp 1666464484
transform 1 0 25200 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1065
timestamp 1666464484
transform 1 0 33152 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1066
timestamp 1666464484
transform 1 0 41104 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1067
timestamp 1666464484
transform 1 0 49056 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1068
timestamp 1666464484
transform 1 0 57008 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1069
timestamp 1666464484
transform 1 0 64960 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1070
timestamp 1666464484
transform 1 0 72912 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1071
timestamp 1666464484
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1072
timestamp 1666464484
transform 1 0 13216 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1073
timestamp 1666464484
transform 1 0 21168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1074
timestamp 1666464484
transform 1 0 29120 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1075
timestamp 1666464484
transform 1 0 37072 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1076
timestamp 1666464484
transform 1 0 45024 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1077
timestamp 1666464484
transform 1 0 52976 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1078
timestamp 1666464484
transform 1 0 60928 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1079
timestamp 1666464484
transform 1 0 68880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1080
timestamp 1666464484
transform 1 0 76832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1081
timestamp 1666464484
transform 1 0 5264 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1082
timestamp 1666464484
transform 1 0 9184 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1083
timestamp 1666464484
transform 1 0 13104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1084
timestamp 1666464484
transform 1 0 17024 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1085
timestamp 1666464484
transform 1 0 20944 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1086
timestamp 1666464484
transform 1 0 24864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1087
timestamp 1666464484
transform 1 0 28784 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1088
timestamp 1666464484
transform 1 0 32704 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1089
timestamp 1666464484
transform 1 0 36624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1090
timestamp 1666464484
transform 1 0 40544 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1091
timestamp 1666464484
transform 1 0 44464 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1092
timestamp 1666464484
transform 1 0 48384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1093
timestamp 1666464484
transform 1 0 52304 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1094
timestamp 1666464484
transform 1 0 56224 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1095
timestamp 1666464484
transform 1 0 60144 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1096
timestamp 1666464484
transform 1 0 64064 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1097
timestamp 1666464484
transform 1 0 67984 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1098
timestamp 1666464484
transform 1 0 71904 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1099
timestamp 1666464484
transform 1 0 75824 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _100_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 69216 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _101_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 19936 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _102_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 25648 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _103_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 25536 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _104_
timestamp 1666464484
transform 1 0 18144 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _105_
timestamp 1666464484
transform 1 0 22736 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _106_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 22512 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _107_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 55440 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _108_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 54656 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _109_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 57344 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _110_
timestamp 1666464484
transform 1 0 67312 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _111_
timestamp 1666464484
transform 1 0 68544 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _112_
timestamp 1666464484
transform 1 0 55888 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _113_
timestamp 1666464484
transform 1 0 55440 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _114_
timestamp 1666464484
transform 1 0 57344 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _115_
timestamp 1666464484
transform 1 0 67200 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _116_
timestamp 1666464484
transform 1 0 69216 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _117_
timestamp 1666464484
transform 1 0 69888 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _118_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 70448 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _119_
timestamp 1666464484
transform 1 0 67872 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _120_
timestamp 1666464484
transform 1 0 68656 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _121_
timestamp 1666464484
transform 1 0 69216 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _122_
timestamp 1666464484
transform 1 0 48272 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _123_
timestamp 1666464484
transform -1 0 56672 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _124_
timestamp 1666464484
transform -1 0 53984 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _125_
timestamp 1666464484
transform -1 0 56560 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_
timestamp 1666464484
transform -1 0 51072 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _127_
timestamp 1666464484
transform -1 0 50736 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _128_
timestamp 1666464484
transform -1 0 50064 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _129_
timestamp 1666464484
transform 1 0 47824 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _130_
timestamp 1666464484
transform -1 0 50064 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _131_
timestamp 1666464484
transform 1 0 49392 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _132_
timestamp 1666464484
transform 1 0 46368 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _133_
timestamp 1666464484
transform -1 0 52528 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _134_
timestamp 1666464484
transform -1 0 51856 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _135_
timestamp 1666464484
transform 1 0 49504 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _136_
timestamp 1666464484
transform -1 0 51968 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _137_
timestamp 1666464484
transform -1 0 51296 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _138_
timestamp 1666464484
transform 1 0 48608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _139_
timestamp 1666464484
transform -1 0 53872 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _140_
timestamp 1666464484
transform 1 0 51408 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _141_
timestamp 1666464484
transform -1 0 59472 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _142_
timestamp 1666464484
transform -1 0 52752 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _143_
timestamp 1666464484
transform 1 0 46816 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _144_
timestamp 1666464484
transform -1 0 60592 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _145_
timestamp 1666464484
transform -1 0 52864 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _146_
timestamp 1666464484
transform 1 0 48160 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _147_
timestamp 1666464484
transform -1 0 56896 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _148_
timestamp 1666464484
transform -1 0 53536 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _149_
timestamp 1666464484
transform 1 0 50064 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _150_
timestamp 1666464484
transform 1 0 53312 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _151_
timestamp 1666464484
transform 1 0 53760 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _152_
timestamp 1666464484
transform 1 0 51968 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _153_
timestamp 1666464484
transform -1 0 56112 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _154_
timestamp 1666464484
transform 1 0 53872 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _155_
timestamp 1666464484
transform 1 0 53648 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _156_
timestamp 1666464484
transform 1 0 54096 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _157_
timestamp 1666464484
transform 1 0 52640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _158_
timestamp 1666464484
transform -1 0 56112 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _159_
timestamp 1666464484
transform -1 0 55440 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _160_
timestamp 1666464484
transform 1 0 50176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _161_
timestamp 1666464484
transform -1 0 56784 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _162_
timestamp 1666464484
transform -1 0 56000 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _163_
timestamp 1666464484
transform 1 0 51968 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _164_
timestamp 1666464484
transform -1 0 56896 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _165_
timestamp 1666464484
transform -1 0 56224 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _166_
timestamp 1666464484
transform 1 0 56560 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _167_
timestamp 1666464484
transform 1 0 57344 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _168_
timestamp 1666464484
transform 1 0 56784 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _169_
timestamp 1666464484
transform -1 0 59360 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _170_
timestamp 1666464484
transform -1 0 58464 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _171_
timestamp 1666464484
transform 1 0 54880 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _172_
timestamp 1666464484
transform -1 0 62944 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _173_
timestamp 1666464484
transform -1 0 58464 0 -1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _174_
timestamp 1666464484
transform 1 0 56000 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _175_
timestamp 1666464484
transform -1 0 59584 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _176_
timestamp 1666464484
transform -1 0 58688 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _177_
timestamp 1666464484
transform 1 0 57120 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _178_
timestamp 1666464484
transform 1 0 58352 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _179_
timestamp 1666464484
transform 1 0 58688 0 -1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _180_
timestamp 1666464484
transform 1 0 58576 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _181_
timestamp 1666464484
transform -1 0 61600 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _182_
timestamp 1666464484
transform 1 0 59248 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _183_
timestamp 1666464484
transform -1 0 61712 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _184_
timestamp 1666464484
transform -1 0 60480 0 -1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _185_
timestamp 1666464484
transform 1 0 57232 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _186_
timestamp 1666464484
transform -1 0 66864 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _187_
timestamp 1666464484
transform -1 0 60816 0 1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _188_
timestamp 1666464484
transform 1 0 57344 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _189_
timestamp 1666464484
transform -1 0 64848 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _190_
timestamp 1666464484
transform -1 0 61488 0 -1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _191_
timestamp 1666464484
transform 1 0 60032 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _192_
timestamp 1666464484
transform 1 0 61264 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _193_
timestamp 1666464484
transform 1 0 61712 0 -1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _194_
timestamp 1666464484
transform 1 0 61264 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _195_
timestamp 1666464484
transform -1 0 63840 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _196_
timestamp 1666464484
transform 1 0 62048 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _197_
timestamp 1666464484
transform -1 0 62944 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _198_
timestamp 1666464484
transform 1 0 62048 0 -1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _199_
timestamp 1666464484
transform 1 0 59584 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _200_
timestamp 1666464484
transform -1 0 68544 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _201_
timestamp 1666464484
transform -1 0 64512 0 -1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _202_
timestamp 1666464484
transform 1 0 59136 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _203_
timestamp 1666464484
transform -1 0 64736 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _204_
timestamp 1666464484
transform -1 0 63952 0 1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _205_
timestamp 1666464484
transform 1 0 60928 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _206_
timestamp 1666464484
transform 1 0 63392 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _207_
timestamp 1666464484
transform -1 0 64064 0 -1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _208_
timestamp 1666464484
transform 1 0 61264 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _209_
timestamp 1666464484
transform -1 0 66976 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _210_
timestamp 1666464484
transform 1 0 65408 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _211_
timestamp 1666464484
transform -1 0 66640 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _212_
timestamp 1666464484
transform -1 0 65968 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _213_
timestamp 1666464484
transform 1 0 61600 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _214_
timestamp 1666464484
transform 1 0 64400 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _215_
timestamp 1666464484
transform 1 0 65296 0 -1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _216_
timestamp 1666464484
transform 1 0 62272 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _217_
timestamp 1666464484
transform -1 0 67200 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _218_
timestamp 1666464484
transform -1 0 66528 0 1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _219_
timestamp 1666464484
transform 1 0 63168 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _220_
timestamp 1666464484
transform -1 0 67312 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _221_
timestamp 1666464484
transform -1 0 66640 0 -1 67424
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _222_
timestamp 1666464484
transform 1 0 66976 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _223_
timestamp 1666464484
transform -1 0 68768 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _224_
timestamp 1666464484
transform -1 0 68544 0 1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _225_
timestamp 1666464484
transform 1 0 67648 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _226_
timestamp 1666464484
transform -1 0 69664 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _227_
timestamp 1666464484
transform -1 0 68880 0 -1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _228_
timestamp 1666464484
transform 1 0 67648 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _229_
timestamp 1666464484
transform 1 0 68544 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _230_
timestamp 1666464484
transform -1 0 69104 0 -1 67424
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _231_
timestamp 1666464484
transform -1 0 73696 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _232_
timestamp 1666464484
transform -1 0 74368 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _233_
timestamp 1666464484
transform -1 0 74368 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _234_
timestamp 1666464484
transform 1 0 73472 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _235_
timestamp 1666464484
transform 1 0 69216 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _236_
timestamp 1666464484
transform 1 0 68992 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _237_
timestamp 1666464484
transform 1 0 5600 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _238_
timestamp 1666464484
transform 1 0 6272 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _239_
timestamp 1666464484
transform 1 0 6720 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _240_
timestamp 1666464484
transform 1 0 7616 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _241_
timestamp 1666464484
transform 1 0 8288 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _242_
timestamp 1666464484
transform 1 0 8960 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _243_
timestamp 1666464484
transform 1 0 9744 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _244_
timestamp 1666464484
transform 1 0 10416 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _245_
timestamp 1666464484
transform 1 0 10976 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _246_
timestamp 1666464484
transform 1 0 11536 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _247_
timestamp 1666464484
transform 1 0 12432 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _248_
timestamp 1666464484
transform 1 0 13104 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _249_
timestamp 1666464484
transform 1 0 57344 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _250_
timestamp 1666464484
transform 1 0 55104 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _251_
timestamp 1666464484
transform 1 0 55664 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _252_
timestamp 1666464484
transform 1 0 55440 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _253_
timestamp 1666464484
transform 1 0 19488 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _254_
timestamp 1666464484
transform 1 0 19376 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _255_
timestamp 1666464484
transform 1 0 18144 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _256_
timestamp 1666464484
transform 1 0 18480 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _257_
timestamp 1666464484
transform 1 0 20608 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _258_
timestamp 1666464484
transform 1 0 21504 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _259_
timestamp 1666464484
transform 1 0 20272 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _260_
timestamp 1666464484
transform 1 0 20720 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _261_
timestamp 1666464484
transform 1 0 23072 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _262_
timestamp 1666464484
transform 1 0 23520 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _263_
timestamp 1666464484
transform 1 0 22848 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _264_
timestamp 1666464484
transform 1 0 23408 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _265_
timestamp 1666464484
transform 1 0 26208 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _266_
timestamp 1666464484
transform 1 0 25312 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _267_
timestamp 1666464484
transform 1 0 25648 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _268_
timestamp 1666464484
transform 1 0 26208 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _269_
timestamp 1666464484
transform -1 0 5152 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _270_
timestamp 1666464484
transform -1 0 5824 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _271_
timestamp 1666464484
transform -1 0 6496 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _272_
timestamp 1666464484
transform -1 0 7056 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _273_
timestamp 1666464484
transform -1 0 7952 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _274_
timestamp 1666464484
transform -1 0 8512 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _275_
timestamp 1666464484
transform -1 0 9184 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _276_
timestamp 1666464484
transform -1 0 9968 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _277_
timestamp 1666464484
transform -1 0 10640 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _278_
timestamp 1666464484
transform -1 0 11312 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _279_
timestamp 1666464484
transform -1 0 11872 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _280_
timestamp 1666464484
transform -1 0 12768 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _281_
timestamp 1666464484
transform -1 0 12992 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _282_
timestamp 1666464484
transform -1 0 13888 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _283_
timestamp 1666464484
transform -1 0 14560 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _284_
timestamp 1666464484
transform -1 0 15232 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _285_
timestamp 1666464484
transform -1 0 16240 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _286_
timestamp 1666464484
transform -1 0 16240 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _287_
timestamp 1666464484
transform -1 0 17136 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _288_
timestamp 1666464484
transform -1 0 18256 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _289_
timestamp 1666464484
transform -1 0 19152 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _290_
timestamp 1666464484
transform -1 0 19152 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _291_
timestamp 1666464484
transform -1 0 20048 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _292_
timestamp 1666464484
transform -1 0 20496 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _293_
timestamp 1666464484
transform -1 0 22176 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _294_
timestamp 1666464484
transform -1 0 22176 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _295_
timestamp 1666464484
transform -1 0 22624 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _296_
timestamp 1666464484
transform -1 0 22960 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _297_
timestamp 1666464484
transform -1 0 24192 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _298_
timestamp 1666464484
transform -1 0 24640 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _299_
timestamp 1666464484
transform -1 0 24864 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _300_
timestamp 1666464484
transform -1 0 25760 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _301_
timestamp 1666464484
transform 1 0 27216 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _302_
timestamp 1666464484
transform 1 0 27888 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _303_
timestamp 1666464484
transform 1 0 28448 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _304_
timestamp 1666464484
transform 1 0 29456 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _305_
timestamp 1666464484
transform 1 0 30352 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _306_
timestamp 1666464484
transform 1 0 30240 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _307_
timestamp 1666464484
transform 1 0 31136 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _308_
timestamp 1666464484
transform 1 0 31808 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _309_
timestamp 1666464484
transform 1 0 32480 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _310_
timestamp 1666464484
transform 1 0 33488 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _311_
timestamp 1666464484
transform 1 0 33936 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _312_
timestamp 1666464484
transform 1 0 34608 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _313_
timestamp 1666464484
transform 1 0 34944 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _314_
timestamp 1666464484
transform 1 0 35840 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _315_
timestamp 1666464484
transform 1 0 36512 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _316_
timestamp 1666464484
transform 1 0 37408 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _317_
timestamp 1666464484
transform 1 0 37856 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _318_
timestamp 1666464484
transform 1 0 38528 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _319_
timestamp 1666464484
transform 1 0 39312 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _320_
timestamp 1666464484
transform 1 0 39536 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _321_
timestamp 1666464484
transform 1 0 40432 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _322_
timestamp 1666464484
transform 1 0 41440 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _323_
timestamp 1666464484
transform 1 0 41888 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _324_
timestamp 1666464484
transform 1 0 42560 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _325_
timestamp 1666464484
transform 1 0 43232 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _326_
timestamp 1666464484
transform 1 0 43904 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _327_
timestamp 1666464484
transform 1 0 45360 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _328_
timestamp 1666464484
transform 1 0 46256 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _329_
timestamp 1666464484
transform 1 0 46032 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _330_
timestamp 1666464484
transform 1 0 46704 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _331_
timestamp 1666464484
transform 1 0 47376 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _332_
timestamp 1666464484
transform 1 0 48048 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _333_
timestamp 1666464484
transform -1 0 26768 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _334_
timestamp 1666464484
transform -1 0 27440 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _335_
timestamp 1666464484
transform -1 0 28112 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _336_
timestamp 1666464484
transform -1 0 28784 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _337_
timestamp 1666464484
transform -1 0 29232 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _338_
timestamp 1666464484
transform -1 0 30128 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _339_
timestamp 1666464484
transform -1 0 30576 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _340_
timestamp 1666464484
transform -1 0 31472 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _341_
timestamp 1666464484
transform -1 0 32144 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _342_
timestamp 1666464484
transform -1 0 32704 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _343_
timestamp 1666464484
transform -1 0 33488 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _344_
timestamp 1666464484
transform -1 0 34160 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _345_
timestamp 1666464484
transform -1 0 34720 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _346_
timestamp 1666464484
transform -1 0 35168 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _347_
timestamp 1666464484
transform -1 0 36064 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _348_
timestamp 1666464484
transform -1 0 36848 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _349_
timestamp 1666464484
transform -1 0 37520 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _350_
timestamp 1666464484
transform -1 0 38192 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _351_
timestamp 1666464484
transform -1 0 38864 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _352_
timestamp 1666464484
transform -1 0 39312 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _353_
timestamp 1666464484
transform -1 0 39872 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _354_
timestamp 1666464484
transform -1 0 40768 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _355_
timestamp 1666464484
transform -1 0 41552 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _356_
timestamp 1666464484
transform -1 0 42224 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _357_
timestamp 1666464484
transform -1 0 42896 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _358_
timestamp 1666464484
transform -1 0 43456 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _359_
timestamp 1666464484
transform -1 0 44240 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _360_
timestamp 1666464484
transform -1 0 44912 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _361_
timestamp 1666464484
transform -1 0 45808 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _362_
timestamp 1666464484
transform -1 0 46368 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _363_
timestamp 1666464484
transform -1 0 47040 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _364_
timestamp 1666464484
transform -1 0 47712 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _365_
timestamp 1666464484
transform 1 0 70784 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _366_
timestamp 1666464484
transform 1 0 71456 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _367_
timestamp 1666464484
transform 1 0 72016 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _368_
timestamp 1666464484
transform 1 0 72800 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _369_
timestamp 1666464484
transform -1 0 70448 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _370_
timestamp 1666464484
transform -1 0 71120 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _371_
timestamp 1666464484
transform -1 0 71680 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _372_
timestamp 1666464484
transform -1 0 72352 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _373_
timestamp 1666464484
transform 1 0 70112 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _374_
timestamp 1666464484
transform -1 0 69888 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1666464484
transform -1 0 78288 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1666464484
transform 1 0 3472 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1666464484
transform 1 0 5376 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1666464484
transform -1 0 12096 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1666464484
transform 1 0 12320 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1666464484
transform 1 0 13440 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1666464484
transform -1 0 14224 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1666464484
transform 1 0 14448 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1666464484
transform 1 0 15456 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1666464484
transform 1 0 15344 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1666464484
transform -1 0 16912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1666464484
transform 1 0 17584 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1666464484
transform -1 0 18144 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1666464484
transform 1 0 5712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1666464484
transform 1 0 18368 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1666464484
transform 1 0 19264 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1666464484
transform 1 0 20160 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1666464484
transform -1 0 20832 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1666464484
transform 1 0 21504 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1666464484
transform 1 0 21392 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1666464484
transform -1 0 22960 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1666464484
transform 1 0 23184 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1666464484
transform 1 0 24192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1666464484
transform -1 0 24752 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1666464484
transform -1 0 7392 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1666464484
transform -1 0 25984 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1666464484
transform 1 0 26208 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1666464484
transform -1 0 7280 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1666464484
transform -1 0 8176 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1666464484
transform -1 0 10304 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1666464484
transform 1 0 8400 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1666464484
transform -1 0 10304 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1666464484
transform 1 0 10528 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1666464484
transform 1 0 11424 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1666464484
transform -1 0 75712 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1666464484
transform -1 0 78288 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1666464484
transform -1 0 78288 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1666464484
transform -1 0 78288 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1666464484
transform -1 0 78288 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1666464484
transform -1 0 78288 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1666464484
transform -1 0 78288 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1666464484
transform -1 0 78288 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1666464484
transform -1 0 77392 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1666464484
transform -1 0 78288 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1666464484
transform -1 0 78288 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1666464484
transform -1 0 78288 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1666464484
transform -1 0 78288 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1666464484
transform -1 0 78288 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1666464484
transform -1 0 78288 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1666464484
transform -1 0 78288 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1666464484
transform -1 0 77392 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1666464484
transform -1 0 78288 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1666464484
transform -1 0 78288 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1666464484
transform -1 0 78288 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1666464484
transform -1 0 78288 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1666464484
transform -1 0 78288 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1666464484
transform -1 0 78288 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1666464484
transform -1 0 78288 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1666464484
transform -1 0 77392 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1666464484
transform -1 0 76720 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1666464484
transform -1 0 78288 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1666464484
transform -1 0 78288 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input63
timestamp 1666464484
transform -1 0 78288 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1666464484
transform -1 0 78288 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input65
timestamp 1666464484
transform -1 0 78288 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input66
timestamp 1666464484
transform -1 0 78288 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input67
timestamp 1666464484
transform -1 0 77392 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input68
timestamp 1666464484
transform 1 0 1680 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input69
timestamp 1666464484
transform 1 0 1680 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input70
timestamp 1666464484
transform 1 0 1680 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input71
timestamp 1666464484
transform 1 0 1680 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input72
timestamp 1666464484
transform 1 0 1680 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input73
timestamp 1666464484
transform 1 0 1680 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1666464484
transform 1 0 1680 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1666464484
transform 1 0 2576 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input76
timestamp 1666464484
transform 1 0 1680 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input77
timestamp 1666464484
transform 1 0 1680 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input78
timestamp 1666464484
transform 1 0 1680 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input79
timestamp 1666464484
transform 1 0 1680 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input80
timestamp 1666464484
transform 1 0 1680 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input81
timestamp 1666464484
transform 1 0 1680 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input82
timestamp 1666464484
transform 1 0 1680 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input83
timestamp 1666464484
transform 1 0 2576 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input84
timestamp 1666464484
transform 1 0 1680 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input85
timestamp 1666464484
transform 1 0 1680 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input86
timestamp 1666464484
transform 1 0 1680 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input87
timestamp 1666464484
transform 1 0 1680 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input88
timestamp 1666464484
transform 1 0 1680 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input89
timestamp 1666464484
transform 1 0 1680 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input90
timestamp 1666464484
transform 1 0 2576 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input91
timestamp 1666464484
transform 1 0 2576 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input92
timestamp 1666464484
transform 1 0 2576 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input93
timestamp 1666464484
transform 1 0 1680 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input94
timestamp 1666464484
transform 1 0 1680 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input95
timestamp 1666464484
transform 1 0 1680 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input96
timestamp 1666464484
transform 1 0 1680 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input97
timestamp 1666464484
transform 1 0 1680 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input98
timestamp 1666464484
transform 1 0 1680 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input99
timestamp 1666464484
transform 1 0 2576 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input100
timestamp 1666464484
transform -1 0 26880 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input101
timestamp 1666464484
transform -1 0 33824 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input102
timestamp 1666464484
transform 1 0 34048 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input103
timestamp 1666464484
transform 1 0 34944 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input104
timestamp 1666464484
transform -1 0 35616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input105
timestamp 1666464484
transform -1 0 36512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input106
timestamp 1666464484
transform 1 0 36960 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input107
timestamp 1666464484
transform -1 0 37744 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input108
timestamp 1666464484
transform 1 0 37968 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input109
timestamp 1666464484
transform 1 0 38976 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input110
timestamp 1666464484
transform -1 0 39536 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input111
timestamp 1666464484
transform -1 0 27776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input112
timestamp 1666464484
transform -1 0 40432 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input113
timestamp 1666464484
transform 1 0 41440 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input114
timestamp 1666464484
transform 1 0 41664 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input115
timestamp 1666464484
transform 1 0 42560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input116
timestamp 1666464484
transform 1 0 43456 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input117
timestamp 1666464484
transform 1 0 43680 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input118
timestamp 1666464484
transform 1 0 44800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input119
timestamp 1666464484
transform 1 0 45696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input120
timestamp 1666464484
transform -1 0 47264 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input121
timestamp 1666464484
transform 1 0 46368 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input122
timestamp 1666464484
transform 1 0 28000 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input123
timestamp 1666464484
transform -1 0 48160 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input124
timestamp 1666464484
transform 1 0 47712 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input125
timestamp 1666464484
transform 1 0 28896 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input126
timestamp 1666464484
transform -1 0 29904 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input127
timestamp 1666464484
transform 1 0 30240 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input128
timestamp 1666464484
transform -1 0 30800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input129
timestamp 1666464484
transform -1 0 31696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input130
timestamp 1666464484
transform 1 0 32256 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input131
timestamp 1666464484
transform -1 0 32592 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input132
timestamp 1666464484
transform -1 0 72912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input133
timestamp 1666464484
transform -1 0 72240 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input134
timestamp 1666464484
transform 1 0 71904 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input135
timestamp 1666464484
transform 1 0 73248 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input136
timestamp 1666464484
transform -1 0 74816 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input137
timestamp 1666464484
transform 1 0 70672 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output138 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 73920 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output139
timestamp 1666464484
transform 1 0 74928 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output140
timestamp 1666464484
transform 1 0 74928 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output141
timestamp 1666464484
transform 1 0 76720 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output142
timestamp 1666464484
transform 1 0 74928 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output143
timestamp 1666464484
transform 1 0 76720 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output144
timestamp 1666464484
transform 1 0 74928 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output145
timestamp 1666464484
transform 1 0 75152 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output146
timestamp 1666464484
transform 1 0 76720 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output147
timestamp 1666464484
transform 1 0 74928 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output148
timestamp 1666464484
transform 1 0 76720 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output149
timestamp 1666464484
transform 1 0 74928 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output150
timestamp 1666464484
transform 1 0 75152 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output151
timestamp 1666464484
transform 1 0 76720 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output152
timestamp 1666464484
transform 1 0 74928 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output153
timestamp 1666464484
transform 1 0 75152 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output154
timestamp 1666464484
transform 1 0 76720 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output155
timestamp 1666464484
transform 1 0 74928 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output156
timestamp 1666464484
transform 1 0 76720 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output157
timestamp 1666464484
transform 1 0 74928 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output158
timestamp 1666464484
transform 1 0 76720 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output159
timestamp 1666464484
transform 1 0 74928 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output160
timestamp 1666464484
transform 1 0 75152 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output161
timestamp 1666464484
transform 1 0 76720 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output162
timestamp 1666464484
transform 1 0 76720 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output163
timestamp 1666464484
transform 1 0 74928 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output164
timestamp 1666464484
transform 1 0 74928 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output165
timestamp 1666464484
transform 1 0 76720 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output166
timestamp 1666464484
transform 1 0 74928 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output167
timestamp 1666464484
transform 1 0 76720 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output168
timestamp 1666464484
transform 1 0 74928 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output169
timestamp 1666464484
transform 1 0 75152 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output170
timestamp 1666464484
transform 1 0 76720 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output171
timestamp 1666464484
transform -1 0 3248 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output172
timestamp 1666464484
transform -1 0 3248 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output173
timestamp 1666464484
transform -1 0 3248 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output174
timestamp 1666464484
transform -1 0 3248 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output175
timestamp 1666464484
transform -1 0 3248 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output176
timestamp 1666464484
transform -1 0 3248 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output177
timestamp 1666464484
transform -1 0 3248 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output178
timestamp 1666464484
transform -1 0 5040 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output179
timestamp 1666464484
transform -1 0 3248 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output180
timestamp 1666464484
transform -1 0 3248 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output181
timestamp 1666464484
transform -1 0 3248 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output182
timestamp 1666464484
transform -1 0 3248 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output183
timestamp 1666464484
transform -1 0 3248 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output184
timestamp 1666464484
transform -1 0 3248 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output185
timestamp 1666464484
transform -1 0 3248 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output186
timestamp 1666464484
transform -1 0 5040 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output187
timestamp 1666464484
transform -1 0 3248 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output188
timestamp 1666464484
transform -1 0 3248 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output189
timestamp 1666464484
transform -1 0 3248 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output190
timestamp 1666464484
transform -1 0 3248 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output191
timestamp 1666464484
transform -1 0 3248 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output192
timestamp 1666464484
transform -1 0 3248 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output193
timestamp 1666464484
transform -1 0 5040 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output194
timestamp 1666464484
transform -1 0 5040 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output195
timestamp 1666464484
transform -1 0 3248 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output196
timestamp 1666464484
transform -1 0 3248 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output197
timestamp 1666464484
transform -1 0 3248 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output198
timestamp 1666464484
transform -1 0 3248 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output199
timestamp 1666464484
transform -1 0 3248 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output200
timestamp 1666464484
transform -1 0 3248 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output201
timestamp 1666464484
transform -1 0 3248 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output202
timestamp 1666464484
transform -1 0 5040 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output203
timestamp 1666464484
transform 1 0 74928 0 -1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output204
timestamp 1666464484
transform -1 0 3248 0 -1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output205
timestamp 1666464484
transform -1 0 50288 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output206
timestamp 1666464484
transform 1 0 55104 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output207
timestamp 1666464484
transform 1 0 57344 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output208
timestamp 1666464484
transform 1 0 58352 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output209
timestamp 1666464484
transform -1 0 58688 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output210
timestamp 1666464484
transform 1 0 59136 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output211
timestamp 1666464484
transform 1 0 60480 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output212
timestamp 1666464484
transform -1 0 60704 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output213
timestamp 1666464484
transform 1 0 60928 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output214
timestamp 1666464484
transform 1 0 62272 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output215
timestamp 1666464484
transform 1 0 61264 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output216
timestamp 1666464484
transform 1 0 49392 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output217
timestamp 1666464484
transform -1 0 64288 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output218
timestamp 1666464484
transform 1 0 64400 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output219
timestamp 1666464484
transform -1 0 64736 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output220
timestamp 1666464484
transform 1 0 65296 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output221
timestamp 1666464484
transform 1 0 66192 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output222
timestamp 1666464484
transform -1 0 66752 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output223
timestamp 1666464484
transform 1 0 67088 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output224
timestamp 1666464484
transform 1 0 68320 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output225
timestamp 1666464484
transform 1 0 67200 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output226
timestamp 1666464484
transform 1 0 68880 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output227
timestamp 1666464484
transform 1 0 50512 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output228
timestamp 1666464484
transform -1 0 71680 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output229
timestamp 1666464484
transform 1 0 69216 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output230
timestamp 1666464484
transform 1 0 51184 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output231
timestamp 1666464484
transform 1 0 52640 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output232
timestamp 1666464484
transform 1 0 52976 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output233
timestamp 1666464484
transform 1 0 54432 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output234
timestamp 1666464484
transform 1 0 53312 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output235
timestamp 1666464484
transform -1 0 56336 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output236
timestamp 1666464484
transform 1 0 56560 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output237
timestamp 1666464484
transform 1 0 76720 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output238
timestamp 1666464484
transform 1 0 74928 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output239
timestamp 1666464484
transform 1 0 75152 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output240
timestamp 1666464484
transform 1 0 76720 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output241
timestamp 1666464484
transform 1 0 74928 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output242
timestamp 1666464484
transform 1 0 76720 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output243
timestamp 1666464484
transform 1 0 74928 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output244
timestamp 1666464484
transform 1 0 76720 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output245
timestamp 1666464484
transform 1 0 74928 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output246
timestamp 1666464484
transform 1 0 75152 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output247
timestamp 1666464484
transform 1 0 76720 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output248
timestamp 1666464484
transform 1 0 74928 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output249
timestamp 1666464484
transform 1 0 74928 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output250
timestamp 1666464484
transform 1 0 76720 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output251
timestamp 1666464484
transform 1 0 74928 0 -1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output252
timestamp 1666464484
transform 1 0 76720 0 -1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output253
timestamp 1666464484
transform 1 0 76720 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output254
timestamp 1666464484
transform 1 0 76720 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output255
timestamp 1666464484
transform 1 0 74928 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output256
timestamp 1666464484
transform 1 0 76720 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output257
timestamp 1666464484
transform 1 0 75152 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output258
timestamp 1666464484
transform 1 0 74928 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output259
timestamp 1666464484
transform 1 0 76720 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output260
timestamp 1666464484
transform 1 0 76720 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output261
timestamp 1666464484
transform 1 0 74928 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output262
timestamp 1666464484
transform 1 0 74928 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output263
timestamp 1666464484
transform 1 0 75152 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output264
timestamp 1666464484
transform 1 0 76720 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output265
timestamp 1666464484
transform 1 0 74928 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output266
timestamp 1666464484
transform 1 0 76720 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output267
timestamp 1666464484
transform 1 0 74928 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output268
timestamp 1666464484
transform 1 0 76720 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output269
timestamp 1666464484
transform -1 0 3248 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output270
timestamp 1666464484
transform -1 0 3248 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output271
timestamp 1666464484
transform -1 0 3248 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output272
timestamp 1666464484
transform -1 0 5040 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output273
timestamp 1666464484
transform -1 0 3248 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output274
timestamp 1666464484
transform -1 0 3248 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output275
timestamp 1666464484
transform -1 0 3248 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output276
timestamp 1666464484
transform -1 0 3248 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output277
timestamp 1666464484
transform -1 0 3248 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output278
timestamp 1666464484
transform -1 0 3248 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output279
timestamp 1666464484
transform -1 0 3248 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output280
timestamp 1666464484
transform -1 0 3248 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output281
timestamp 1666464484
transform -1 0 3248 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output282
timestamp 1666464484
transform -1 0 3248 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output283
timestamp 1666464484
transform -1 0 3248 0 -1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output284
timestamp 1666464484
transform -1 0 3248 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output285
timestamp 1666464484
transform -1 0 3248 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output286
timestamp 1666464484
transform -1 0 3248 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output287
timestamp 1666464484
transform -1 0 3248 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output288
timestamp 1666464484
transform -1 0 3248 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output289
timestamp 1666464484
transform -1 0 3248 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output290
timestamp 1666464484
transform -1 0 3248 0 1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output291
timestamp 1666464484
transform -1 0 3248 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output292
timestamp 1666464484
transform -1 0 3248 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output293
timestamp 1666464484
transform -1 0 3248 0 1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output294
timestamp 1666464484
transform -1 0 3248 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output295
timestamp 1666464484
transform -1 0 3248 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output296
timestamp 1666464484
transform -1 0 5040 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output297
timestamp 1666464484
transform -1 0 3248 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output298
timestamp 1666464484
transform -1 0 3248 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output299
timestamp 1666464484
transform -1 0 3248 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output300
timestamp 1666464484
transform -1 0 3248 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output301
timestamp 1666464484
transform 1 0 76720 0 -1 72128
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output302
timestamp 1666464484
transform 1 0 74928 0 -1 72128
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output303
timestamp 1666464484
transform 1 0 76720 0 -1 73696
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output304
timestamp 1666464484
transform 1 0 74928 0 -1 73696
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output305
timestamp 1666464484
transform -1 0 3248 0 1 70560
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output306
timestamp 1666464484
transform -1 0 3248 0 -1 72128
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output307
timestamp 1666464484
transform -1 0 3248 0 1 72128
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output308
timestamp 1666464484
transform -1 0 3248 0 -1 73696
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output309
timestamp 1666464484
transform 1 0 76720 0 -1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output310
timestamp 1666464484
transform -1 0 3248 0 1 73696
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output311
timestamp 1666464484
transform 1 0 76720 0 -1 70560
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output312
timestamp 1666464484
transform -1 0 3248 0 -1 70560
box -86 -86 1654 870
<< labels >>
flabel metal2 s 73808 0 73920 800 0 FreeSans 448 90 0 0 io_wbs_ack
port 0 nsew signal tristate
flabel metal3 s 79200 73808 80000 73920 0 FreeSans 448 0 0 0 io_wbs_ack_0
port 1 nsew signal input
flabel metal3 s 0 73808 800 73920 0 FreeSans 448 0 0 0 io_wbs_ack_1
port 2 nsew signal input
flabel metal2 s 5264 0 5376 800 0 FreeSans 448 90 0 0 io_wbs_adr[0]
port 3 nsew signal input
flabel metal2 s 11984 0 12096 800 0 FreeSans 448 90 0 0 io_wbs_adr[10]
port 4 nsew signal input
flabel metal2 s 12656 0 12768 800 0 FreeSans 448 90 0 0 io_wbs_adr[11]
port 5 nsew signal input
flabel metal2 s 13328 0 13440 800 0 FreeSans 448 90 0 0 io_wbs_adr[12]
port 6 nsew signal input
flabel metal2 s 14000 0 14112 800 0 FreeSans 448 90 0 0 io_wbs_adr[13]
port 7 nsew signal input
flabel metal2 s 14672 0 14784 800 0 FreeSans 448 90 0 0 io_wbs_adr[14]
port 8 nsew signal input
flabel metal2 s 15344 0 15456 800 0 FreeSans 448 90 0 0 io_wbs_adr[15]
port 9 nsew signal input
flabel metal2 s 16016 0 16128 800 0 FreeSans 448 90 0 0 io_wbs_adr[16]
port 10 nsew signal input
flabel metal2 s 16688 0 16800 800 0 FreeSans 448 90 0 0 io_wbs_adr[17]
port 11 nsew signal input
flabel metal2 s 17360 0 17472 800 0 FreeSans 448 90 0 0 io_wbs_adr[18]
port 12 nsew signal input
flabel metal2 s 18032 0 18144 800 0 FreeSans 448 90 0 0 io_wbs_adr[19]
port 13 nsew signal input
flabel metal2 s 5936 0 6048 800 0 FreeSans 448 90 0 0 io_wbs_adr[1]
port 14 nsew signal input
flabel metal2 s 18704 0 18816 800 0 FreeSans 448 90 0 0 io_wbs_adr[20]
port 15 nsew signal input
flabel metal2 s 19376 0 19488 800 0 FreeSans 448 90 0 0 io_wbs_adr[21]
port 16 nsew signal input
flabel metal2 s 20048 0 20160 800 0 FreeSans 448 90 0 0 io_wbs_adr[22]
port 17 nsew signal input
flabel metal2 s 20720 0 20832 800 0 FreeSans 448 90 0 0 io_wbs_adr[23]
port 18 nsew signal input
flabel metal2 s 21392 0 21504 800 0 FreeSans 448 90 0 0 io_wbs_adr[24]
port 19 nsew signal input
flabel metal2 s 22064 0 22176 800 0 FreeSans 448 90 0 0 io_wbs_adr[25]
port 20 nsew signal input
flabel metal2 s 22736 0 22848 800 0 FreeSans 448 90 0 0 io_wbs_adr[26]
port 21 nsew signal input
flabel metal2 s 23408 0 23520 800 0 FreeSans 448 90 0 0 io_wbs_adr[27]
port 22 nsew signal input
flabel metal2 s 24080 0 24192 800 0 FreeSans 448 90 0 0 io_wbs_adr[28]
port 23 nsew signal input
flabel metal2 s 24752 0 24864 800 0 FreeSans 448 90 0 0 io_wbs_adr[29]
port 24 nsew signal input
flabel metal2 s 6608 0 6720 800 0 FreeSans 448 90 0 0 io_wbs_adr[2]
port 25 nsew signal input
flabel metal2 s 25424 0 25536 800 0 FreeSans 448 90 0 0 io_wbs_adr[30]
port 26 nsew signal input
flabel metal2 s 26096 0 26208 800 0 FreeSans 448 90 0 0 io_wbs_adr[31]
port 27 nsew signal input
flabel metal2 s 7280 0 7392 800 0 FreeSans 448 90 0 0 io_wbs_adr[3]
port 28 nsew signal input
flabel metal2 s 7952 0 8064 800 0 FreeSans 448 90 0 0 io_wbs_adr[4]
port 29 nsew signal input
flabel metal2 s 8624 0 8736 800 0 FreeSans 448 90 0 0 io_wbs_adr[5]
port 30 nsew signal input
flabel metal2 s 9296 0 9408 800 0 FreeSans 448 90 0 0 io_wbs_adr[6]
port 31 nsew signal input
flabel metal2 s 9968 0 10080 800 0 FreeSans 448 90 0 0 io_wbs_adr[7]
port 32 nsew signal input
flabel metal2 s 10640 0 10752 800 0 FreeSans 448 90 0 0 io_wbs_adr[8]
port 33 nsew signal input
flabel metal2 s 11312 0 11424 800 0 FreeSans 448 90 0 0 io_wbs_adr[9]
port 34 nsew signal input
flabel metal3 s 79200 5264 80000 5376 0 FreeSans 448 0 0 0 io_wbs_adr_0[0]
port 35 nsew signal tristate
flabel metal3 s 79200 11984 80000 12096 0 FreeSans 448 0 0 0 io_wbs_adr_0[10]
port 36 nsew signal tristate
flabel metal3 s 79200 12656 80000 12768 0 FreeSans 448 0 0 0 io_wbs_adr_0[11]
port 37 nsew signal tristate
flabel metal3 s 79200 13328 80000 13440 0 FreeSans 448 0 0 0 io_wbs_adr_0[12]
port 38 nsew signal tristate
flabel metal3 s 79200 14000 80000 14112 0 FreeSans 448 0 0 0 io_wbs_adr_0[13]
port 39 nsew signal tristate
flabel metal3 s 79200 14672 80000 14784 0 FreeSans 448 0 0 0 io_wbs_adr_0[14]
port 40 nsew signal tristate
flabel metal3 s 79200 15344 80000 15456 0 FreeSans 448 0 0 0 io_wbs_adr_0[15]
port 41 nsew signal tristate
flabel metal3 s 79200 16016 80000 16128 0 FreeSans 448 0 0 0 io_wbs_adr_0[16]
port 42 nsew signal tristate
flabel metal3 s 79200 16688 80000 16800 0 FreeSans 448 0 0 0 io_wbs_adr_0[17]
port 43 nsew signal tristate
flabel metal3 s 79200 17360 80000 17472 0 FreeSans 448 0 0 0 io_wbs_adr_0[18]
port 44 nsew signal tristate
flabel metal3 s 79200 18032 80000 18144 0 FreeSans 448 0 0 0 io_wbs_adr_0[19]
port 45 nsew signal tristate
flabel metal3 s 79200 5936 80000 6048 0 FreeSans 448 0 0 0 io_wbs_adr_0[1]
port 46 nsew signal tristate
flabel metal3 s 79200 18704 80000 18816 0 FreeSans 448 0 0 0 io_wbs_adr_0[20]
port 47 nsew signal tristate
flabel metal3 s 79200 19376 80000 19488 0 FreeSans 448 0 0 0 io_wbs_adr_0[21]
port 48 nsew signal tristate
flabel metal3 s 79200 20048 80000 20160 0 FreeSans 448 0 0 0 io_wbs_adr_0[22]
port 49 nsew signal tristate
flabel metal3 s 79200 20720 80000 20832 0 FreeSans 448 0 0 0 io_wbs_adr_0[23]
port 50 nsew signal tristate
flabel metal3 s 79200 21392 80000 21504 0 FreeSans 448 0 0 0 io_wbs_adr_0[24]
port 51 nsew signal tristate
flabel metal3 s 79200 22064 80000 22176 0 FreeSans 448 0 0 0 io_wbs_adr_0[25]
port 52 nsew signal tristate
flabel metal3 s 79200 22736 80000 22848 0 FreeSans 448 0 0 0 io_wbs_adr_0[26]
port 53 nsew signal tristate
flabel metal3 s 79200 23408 80000 23520 0 FreeSans 448 0 0 0 io_wbs_adr_0[27]
port 54 nsew signal tristate
flabel metal3 s 79200 24080 80000 24192 0 FreeSans 448 0 0 0 io_wbs_adr_0[28]
port 55 nsew signal tristate
flabel metal3 s 79200 24752 80000 24864 0 FreeSans 448 0 0 0 io_wbs_adr_0[29]
port 56 nsew signal tristate
flabel metal3 s 79200 6608 80000 6720 0 FreeSans 448 0 0 0 io_wbs_adr_0[2]
port 57 nsew signal tristate
flabel metal3 s 79200 25424 80000 25536 0 FreeSans 448 0 0 0 io_wbs_adr_0[30]
port 58 nsew signal tristate
flabel metal3 s 79200 26096 80000 26208 0 FreeSans 448 0 0 0 io_wbs_adr_0[31]
port 59 nsew signal tristate
flabel metal3 s 79200 7280 80000 7392 0 FreeSans 448 0 0 0 io_wbs_adr_0[3]
port 60 nsew signal tristate
flabel metal3 s 79200 7952 80000 8064 0 FreeSans 448 0 0 0 io_wbs_adr_0[4]
port 61 nsew signal tristate
flabel metal3 s 79200 8624 80000 8736 0 FreeSans 448 0 0 0 io_wbs_adr_0[5]
port 62 nsew signal tristate
flabel metal3 s 79200 9296 80000 9408 0 FreeSans 448 0 0 0 io_wbs_adr_0[6]
port 63 nsew signal tristate
flabel metal3 s 79200 9968 80000 10080 0 FreeSans 448 0 0 0 io_wbs_adr_0[7]
port 64 nsew signal tristate
flabel metal3 s 79200 10640 80000 10752 0 FreeSans 448 0 0 0 io_wbs_adr_0[8]
port 65 nsew signal tristate
flabel metal3 s 79200 11312 80000 11424 0 FreeSans 448 0 0 0 io_wbs_adr_0[9]
port 66 nsew signal tristate
flabel metal3 s 0 5264 800 5376 0 FreeSans 448 0 0 0 io_wbs_adr_1[0]
port 67 nsew signal tristate
flabel metal3 s 0 11984 800 12096 0 FreeSans 448 0 0 0 io_wbs_adr_1[10]
port 68 nsew signal tristate
flabel metal3 s 0 12656 800 12768 0 FreeSans 448 0 0 0 io_wbs_adr_1[11]
port 69 nsew signal tristate
flabel metal3 s 0 13328 800 13440 0 FreeSans 448 0 0 0 io_wbs_adr_1[12]
port 70 nsew signal tristate
flabel metal3 s 0 14000 800 14112 0 FreeSans 448 0 0 0 io_wbs_adr_1[13]
port 71 nsew signal tristate
flabel metal3 s 0 14672 800 14784 0 FreeSans 448 0 0 0 io_wbs_adr_1[14]
port 72 nsew signal tristate
flabel metal3 s 0 15344 800 15456 0 FreeSans 448 0 0 0 io_wbs_adr_1[15]
port 73 nsew signal tristate
flabel metal3 s 0 16016 800 16128 0 FreeSans 448 0 0 0 io_wbs_adr_1[16]
port 74 nsew signal tristate
flabel metal3 s 0 16688 800 16800 0 FreeSans 448 0 0 0 io_wbs_adr_1[17]
port 75 nsew signal tristate
flabel metal3 s 0 17360 800 17472 0 FreeSans 448 0 0 0 io_wbs_adr_1[18]
port 76 nsew signal tristate
flabel metal3 s 0 18032 800 18144 0 FreeSans 448 0 0 0 io_wbs_adr_1[19]
port 77 nsew signal tristate
flabel metal3 s 0 5936 800 6048 0 FreeSans 448 0 0 0 io_wbs_adr_1[1]
port 78 nsew signal tristate
flabel metal3 s 0 18704 800 18816 0 FreeSans 448 0 0 0 io_wbs_adr_1[20]
port 79 nsew signal tristate
flabel metal3 s 0 19376 800 19488 0 FreeSans 448 0 0 0 io_wbs_adr_1[21]
port 80 nsew signal tristate
flabel metal3 s 0 20048 800 20160 0 FreeSans 448 0 0 0 io_wbs_adr_1[22]
port 81 nsew signal tristate
flabel metal3 s 0 20720 800 20832 0 FreeSans 448 0 0 0 io_wbs_adr_1[23]
port 82 nsew signal tristate
flabel metal3 s 0 21392 800 21504 0 FreeSans 448 0 0 0 io_wbs_adr_1[24]
port 83 nsew signal tristate
flabel metal3 s 0 22064 800 22176 0 FreeSans 448 0 0 0 io_wbs_adr_1[25]
port 84 nsew signal tristate
flabel metal3 s 0 22736 800 22848 0 FreeSans 448 0 0 0 io_wbs_adr_1[26]
port 85 nsew signal tristate
flabel metal3 s 0 23408 800 23520 0 FreeSans 448 0 0 0 io_wbs_adr_1[27]
port 86 nsew signal tristate
flabel metal3 s 0 24080 800 24192 0 FreeSans 448 0 0 0 io_wbs_adr_1[28]
port 87 nsew signal tristate
flabel metal3 s 0 24752 800 24864 0 FreeSans 448 0 0 0 io_wbs_adr_1[29]
port 88 nsew signal tristate
flabel metal3 s 0 6608 800 6720 0 FreeSans 448 0 0 0 io_wbs_adr_1[2]
port 89 nsew signal tristate
flabel metal3 s 0 25424 800 25536 0 FreeSans 448 0 0 0 io_wbs_adr_1[30]
port 90 nsew signal tristate
flabel metal3 s 0 26096 800 26208 0 FreeSans 448 0 0 0 io_wbs_adr_1[31]
port 91 nsew signal tristate
flabel metal3 s 0 7280 800 7392 0 FreeSans 448 0 0 0 io_wbs_adr_1[3]
port 92 nsew signal tristate
flabel metal3 s 0 7952 800 8064 0 FreeSans 448 0 0 0 io_wbs_adr_1[4]
port 93 nsew signal tristate
flabel metal3 s 0 8624 800 8736 0 FreeSans 448 0 0 0 io_wbs_adr_1[5]
port 94 nsew signal tristate
flabel metal3 s 0 9296 800 9408 0 FreeSans 448 0 0 0 io_wbs_adr_1[6]
port 95 nsew signal tristate
flabel metal3 s 0 9968 800 10080 0 FreeSans 448 0 0 0 io_wbs_adr_1[7]
port 96 nsew signal tristate
flabel metal3 s 0 10640 800 10752 0 FreeSans 448 0 0 0 io_wbs_adr_1[8]
port 97 nsew signal tristate
flabel metal3 s 0 11312 800 11424 0 FreeSans 448 0 0 0 io_wbs_adr_1[9]
port 98 nsew signal tristate
flabel metal2 s 74480 0 74592 800 0 FreeSans 448 90 0 0 io_wbs_cyc
port 99 nsew signal input
flabel metal3 s 79200 74480 80000 74592 0 FreeSans 448 0 0 0 io_wbs_cyc_0
port 100 nsew signal tristate
flabel metal3 s 0 74480 800 74592 0 FreeSans 448 0 0 0 io_wbs_cyc_1
port 101 nsew signal tristate
flabel metal2 s 48272 0 48384 800 0 FreeSans 448 90 0 0 io_wbs_datrd[0]
port 102 nsew signal tristate
flabel metal2 s 54992 0 55104 800 0 FreeSans 448 90 0 0 io_wbs_datrd[10]
port 103 nsew signal tristate
flabel metal2 s 55664 0 55776 800 0 FreeSans 448 90 0 0 io_wbs_datrd[11]
port 104 nsew signal tristate
flabel metal2 s 56336 0 56448 800 0 FreeSans 448 90 0 0 io_wbs_datrd[12]
port 105 nsew signal tristate
flabel metal2 s 57008 0 57120 800 0 FreeSans 448 90 0 0 io_wbs_datrd[13]
port 106 nsew signal tristate
flabel metal2 s 57680 0 57792 800 0 FreeSans 448 90 0 0 io_wbs_datrd[14]
port 107 nsew signal tristate
flabel metal2 s 58352 0 58464 800 0 FreeSans 448 90 0 0 io_wbs_datrd[15]
port 108 nsew signal tristate
flabel metal2 s 59024 0 59136 800 0 FreeSans 448 90 0 0 io_wbs_datrd[16]
port 109 nsew signal tristate
flabel metal2 s 59696 0 59808 800 0 FreeSans 448 90 0 0 io_wbs_datrd[17]
port 110 nsew signal tristate
flabel metal2 s 60368 0 60480 800 0 FreeSans 448 90 0 0 io_wbs_datrd[18]
port 111 nsew signal tristate
flabel metal2 s 61040 0 61152 800 0 FreeSans 448 90 0 0 io_wbs_datrd[19]
port 112 nsew signal tristate
flabel metal2 s 48944 0 49056 800 0 FreeSans 448 90 0 0 io_wbs_datrd[1]
port 113 nsew signal tristate
flabel metal2 s 61712 0 61824 800 0 FreeSans 448 90 0 0 io_wbs_datrd[20]
port 114 nsew signal tristate
flabel metal2 s 62384 0 62496 800 0 FreeSans 448 90 0 0 io_wbs_datrd[21]
port 115 nsew signal tristate
flabel metal2 s 63056 0 63168 800 0 FreeSans 448 90 0 0 io_wbs_datrd[22]
port 116 nsew signal tristate
flabel metal2 s 63728 0 63840 800 0 FreeSans 448 90 0 0 io_wbs_datrd[23]
port 117 nsew signal tristate
flabel metal2 s 64400 0 64512 800 0 FreeSans 448 90 0 0 io_wbs_datrd[24]
port 118 nsew signal tristate
flabel metal2 s 65072 0 65184 800 0 FreeSans 448 90 0 0 io_wbs_datrd[25]
port 119 nsew signal tristate
flabel metal2 s 65744 0 65856 800 0 FreeSans 448 90 0 0 io_wbs_datrd[26]
port 120 nsew signal tristate
flabel metal2 s 66416 0 66528 800 0 FreeSans 448 90 0 0 io_wbs_datrd[27]
port 121 nsew signal tristate
flabel metal2 s 67088 0 67200 800 0 FreeSans 448 90 0 0 io_wbs_datrd[28]
port 122 nsew signal tristate
flabel metal2 s 67760 0 67872 800 0 FreeSans 448 90 0 0 io_wbs_datrd[29]
port 123 nsew signal tristate
flabel metal2 s 49616 0 49728 800 0 FreeSans 448 90 0 0 io_wbs_datrd[2]
port 124 nsew signal tristate
flabel metal2 s 68432 0 68544 800 0 FreeSans 448 90 0 0 io_wbs_datrd[30]
port 125 nsew signal tristate
flabel metal2 s 69104 0 69216 800 0 FreeSans 448 90 0 0 io_wbs_datrd[31]
port 126 nsew signal tristate
flabel metal2 s 50288 0 50400 800 0 FreeSans 448 90 0 0 io_wbs_datrd[3]
port 127 nsew signal tristate
flabel metal2 s 50960 0 51072 800 0 FreeSans 448 90 0 0 io_wbs_datrd[4]
port 128 nsew signal tristate
flabel metal2 s 51632 0 51744 800 0 FreeSans 448 90 0 0 io_wbs_datrd[5]
port 129 nsew signal tristate
flabel metal2 s 52304 0 52416 800 0 FreeSans 448 90 0 0 io_wbs_datrd[6]
port 130 nsew signal tristate
flabel metal2 s 52976 0 53088 800 0 FreeSans 448 90 0 0 io_wbs_datrd[7]
port 131 nsew signal tristate
flabel metal2 s 53648 0 53760 800 0 FreeSans 448 90 0 0 io_wbs_datrd[8]
port 132 nsew signal tristate
flabel metal2 s 54320 0 54432 800 0 FreeSans 448 90 0 0 io_wbs_datrd[9]
port 133 nsew signal tristate
flabel metal3 s 79200 48272 80000 48384 0 FreeSans 448 0 0 0 io_wbs_datrd_0[0]
port 134 nsew signal input
flabel metal3 s 79200 54992 80000 55104 0 FreeSans 448 0 0 0 io_wbs_datrd_0[10]
port 135 nsew signal input
flabel metal3 s 79200 55664 80000 55776 0 FreeSans 448 0 0 0 io_wbs_datrd_0[11]
port 136 nsew signal input
flabel metal3 s 79200 56336 80000 56448 0 FreeSans 448 0 0 0 io_wbs_datrd_0[12]
port 137 nsew signal input
flabel metal3 s 79200 57008 80000 57120 0 FreeSans 448 0 0 0 io_wbs_datrd_0[13]
port 138 nsew signal input
flabel metal3 s 79200 57680 80000 57792 0 FreeSans 448 0 0 0 io_wbs_datrd_0[14]
port 139 nsew signal input
flabel metal3 s 79200 58352 80000 58464 0 FreeSans 448 0 0 0 io_wbs_datrd_0[15]
port 140 nsew signal input
flabel metal3 s 79200 59024 80000 59136 0 FreeSans 448 0 0 0 io_wbs_datrd_0[16]
port 141 nsew signal input
flabel metal3 s 79200 59696 80000 59808 0 FreeSans 448 0 0 0 io_wbs_datrd_0[17]
port 142 nsew signal input
flabel metal3 s 79200 60368 80000 60480 0 FreeSans 448 0 0 0 io_wbs_datrd_0[18]
port 143 nsew signal input
flabel metal3 s 79200 61040 80000 61152 0 FreeSans 448 0 0 0 io_wbs_datrd_0[19]
port 144 nsew signal input
flabel metal3 s 79200 48944 80000 49056 0 FreeSans 448 0 0 0 io_wbs_datrd_0[1]
port 145 nsew signal input
flabel metal3 s 79200 61712 80000 61824 0 FreeSans 448 0 0 0 io_wbs_datrd_0[20]
port 146 nsew signal input
flabel metal3 s 79200 62384 80000 62496 0 FreeSans 448 0 0 0 io_wbs_datrd_0[21]
port 147 nsew signal input
flabel metal3 s 79200 63056 80000 63168 0 FreeSans 448 0 0 0 io_wbs_datrd_0[22]
port 148 nsew signal input
flabel metal3 s 79200 63728 80000 63840 0 FreeSans 448 0 0 0 io_wbs_datrd_0[23]
port 149 nsew signal input
flabel metal3 s 79200 64400 80000 64512 0 FreeSans 448 0 0 0 io_wbs_datrd_0[24]
port 150 nsew signal input
flabel metal3 s 79200 65072 80000 65184 0 FreeSans 448 0 0 0 io_wbs_datrd_0[25]
port 151 nsew signal input
flabel metal3 s 79200 65744 80000 65856 0 FreeSans 448 0 0 0 io_wbs_datrd_0[26]
port 152 nsew signal input
flabel metal3 s 79200 66416 80000 66528 0 FreeSans 448 0 0 0 io_wbs_datrd_0[27]
port 153 nsew signal input
flabel metal3 s 79200 67088 80000 67200 0 FreeSans 448 0 0 0 io_wbs_datrd_0[28]
port 154 nsew signal input
flabel metal3 s 79200 67760 80000 67872 0 FreeSans 448 0 0 0 io_wbs_datrd_0[29]
port 155 nsew signal input
flabel metal3 s 79200 49616 80000 49728 0 FreeSans 448 0 0 0 io_wbs_datrd_0[2]
port 156 nsew signal input
flabel metal3 s 79200 68432 80000 68544 0 FreeSans 448 0 0 0 io_wbs_datrd_0[30]
port 157 nsew signal input
flabel metal3 s 79200 69104 80000 69216 0 FreeSans 448 0 0 0 io_wbs_datrd_0[31]
port 158 nsew signal input
flabel metal3 s 79200 50288 80000 50400 0 FreeSans 448 0 0 0 io_wbs_datrd_0[3]
port 159 nsew signal input
flabel metal3 s 79200 50960 80000 51072 0 FreeSans 448 0 0 0 io_wbs_datrd_0[4]
port 160 nsew signal input
flabel metal3 s 79200 51632 80000 51744 0 FreeSans 448 0 0 0 io_wbs_datrd_0[5]
port 161 nsew signal input
flabel metal3 s 79200 52304 80000 52416 0 FreeSans 448 0 0 0 io_wbs_datrd_0[6]
port 162 nsew signal input
flabel metal3 s 79200 52976 80000 53088 0 FreeSans 448 0 0 0 io_wbs_datrd_0[7]
port 163 nsew signal input
flabel metal3 s 79200 53648 80000 53760 0 FreeSans 448 0 0 0 io_wbs_datrd_0[8]
port 164 nsew signal input
flabel metal3 s 79200 54320 80000 54432 0 FreeSans 448 0 0 0 io_wbs_datrd_0[9]
port 165 nsew signal input
flabel metal3 s 0 48272 800 48384 0 FreeSans 448 0 0 0 io_wbs_datrd_1[0]
port 166 nsew signal input
flabel metal3 s 0 54992 800 55104 0 FreeSans 448 0 0 0 io_wbs_datrd_1[10]
port 167 nsew signal input
flabel metal3 s 0 55664 800 55776 0 FreeSans 448 0 0 0 io_wbs_datrd_1[11]
port 168 nsew signal input
flabel metal3 s 0 56336 800 56448 0 FreeSans 448 0 0 0 io_wbs_datrd_1[12]
port 169 nsew signal input
flabel metal3 s 0 57008 800 57120 0 FreeSans 448 0 0 0 io_wbs_datrd_1[13]
port 170 nsew signal input
flabel metal3 s 0 57680 800 57792 0 FreeSans 448 0 0 0 io_wbs_datrd_1[14]
port 171 nsew signal input
flabel metal3 s 0 58352 800 58464 0 FreeSans 448 0 0 0 io_wbs_datrd_1[15]
port 172 nsew signal input
flabel metal3 s 0 59024 800 59136 0 FreeSans 448 0 0 0 io_wbs_datrd_1[16]
port 173 nsew signal input
flabel metal3 s 0 59696 800 59808 0 FreeSans 448 0 0 0 io_wbs_datrd_1[17]
port 174 nsew signal input
flabel metal3 s 0 60368 800 60480 0 FreeSans 448 0 0 0 io_wbs_datrd_1[18]
port 175 nsew signal input
flabel metal3 s 0 61040 800 61152 0 FreeSans 448 0 0 0 io_wbs_datrd_1[19]
port 176 nsew signal input
flabel metal3 s 0 48944 800 49056 0 FreeSans 448 0 0 0 io_wbs_datrd_1[1]
port 177 nsew signal input
flabel metal3 s 0 61712 800 61824 0 FreeSans 448 0 0 0 io_wbs_datrd_1[20]
port 178 nsew signal input
flabel metal3 s 0 62384 800 62496 0 FreeSans 448 0 0 0 io_wbs_datrd_1[21]
port 179 nsew signal input
flabel metal3 s 0 63056 800 63168 0 FreeSans 448 0 0 0 io_wbs_datrd_1[22]
port 180 nsew signal input
flabel metal3 s 0 63728 800 63840 0 FreeSans 448 0 0 0 io_wbs_datrd_1[23]
port 181 nsew signal input
flabel metal3 s 0 64400 800 64512 0 FreeSans 448 0 0 0 io_wbs_datrd_1[24]
port 182 nsew signal input
flabel metal3 s 0 65072 800 65184 0 FreeSans 448 0 0 0 io_wbs_datrd_1[25]
port 183 nsew signal input
flabel metal3 s 0 65744 800 65856 0 FreeSans 448 0 0 0 io_wbs_datrd_1[26]
port 184 nsew signal input
flabel metal3 s 0 66416 800 66528 0 FreeSans 448 0 0 0 io_wbs_datrd_1[27]
port 185 nsew signal input
flabel metal3 s 0 67088 800 67200 0 FreeSans 448 0 0 0 io_wbs_datrd_1[28]
port 186 nsew signal input
flabel metal3 s 0 67760 800 67872 0 FreeSans 448 0 0 0 io_wbs_datrd_1[29]
port 187 nsew signal input
flabel metal3 s 0 49616 800 49728 0 FreeSans 448 0 0 0 io_wbs_datrd_1[2]
port 188 nsew signal input
flabel metal3 s 0 68432 800 68544 0 FreeSans 448 0 0 0 io_wbs_datrd_1[30]
port 189 nsew signal input
flabel metal3 s 0 69104 800 69216 0 FreeSans 448 0 0 0 io_wbs_datrd_1[31]
port 190 nsew signal input
flabel metal3 s 0 50288 800 50400 0 FreeSans 448 0 0 0 io_wbs_datrd_1[3]
port 191 nsew signal input
flabel metal3 s 0 50960 800 51072 0 FreeSans 448 0 0 0 io_wbs_datrd_1[4]
port 192 nsew signal input
flabel metal3 s 0 51632 800 51744 0 FreeSans 448 0 0 0 io_wbs_datrd_1[5]
port 193 nsew signal input
flabel metal3 s 0 52304 800 52416 0 FreeSans 448 0 0 0 io_wbs_datrd_1[6]
port 194 nsew signal input
flabel metal3 s 0 52976 800 53088 0 FreeSans 448 0 0 0 io_wbs_datrd_1[7]
port 195 nsew signal input
flabel metal3 s 0 53648 800 53760 0 FreeSans 448 0 0 0 io_wbs_datrd_1[8]
port 196 nsew signal input
flabel metal3 s 0 54320 800 54432 0 FreeSans 448 0 0 0 io_wbs_datrd_1[9]
port 197 nsew signal input
flabel metal2 s 26768 0 26880 800 0 FreeSans 448 90 0 0 io_wbs_datwr[0]
port 198 nsew signal input
flabel metal2 s 33488 0 33600 800 0 FreeSans 448 90 0 0 io_wbs_datwr[10]
port 199 nsew signal input
flabel metal2 s 34160 0 34272 800 0 FreeSans 448 90 0 0 io_wbs_datwr[11]
port 200 nsew signal input
flabel metal2 s 34832 0 34944 800 0 FreeSans 448 90 0 0 io_wbs_datwr[12]
port 201 nsew signal input
flabel metal2 s 35504 0 35616 800 0 FreeSans 448 90 0 0 io_wbs_datwr[13]
port 202 nsew signal input
flabel metal2 s 36176 0 36288 800 0 FreeSans 448 90 0 0 io_wbs_datwr[14]
port 203 nsew signal input
flabel metal2 s 36848 0 36960 800 0 FreeSans 448 90 0 0 io_wbs_datwr[15]
port 204 nsew signal input
flabel metal2 s 37520 0 37632 800 0 FreeSans 448 90 0 0 io_wbs_datwr[16]
port 205 nsew signal input
flabel metal2 s 38192 0 38304 800 0 FreeSans 448 90 0 0 io_wbs_datwr[17]
port 206 nsew signal input
flabel metal2 s 38864 0 38976 800 0 FreeSans 448 90 0 0 io_wbs_datwr[18]
port 207 nsew signal input
flabel metal2 s 39536 0 39648 800 0 FreeSans 448 90 0 0 io_wbs_datwr[19]
port 208 nsew signal input
flabel metal2 s 27440 0 27552 800 0 FreeSans 448 90 0 0 io_wbs_datwr[1]
port 209 nsew signal input
flabel metal2 s 40208 0 40320 800 0 FreeSans 448 90 0 0 io_wbs_datwr[20]
port 210 nsew signal input
flabel metal2 s 40880 0 40992 800 0 FreeSans 448 90 0 0 io_wbs_datwr[21]
port 211 nsew signal input
flabel metal2 s 41552 0 41664 800 0 FreeSans 448 90 0 0 io_wbs_datwr[22]
port 212 nsew signal input
flabel metal2 s 42224 0 42336 800 0 FreeSans 448 90 0 0 io_wbs_datwr[23]
port 213 nsew signal input
flabel metal2 s 42896 0 43008 800 0 FreeSans 448 90 0 0 io_wbs_datwr[24]
port 214 nsew signal input
flabel metal2 s 43568 0 43680 800 0 FreeSans 448 90 0 0 io_wbs_datwr[25]
port 215 nsew signal input
flabel metal2 s 44240 0 44352 800 0 FreeSans 448 90 0 0 io_wbs_datwr[26]
port 216 nsew signal input
flabel metal2 s 44912 0 45024 800 0 FreeSans 448 90 0 0 io_wbs_datwr[27]
port 217 nsew signal input
flabel metal2 s 45584 0 45696 800 0 FreeSans 448 90 0 0 io_wbs_datwr[28]
port 218 nsew signal input
flabel metal2 s 46256 0 46368 800 0 FreeSans 448 90 0 0 io_wbs_datwr[29]
port 219 nsew signal input
flabel metal2 s 28112 0 28224 800 0 FreeSans 448 90 0 0 io_wbs_datwr[2]
port 220 nsew signal input
flabel metal2 s 46928 0 47040 800 0 FreeSans 448 90 0 0 io_wbs_datwr[30]
port 221 nsew signal input
flabel metal2 s 47600 0 47712 800 0 FreeSans 448 90 0 0 io_wbs_datwr[31]
port 222 nsew signal input
flabel metal2 s 28784 0 28896 800 0 FreeSans 448 90 0 0 io_wbs_datwr[3]
port 223 nsew signal input
flabel metal2 s 29456 0 29568 800 0 FreeSans 448 90 0 0 io_wbs_datwr[4]
port 224 nsew signal input
flabel metal2 s 30128 0 30240 800 0 FreeSans 448 90 0 0 io_wbs_datwr[5]
port 225 nsew signal input
flabel metal2 s 30800 0 30912 800 0 FreeSans 448 90 0 0 io_wbs_datwr[6]
port 226 nsew signal input
flabel metal2 s 31472 0 31584 800 0 FreeSans 448 90 0 0 io_wbs_datwr[7]
port 227 nsew signal input
flabel metal2 s 32144 0 32256 800 0 FreeSans 448 90 0 0 io_wbs_datwr[8]
port 228 nsew signal input
flabel metal2 s 32816 0 32928 800 0 FreeSans 448 90 0 0 io_wbs_datwr[9]
port 229 nsew signal input
flabel metal3 s 79200 26768 80000 26880 0 FreeSans 448 0 0 0 io_wbs_datwr_0[0]
port 230 nsew signal tristate
flabel metal3 s 79200 33488 80000 33600 0 FreeSans 448 0 0 0 io_wbs_datwr_0[10]
port 231 nsew signal tristate
flabel metal3 s 79200 34160 80000 34272 0 FreeSans 448 0 0 0 io_wbs_datwr_0[11]
port 232 nsew signal tristate
flabel metal3 s 79200 34832 80000 34944 0 FreeSans 448 0 0 0 io_wbs_datwr_0[12]
port 233 nsew signal tristate
flabel metal3 s 79200 35504 80000 35616 0 FreeSans 448 0 0 0 io_wbs_datwr_0[13]
port 234 nsew signal tristate
flabel metal3 s 79200 36176 80000 36288 0 FreeSans 448 0 0 0 io_wbs_datwr_0[14]
port 235 nsew signal tristate
flabel metal3 s 79200 36848 80000 36960 0 FreeSans 448 0 0 0 io_wbs_datwr_0[15]
port 236 nsew signal tristate
flabel metal3 s 79200 37520 80000 37632 0 FreeSans 448 0 0 0 io_wbs_datwr_0[16]
port 237 nsew signal tristate
flabel metal3 s 79200 38192 80000 38304 0 FreeSans 448 0 0 0 io_wbs_datwr_0[17]
port 238 nsew signal tristate
flabel metal3 s 79200 38864 80000 38976 0 FreeSans 448 0 0 0 io_wbs_datwr_0[18]
port 239 nsew signal tristate
flabel metal3 s 79200 39536 80000 39648 0 FreeSans 448 0 0 0 io_wbs_datwr_0[19]
port 240 nsew signal tristate
flabel metal3 s 79200 27440 80000 27552 0 FreeSans 448 0 0 0 io_wbs_datwr_0[1]
port 241 nsew signal tristate
flabel metal3 s 79200 40208 80000 40320 0 FreeSans 448 0 0 0 io_wbs_datwr_0[20]
port 242 nsew signal tristate
flabel metal3 s 79200 40880 80000 40992 0 FreeSans 448 0 0 0 io_wbs_datwr_0[21]
port 243 nsew signal tristate
flabel metal3 s 79200 41552 80000 41664 0 FreeSans 448 0 0 0 io_wbs_datwr_0[22]
port 244 nsew signal tristate
flabel metal3 s 79200 42224 80000 42336 0 FreeSans 448 0 0 0 io_wbs_datwr_0[23]
port 245 nsew signal tristate
flabel metal3 s 79200 42896 80000 43008 0 FreeSans 448 0 0 0 io_wbs_datwr_0[24]
port 246 nsew signal tristate
flabel metal3 s 79200 43568 80000 43680 0 FreeSans 448 0 0 0 io_wbs_datwr_0[25]
port 247 nsew signal tristate
flabel metal3 s 79200 44240 80000 44352 0 FreeSans 448 0 0 0 io_wbs_datwr_0[26]
port 248 nsew signal tristate
flabel metal3 s 79200 44912 80000 45024 0 FreeSans 448 0 0 0 io_wbs_datwr_0[27]
port 249 nsew signal tristate
flabel metal3 s 79200 45584 80000 45696 0 FreeSans 448 0 0 0 io_wbs_datwr_0[28]
port 250 nsew signal tristate
flabel metal3 s 79200 46256 80000 46368 0 FreeSans 448 0 0 0 io_wbs_datwr_0[29]
port 251 nsew signal tristate
flabel metal3 s 79200 28112 80000 28224 0 FreeSans 448 0 0 0 io_wbs_datwr_0[2]
port 252 nsew signal tristate
flabel metal3 s 79200 46928 80000 47040 0 FreeSans 448 0 0 0 io_wbs_datwr_0[30]
port 253 nsew signal tristate
flabel metal3 s 79200 47600 80000 47712 0 FreeSans 448 0 0 0 io_wbs_datwr_0[31]
port 254 nsew signal tristate
flabel metal3 s 79200 28784 80000 28896 0 FreeSans 448 0 0 0 io_wbs_datwr_0[3]
port 255 nsew signal tristate
flabel metal3 s 79200 29456 80000 29568 0 FreeSans 448 0 0 0 io_wbs_datwr_0[4]
port 256 nsew signal tristate
flabel metal3 s 79200 30128 80000 30240 0 FreeSans 448 0 0 0 io_wbs_datwr_0[5]
port 257 nsew signal tristate
flabel metal3 s 79200 30800 80000 30912 0 FreeSans 448 0 0 0 io_wbs_datwr_0[6]
port 258 nsew signal tristate
flabel metal3 s 79200 31472 80000 31584 0 FreeSans 448 0 0 0 io_wbs_datwr_0[7]
port 259 nsew signal tristate
flabel metal3 s 79200 32144 80000 32256 0 FreeSans 448 0 0 0 io_wbs_datwr_0[8]
port 260 nsew signal tristate
flabel metal3 s 79200 32816 80000 32928 0 FreeSans 448 0 0 0 io_wbs_datwr_0[9]
port 261 nsew signal tristate
flabel metal3 s 0 26768 800 26880 0 FreeSans 448 0 0 0 io_wbs_datwr_1[0]
port 262 nsew signal tristate
flabel metal3 s 0 33488 800 33600 0 FreeSans 448 0 0 0 io_wbs_datwr_1[10]
port 263 nsew signal tristate
flabel metal3 s 0 34160 800 34272 0 FreeSans 448 0 0 0 io_wbs_datwr_1[11]
port 264 nsew signal tristate
flabel metal3 s 0 34832 800 34944 0 FreeSans 448 0 0 0 io_wbs_datwr_1[12]
port 265 nsew signal tristate
flabel metal3 s 0 35504 800 35616 0 FreeSans 448 0 0 0 io_wbs_datwr_1[13]
port 266 nsew signal tristate
flabel metal3 s 0 36176 800 36288 0 FreeSans 448 0 0 0 io_wbs_datwr_1[14]
port 267 nsew signal tristate
flabel metal3 s 0 36848 800 36960 0 FreeSans 448 0 0 0 io_wbs_datwr_1[15]
port 268 nsew signal tristate
flabel metal3 s 0 37520 800 37632 0 FreeSans 448 0 0 0 io_wbs_datwr_1[16]
port 269 nsew signal tristate
flabel metal3 s 0 38192 800 38304 0 FreeSans 448 0 0 0 io_wbs_datwr_1[17]
port 270 nsew signal tristate
flabel metal3 s 0 38864 800 38976 0 FreeSans 448 0 0 0 io_wbs_datwr_1[18]
port 271 nsew signal tristate
flabel metal3 s 0 39536 800 39648 0 FreeSans 448 0 0 0 io_wbs_datwr_1[19]
port 272 nsew signal tristate
flabel metal3 s 0 27440 800 27552 0 FreeSans 448 0 0 0 io_wbs_datwr_1[1]
port 273 nsew signal tristate
flabel metal3 s 0 40208 800 40320 0 FreeSans 448 0 0 0 io_wbs_datwr_1[20]
port 274 nsew signal tristate
flabel metal3 s 0 40880 800 40992 0 FreeSans 448 0 0 0 io_wbs_datwr_1[21]
port 275 nsew signal tristate
flabel metal3 s 0 41552 800 41664 0 FreeSans 448 0 0 0 io_wbs_datwr_1[22]
port 276 nsew signal tristate
flabel metal3 s 0 42224 800 42336 0 FreeSans 448 0 0 0 io_wbs_datwr_1[23]
port 277 nsew signal tristate
flabel metal3 s 0 42896 800 43008 0 FreeSans 448 0 0 0 io_wbs_datwr_1[24]
port 278 nsew signal tristate
flabel metal3 s 0 43568 800 43680 0 FreeSans 448 0 0 0 io_wbs_datwr_1[25]
port 279 nsew signal tristate
flabel metal3 s 0 44240 800 44352 0 FreeSans 448 0 0 0 io_wbs_datwr_1[26]
port 280 nsew signal tristate
flabel metal3 s 0 44912 800 45024 0 FreeSans 448 0 0 0 io_wbs_datwr_1[27]
port 281 nsew signal tristate
flabel metal3 s 0 45584 800 45696 0 FreeSans 448 0 0 0 io_wbs_datwr_1[28]
port 282 nsew signal tristate
flabel metal3 s 0 46256 800 46368 0 FreeSans 448 0 0 0 io_wbs_datwr_1[29]
port 283 nsew signal tristate
flabel metal3 s 0 28112 800 28224 0 FreeSans 448 0 0 0 io_wbs_datwr_1[2]
port 284 nsew signal tristate
flabel metal3 s 0 46928 800 47040 0 FreeSans 448 0 0 0 io_wbs_datwr_1[30]
port 285 nsew signal tristate
flabel metal3 s 0 47600 800 47712 0 FreeSans 448 0 0 0 io_wbs_datwr_1[31]
port 286 nsew signal tristate
flabel metal3 s 0 28784 800 28896 0 FreeSans 448 0 0 0 io_wbs_datwr_1[3]
port 287 nsew signal tristate
flabel metal3 s 0 29456 800 29568 0 FreeSans 448 0 0 0 io_wbs_datwr_1[4]
port 288 nsew signal tristate
flabel metal3 s 0 30128 800 30240 0 FreeSans 448 0 0 0 io_wbs_datwr_1[5]
port 289 nsew signal tristate
flabel metal3 s 0 30800 800 30912 0 FreeSans 448 0 0 0 io_wbs_datwr_1[6]
port 290 nsew signal tristate
flabel metal3 s 0 31472 800 31584 0 FreeSans 448 0 0 0 io_wbs_datwr_1[7]
port 291 nsew signal tristate
flabel metal3 s 0 32144 800 32256 0 FreeSans 448 0 0 0 io_wbs_datwr_1[8]
port 292 nsew signal tristate
flabel metal3 s 0 32816 800 32928 0 FreeSans 448 0 0 0 io_wbs_datwr_1[9]
port 293 nsew signal tristate
flabel metal2 s 70448 0 70560 800 0 FreeSans 448 90 0 0 io_wbs_sel[0]
port 294 nsew signal input
flabel metal2 s 71120 0 71232 800 0 FreeSans 448 90 0 0 io_wbs_sel[1]
port 295 nsew signal input
flabel metal2 s 71792 0 71904 800 0 FreeSans 448 90 0 0 io_wbs_sel[2]
port 296 nsew signal input
flabel metal2 s 72464 0 72576 800 0 FreeSans 448 90 0 0 io_wbs_sel[3]
port 297 nsew signal input
flabel metal3 s 79200 70448 80000 70560 0 FreeSans 448 0 0 0 io_wbs_sel_0[0]
port 298 nsew signal tristate
flabel metal3 s 79200 71120 80000 71232 0 FreeSans 448 0 0 0 io_wbs_sel_0[1]
port 299 nsew signal tristate
flabel metal3 s 79200 71792 80000 71904 0 FreeSans 448 0 0 0 io_wbs_sel_0[2]
port 300 nsew signal tristate
flabel metal3 s 79200 72464 80000 72576 0 FreeSans 448 0 0 0 io_wbs_sel_0[3]
port 301 nsew signal tristate
flabel metal3 s 0 70448 800 70560 0 FreeSans 448 0 0 0 io_wbs_sel_1[0]
port 302 nsew signal tristate
flabel metal3 s 0 71120 800 71232 0 FreeSans 448 0 0 0 io_wbs_sel_1[1]
port 303 nsew signal tristate
flabel metal3 s 0 71792 800 71904 0 FreeSans 448 0 0 0 io_wbs_sel_1[2]
port 304 nsew signal tristate
flabel metal3 s 0 72464 800 72576 0 FreeSans 448 0 0 0 io_wbs_sel_1[3]
port 305 nsew signal tristate
flabel metal2 s 73136 0 73248 800 0 FreeSans 448 90 0 0 io_wbs_stb
port 306 nsew signal input
flabel metal3 s 79200 73136 80000 73248 0 FreeSans 448 0 0 0 io_wbs_stb_0
port 307 nsew signal tristate
flabel metal3 s 0 73136 800 73248 0 FreeSans 448 0 0 0 io_wbs_stb_1
port 308 nsew signal tristate
flabel metal2 s 69776 0 69888 800 0 FreeSans 448 90 0 0 io_wbs_we
port 309 nsew signal input
flabel metal3 s 79200 69776 80000 69888 0 FreeSans 448 0 0 0 io_wbs_we_0
port 310 nsew signal tristate
flabel metal3 s 0 69776 800 69888 0 FreeSans 448 0 0 0 io_wbs_we_1
port 311 nsew signal tristate
flabel metal4 s 4448 3076 4768 76892 0 FreeSans 1280 90 0 0 vdd
port 312 nsew power bidirectional
flabel metal4 s 35168 3076 35488 76892 0 FreeSans 1280 90 0 0 vdd
port 312 nsew power bidirectional
flabel metal4 s 65888 3076 66208 76892 0 FreeSans 1280 90 0 0 vdd
port 312 nsew power bidirectional
flabel metal4 s 19808 3076 20128 76892 0 FreeSans 1280 90 0 0 vss
port 313 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 76892 0 FreeSans 1280 90 0 0 vss
port 313 nsew ground bidirectional
rlabel metal1 39984 76048 39984 76048 0 vdd
rlabel metal1 39984 76832 39984 76832 0 vss
rlabel metal2 69496 50176 69496 50176 0 _000_
rlabel metal2 20888 17360 20888 17360 0 _001_
rlabel metal2 26208 16856 26208 16856 0 _002_
rlabel metal2 55272 17136 55272 17136 0 _003_
rlabel metal3 20888 16072 20888 16072 0 _004_
rlabel metal2 22904 16688 22904 16688 0 _005_
rlabel metal2 23240 16800 23240 16800 0 _006_
rlabel metal2 54824 16856 54824 16856 0 _007_
rlabel metal2 55664 17752 55664 17752 0 _008_
rlabel metal2 67480 65016 67480 65016 0 _009_
rlabel metal3 68264 64456 68264 64456 0 _010_
rlabel metal2 69272 72408 69272 72408 0 _011_
rlabel metal2 56224 17864 56224 17864 0 _012_
rlabel metal3 56560 52136 56560 52136 0 _013_
rlabel metal2 62216 64064 62216 64064 0 _014_
rlabel metal2 68488 64736 68488 64736 0 _015_
rlabel metal3 72016 72632 72016 72632 0 _016_
rlabel metal2 70168 50064 70168 50064 0 _017_
rlabel metal3 68992 48776 68992 48776 0 _018_
rlabel metal2 68936 48720 68936 48720 0 _019_
rlabel metal2 48608 48440 48608 48440 0 _020_
rlabel metal3 56560 53704 56560 53704 0 _021_
rlabel metal2 51016 50064 51016 50064 0 _022_
rlabel metal2 56952 55104 56952 55104 0 _023_
rlabel metal2 49728 49672 49728 49672 0 _024_
rlabel metal3 50176 49000 50176 49000 0 _025_
rlabel metal3 49056 49224 49056 49224 0 _026_
rlabel metal2 49672 48440 49672 48440 0 _027_
rlabel metal3 48944 50008 48944 50008 0 _028_
rlabel metal3 51968 49560 51968 49560 0 _029_
rlabel metal3 50232 50456 50232 50456 0 _030_
rlabel metal2 51408 50568 51408 50568 0 _031_
rlabel metal2 48888 51744 48888 51744 0 _032_
rlabel metal3 53592 53144 53592 53144 0 _033_
rlabel metal3 53648 52808 53648 52808 0 _034_
rlabel metal2 52584 51800 52584 51800 0 _035_
rlabel metal3 49672 52024 49672 52024 0 _036_
rlabel metal3 56504 52360 56504 52360 0 _037_
rlabel metal3 50680 52920 50680 52920 0 _038_
rlabel metal3 54992 52696 54992 52696 0 _039_
rlabel metal3 52360 53032 52360 53032 0 _040_
rlabel metal2 53928 53200 53928 53200 0 _041_
rlabel metal3 53480 53704 53480 53704 0 _042_
rlabel metal2 55272 55272 55272 55272 0 _043_
rlabel metal2 55664 55384 55664 55384 0 _044_
rlabel metal2 54264 54096 54264 54096 0 _045_
rlabel metal3 53872 54488 53872 54488 0 _046_
rlabel metal3 55552 54264 55552 54264 0 _047_
rlabel metal3 52920 55048 52920 55048 0 _048_
rlabel metal2 56504 54824 56504 54824 0 _049_
rlabel metal3 53928 56056 53928 56056 0 _050_
rlabel metal2 56056 56224 56056 56224 0 _051_
rlabel metal3 57344 56280 57344 56280 0 _052_
rlabel metal2 57624 57904 57624 57904 0 _053_
rlabel metal2 58072 55552 58072 55552 0 _054_
rlabel metal3 58688 56056 58688 56056 0 _055_
rlabel metal3 56504 57624 56504 57624 0 _056_
rlabel metal3 60480 57400 60480 57400 0 _057_
rlabel metal2 58072 56896 58072 56896 0 _058_
rlabel metal2 58520 57456 58520 57456 0 _059_
rlabel metal3 59304 57680 59304 57680 0 _060_
rlabel metal2 58744 57624 58744 57624 0 _061_
rlabel metal2 59864 59472 59864 59472 0 _062_
rlabel metal2 61040 59416 61040 59416 0 _063_
rlabel metal3 61600 60648 61600 60648 0 _064_
rlabel metal2 60312 59472 60312 59472 0 _065_
rlabel metal3 58856 59864 58856 59864 0 _066_
rlabel metal3 63616 59976 63616 59976 0 _067_
rlabel metal3 59248 60760 59248 60760 0 _068_
rlabel metal3 62944 60536 62944 60536 0 _069_
rlabel metal2 60312 61152 60312 61152 0 _070_
rlabel metal2 61880 61040 61880 61040 0 _071_
rlabel metal3 62104 62552 62104 62552 0 _072_
rlabel metal2 63168 63112 63168 63112 0 _073_
rlabel metal3 63112 63784 63112 63784 0 _074_
rlabel metal2 62664 61936 62664 61936 0 _075_
rlabel metal3 61880 62328 61880 62328 0 _076_
rlabel metal3 66304 62216 66304 62216 0 _077_
rlabel metal2 63336 62832 63336 62832 0 _078_
rlabel metal2 63784 63392 63784 63392 0 _079_
rlabel metal3 62328 64008 62328 64008 0 _080_
rlabel metal2 63840 63784 63840 63784 0 _081_
rlabel metal3 63448 64456 63448 64456 0 _082_
rlabel metal2 65128 64400 65128 64400 0 _083_
rlabel metal2 66136 66416 66136 66416 0 _084_
rlabel metal3 66080 64568 66080 64568 0 _085_
rlabel metal2 61880 65520 61880 65520 0 _086_
rlabel metal2 65072 65240 65072 65240 0 _087_
rlabel metal3 64232 66136 64232 66136 0 _088_
rlabel metal2 66640 66248 66640 66248 0 _089_
rlabel metal2 63448 66752 63448 66752 0 _090_
rlabel metal2 66752 66808 66752 66808 0 _091_
rlabel metal2 67256 67396 67256 67396 0 _092_
rlabel metal2 68544 67368 68544 67368 0 _093_
rlabel metal2 67928 67396 67928 67396 0 _094_
rlabel metal2 69384 67396 69384 67396 0 _095_
rlabel metal2 68152 68376 68152 68376 0 _096_
rlabel metal2 68880 67032 68880 67032 0 _097_
rlabel metal3 71512 71960 71512 71960 0 _098_
rlabel metal3 71624 73416 71624 73416 0 _099_
rlabel metal2 73864 2086 73864 2086 0 io_wbs_ack
rlabel metal3 78120 73920 78120 73920 0 io_wbs_ack_0
rlabel metal2 3640 73920 3640 73920 0 io_wbs_ack_1
rlabel metal2 5208 4200 5208 4200 0 io_wbs_adr[0]
rlabel metal2 11984 3416 11984 3416 0 io_wbs_adr[10]
rlabel metal2 12656 3528 12656 3528 0 io_wbs_adr[11]
rlabel metal2 13272 4200 13272 4200 0 io_wbs_adr[12]
rlabel metal2 14056 2086 14056 2086 0 io_wbs_adr[13]
rlabel metal2 14728 2142 14728 2142 0 io_wbs_adr[14]
rlabel via2 15400 4312 15400 4312 0 io_wbs_adr[15]
rlabel metal2 15848 3080 15848 3080 0 io_wbs_adr[16]
rlabel metal2 16744 2058 16744 2058 0 io_wbs_adr[17]
rlabel via2 17416 4312 17416 4312 0 io_wbs_adr[18]
rlabel metal2 18088 3528 18088 3528 0 io_wbs_adr[19]
rlabel metal2 5992 2142 5992 2142 0 io_wbs_adr[1]
rlabel metal2 18760 2058 18760 2058 0 io_wbs_adr[20]
rlabel metal2 19432 3864 19432 3864 0 io_wbs_adr[21]
rlabel metal2 20104 1862 20104 1862 0 io_wbs_adr[22]
rlabel metal2 20720 3528 20720 3528 0 io_wbs_adr[23]
rlabel via2 21448 4312 21448 4312 0 io_wbs_adr[24]
rlabel metal3 22064 3528 22064 3528 0 io_wbs_adr[25]
rlabel metal2 22848 3528 22848 3528 0 io_wbs_adr[26]
rlabel metal2 23464 3864 23464 3864 0 io_wbs_adr[27]
rlabel via2 24136 4312 24136 4312 0 io_wbs_adr[28]
rlabel metal2 24696 3528 24696 3528 0 io_wbs_adr[29]
rlabel metal2 6440 3976 6440 3976 0 io_wbs_adr[2]
rlabel metal2 25480 854 25480 854 0 io_wbs_adr[30]
rlabel via2 26152 4312 26152 4312 0 io_wbs_adr[31]
rlabel metal2 7224 3416 7224 3416 0 io_wbs_adr[3]
rlabel metal2 8008 2086 8008 2086 0 io_wbs_adr[4]
rlabel metal2 9016 3528 9016 3528 0 io_wbs_adr[5]
rlabel metal3 8960 3416 8960 3416 0 io_wbs_adr[6]
rlabel metal2 10080 3416 10080 3416 0 io_wbs_adr[7]
rlabel metal2 10696 2086 10696 2086 0 io_wbs_adr[8]
rlabel metal2 11256 4200 11256 4200 0 io_wbs_adr[9]
rlabel metal2 76104 5544 76104 5544 0 io_wbs_adr_0[0]
rlabel metal3 77658 12040 77658 12040 0 io_wbs_adr_0[10]
rlabel metal2 77784 12488 77784 12488 0 io_wbs_adr_0[11]
rlabel metal2 76104 13552 76104 13552 0 io_wbs_adr_0[12]
rlabel metal2 77784 13944 77784 13944 0 io_wbs_adr_0[13]
rlabel metal2 76104 14952 76104 14952 0 io_wbs_adr_0[14]
rlabel metal2 76216 15680 76216 15680 0 io_wbs_adr_0[15]
rlabel metal2 77784 15736 77784 15736 0 io_wbs_adr_0[16]
rlabel metal3 75992 16800 75992 16800 0 io_wbs_adr_0[17]
rlabel metal2 77784 17192 77784 17192 0 io_wbs_adr_0[18]
rlabel metal2 76104 18200 76104 18200 0 io_wbs_adr_0[19]
rlabel metal2 76216 6272 76216 6272 0 io_wbs_adr_0[1]
rlabel metal3 77840 18424 77840 18424 0 io_wbs_adr_0[20]
rlabel metal2 76104 19656 76104 19656 0 io_wbs_adr_0[21]
rlabel metal3 76328 20216 76328 20216 0 io_wbs_adr_0[22]
rlabel metal3 78554 20776 78554 20776 0 io_wbs_adr_0[23]
rlabel metal3 77658 21448 77658 21448 0 io_wbs_adr_0[24]
rlabel metal2 77784 21896 77784 21896 0 io_wbs_adr_0[25]
rlabel metal2 76104 22904 76104 22904 0 io_wbs_adr_0[26]
rlabel metal2 77784 23352 77784 23352 0 io_wbs_adr_0[27]
rlabel metal2 76104 24360 76104 24360 0 io_wbs_adr_0[28]
rlabel metal2 76216 25088 76216 25088 0 io_wbs_adr_0[29]
rlabel metal2 77784 6328 77784 6328 0 io_wbs_adr_0[2]
rlabel metal2 77784 25144 77784 25144 0 io_wbs_adr_0[30]
rlabel metal3 77658 26152 77658 26152 0 io_wbs_adr_0[31]
rlabel metal3 77658 7336 77658 7336 0 io_wbs_adr_0[3]
rlabel metal2 77784 7784 77784 7784 0 io_wbs_adr_0[4]
rlabel metal2 76104 8792 76104 8792 0 io_wbs_adr_0[5]
rlabel metal2 77784 9240 77784 9240 0 io_wbs_adr_0[6]
rlabel metal2 76104 10304 76104 10304 0 io_wbs_adr_0[7]
rlabel metal2 76216 10976 76216 10976 0 io_wbs_adr_0[8]
rlabel metal2 77784 11032 77784 11032 0 io_wbs_adr_0[9]
rlabel metal3 1414 5320 1414 5320 0 io_wbs_adr_1[0]
rlabel metal2 2072 11760 2072 11760 0 io_wbs_adr_1[10]
rlabel metal3 1470 12712 1470 12712 0 io_wbs_adr_1[11]
rlabel metal2 2072 13216 2072 13216 0 io_wbs_adr_1[12]
rlabel metal3 1470 14056 1470 14056 0 io_wbs_adr_1[13]
rlabel metal3 1414 14728 1414 14728 0 io_wbs_adr_1[14]
rlabel metal3 1470 15400 1470 15400 0 io_wbs_adr_1[15]
rlabel metal3 2310 16072 2310 16072 0 io_wbs_adr_1[16]
rlabel metal2 2072 16464 2072 16464 0 io_wbs_adr_1[17]
rlabel metal3 1470 17416 1470 17416 0 io_wbs_adr_1[18]
rlabel metal2 2072 17920 2072 17920 0 io_wbs_adr_1[19]
rlabel metal3 1470 5992 1470 5992 0 io_wbs_adr_1[1]
rlabel metal3 1470 18760 1470 18760 0 io_wbs_adr_1[20]
rlabel metal3 1414 19432 1414 19432 0 io_wbs_adr_1[21]
rlabel metal3 1470 20104 1470 20104 0 io_wbs_adr_1[22]
rlabel metal3 2310 20776 2310 20776 0 io_wbs_adr_1[23]
rlabel metal2 2072 21168 2072 21168 0 io_wbs_adr_1[24]
rlabel metal3 1470 22120 1470 22120 0 io_wbs_adr_1[25]
rlabel metal2 2072 22624 2072 22624 0 io_wbs_adr_1[26]
rlabel metal3 1470 23464 1470 23464 0 io_wbs_adr_1[27]
rlabel metal3 1414 24136 1414 24136 0 io_wbs_adr_1[28]
rlabel metal3 1470 24808 1470 24808 0 io_wbs_adr_1[29]
rlabel metal3 2310 6664 2310 6664 0 io_wbs_adr_1[2]
rlabel metal3 2310 25480 2310 25480 0 io_wbs_adr_1[30]
rlabel metal2 2072 25872 2072 25872 0 io_wbs_adr_1[31]
rlabel metal2 2184 7000 2184 7000 0 io_wbs_adr_1[3]
rlabel metal3 1470 8008 1470 8008 0 io_wbs_adr_1[4]
rlabel metal3 1414 8680 1414 8680 0 io_wbs_adr_1[5]
rlabel metal3 1470 9352 1470 9352 0 io_wbs_adr_1[6]
rlabel metal3 1414 10024 1414 10024 0 io_wbs_adr_1[7]
rlabel metal3 1470 10696 1470 10696 0 io_wbs_adr_1[8]
rlabel metal3 2310 11368 2310 11368 0 io_wbs_adr_1[9]
rlabel metal2 75432 2520 75432 2520 0 io_wbs_cyc
rlabel metal2 76104 74648 76104 74648 0 io_wbs_cyc_0
rlabel metal3 1414 74536 1414 74536 0 io_wbs_cyc_1
rlabel metal3 48776 3416 48776 3416 0 io_wbs_datrd[0]
rlabel metal2 55048 2982 55048 2982 0 io_wbs_datrd[10]
rlabel metal2 55720 2142 55720 2142 0 io_wbs_datrd[11]
rlabel metal2 56392 2086 56392 2086 0 io_wbs_datrd[12]
rlabel metal2 57064 2982 57064 2982 0 io_wbs_datrd[13]
rlabel metal2 57736 2478 57736 2478 0 io_wbs_datrd[14]
rlabel metal2 58408 2198 58408 2198 0 io_wbs_datrd[15]
rlabel metal2 59080 1694 59080 1694 0 io_wbs_datrd[16]
rlabel metal2 59752 2142 59752 2142 0 io_wbs_datrd[17]
rlabel metal2 60424 2086 60424 2086 0 io_wbs_datrd[18]
rlabel metal2 61096 1638 61096 1638 0 io_wbs_datrd[19]
rlabel metal3 49616 4200 49616 4200 0 io_wbs_datrd[1]
rlabel metal2 61768 2478 61768 2478 0 io_wbs_datrd[20]
rlabel metal2 62440 1246 62440 1246 0 io_wbs_datrd[21]
rlabel metal2 63112 1638 63112 1638 0 io_wbs_datrd[22]
rlabel metal2 63784 2478 63784 2478 0 io_wbs_datrd[23]
rlabel metal2 64456 2142 64456 2142 0 io_wbs_datrd[24]
rlabel metal2 65128 2982 65128 2982 0 io_wbs_datrd[25]
rlabel metal2 67928 3864 67928 3864 0 io_wbs_datrd[26]
rlabel metal2 66472 2086 66472 2086 0 io_wbs_datrd[27]
rlabel metal2 67144 2982 67144 2982 0 io_wbs_datrd[28]
rlabel metal2 67816 2478 67816 2478 0 io_wbs_datrd[29]
rlabel metal2 49672 2086 49672 2086 0 io_wbs_datrd[2]
rlabel metal2 68488 1246 68488 1246 0 io_wbs_datrd[30]
rlabel metal2 69160 1694 69160 1694 0 io_wbs_datrd[31]
rlabel metal2 52136 3864 52136 3864 0 io_wbs_datrd[3]
rlabel metal2 51016 2198 51016 2198 0 io_wbs_datrd[4]
rlabel metal2 51688 2254 51688 2254 0 io_wbs_datrd[5]
rlabel metal2 52360 2086 52360 2086 0 io_wbs_datrd[6]
rlabel metal2 53032 1694 53032 1694 0 io_wbs_datrd[7]
rlabel metal2 53704 2478 53704 2478 0 io_wbs_datrd[8]
rlabel metal2 54376 2198 54376 2198 0 io_wbs_datrd[9]
rlabel metal2 78120 48608 78120 48608 0 io_wbs_datrd_0[0]
rlabel metal3 79128 55384 79128 55384 0 io_wbs_datrd_0[10]
rlabel metal2 78008 56280 78008 56280 0 io_wbs_datrd_0[11]
rlabel metal2 78120 57008 78120 57008 0 io_wbs_datrd_0[12]
rlabel metal2 78008 57848 78008 57848 0 io_wbs_datrd_0[13]
rlabel metal2 78120 58520 78120 58520 0 io_wbs_datrd_0[14]
rlabel metal2 78008 59416 78008 59416 0 io_wbs_datrd_0[15]
rlabel metal2 77224 59136 77224 59136 0 io_wbs_datrd_0[16]
rlabel metal2 78120 60312 78120 60312 0 io_wbs_datrd_0[17]
rlabel metal2 78176 61432 78176 61432 0 io_wbs_datrd_0[18]
rlabel metal2 78008 61712 78008 61712 0 io_wbs_datrd_0[19]
rlabel metal2 78008 49392 78008 49392 0 io_wbs_datrd_0[1]
rlabel metal2 78120 62384 78120 62384 0 io_wbs_datrd_0[20]
rlabel metal2 78008 63224 78008 63224 0 io_wbs_datrd_0[21]
rlabel metal2 78120 63896 78120 63896 0 io_wbs_datrd_0[22]
rlabel metal3 77224 63840 77224 63840 0 io_wbs_datrd_0[23]
rlabel metal2 78008 64960 78008 64960 0 io_wbs_datrd_0[24]
rlabel metal2 78120 65632 78120 65632 0 io_wbs_datrd_0[25]
rlabel metal2 78176 67032 78176 67032 0 io_wbs_datrd_0[26]
rlabel metal3 77672 67816 77672 67816 0 io_wbs_datrd_0[27]
rlabel metal3 77000 68600 77000 68600 0 io_wbs_datrd_0[28]
rlabel metal2 78176 69272 78176 69272 0 io_wbs_datrd_0[29]
rlabel metal2 78120 50120 78120 50120 0 io_wbs_datrd_0[2]
rlabel metal2 77224 68544 77224 68544 0 io_wbs_datrd_0[30]
rlabel metal3 78274 69160 78274 69160 0 io_wbs_datrd_0[31]
rlabel metal2 78008 50904 78008 50904 0 io_wbs_datrd_0[3]
rlabel metal2 78120 51520 78120 51520 0 io_wbs_datrd_0[4]
rlabel metal2 78008 52304 78008 52304 0 io_wbs_datrd_0[5]
rlabel metal2 78120 52976 78120 52976 0 io_wbs_datrd_0[6]
rlabel metal2 78176 54488 78176 54488 0 io_wbs_datrd_0[7]
rlabel metal2 78008 54544 78008 54544 0 io_wbs_datrd_0[8]
rlabel metal2 77224 54432 77224 54432 0 io_wbs_datrd_0[9]
rlabel metal2 1848 49056 1848 49056 0 io_wbs_datrd_1[0]
rlabel metal3 1358 55048 1358 55048 0 io_wbs_datrd_1[10]
rlabel metal2 1848 56224 1848 56224 0 io_wbs_datrd_1[11]
rlabel metal2 1960 57008 1960 57008 0 io_wbs_datrd_1[12]
rlabel metal2 1848 57680 1848 57680 0 io_wbs_datrd_1[13]
rlabel metal2 1960 58520 1960 58520 0 io_wbs_datrd_1[14]
rlabel metal2 1792 59864 1792 59864 0 io_wbs_datrd_1[15]
rlabel metal2 2744 59136 2744 59136 0 io_wbs_datrd_1[16]
rlabel metal2 1960 60256 1960 60256 0 io_wbs_datrd_1[17]
rlabel metal2 1792 61432 1792 61432 0 io_wbs_datrd_1[18]
rlabel metal2 1960 61712 1960 61712 0 io_wbs_datrd_1[19]
rlabel metal2 1792 50456 1792 50456 0 io_wbs_datrd_1[1]
rlabel metal2 1848 62384 1848 62384 0 io_wbs_datrd_1[20]
rlabel metal2 1960 63224 1960 63224 0 io_wbs_datrd_1[21]
rlabel metal2 1792 64568 1792 64568 0 io_wbs_datrd_1[22]
rlabel metal2 2744 63840 2744 63840 0 io_wbs_datrd_1[23]
rlabel metal2 1960 64960 1960 64960 0 io_wbs_datrd_1[24]
rlabel metal2 1848 65632 1848 65632 0 io_wbs_datrd_1[25]
rlabel metal2 1960 66416 1960 66416 0 io_wbs_datrd_1[26]
rlabel metal3 1302 66472 1302 66472 0 io_wbs_datrd_1[27]
rlabel metal3 2744 68600 2744 68600 0 io_wbs_datrd_1[28]
rlabel metal2 1848 68600 1848 68600 0 io_wbs_datrd_1[29]
rlabel metal2 2744 49728 2744 49728 0 io_wbs_datrd_1[2]
rlabel metal2 2744 68544 2744 68544 0 io_wbs_datrd_1[30]
rlabel metal2 2744 69216 2744 69216 0 io_wbs_datrd_1[31]
rlabel metal2 1960 50848 1960 50848 0 io_wbs_datrd_1[3]
rlabel metal2 1848 51520 1848 51520 0 io_wbs_datrd_1[4]
rlabel metal2 1960 52304 1960 52304 0 io_wbs_datrd_1[5]
rlabel metal2 1848 52976 1848 52976 0 io_wbs_datrd_1[6]
rlabel metal2 1960 53816 1960 53816 0 io_wbs_datrd_1[7]
rlabel metal2 1792 55160 1792 55160 0 io_wbs_datrd_1[8]
rlabel metal2 2744 54432 2744 54432 0 io_wbs_datrd_1[9]
rlabel metal2 26768 3528 26768 3528 0 io_wbs_datwr[0]
rlabel metal2 33600 3416 33600 3416 0 io_wbs_datwr[10]
rlabel metal2 34216 2086 34216 2086 0 io_wbs_datwr[11]
rlabel metal2 34776 4200 34776 4200 0 io_wbs_datwr[12]
rlabel metal2 35504 3416 35504 3416 0 io_wbs_datwr[13]
rlabel metal2 36232 2142 36232 2142 0 io_wbs_datwr[14]
rlabel metal2 36792 4200 36792 4200 0 io_wbs_datwr[15]
rlabel metal2 37576 2086 37576 2086 0 io_wbs_datwr[16]
rlabel metal2 38248 2142 38248 2142 0 io_wbs_datwr[17]
rlabel via2 38920 4312 38920 4312 0 io_wbs_datwr[18]
rlabel metal2 39760 4200 39760 4200 0 io_wbs_datwr[19]
rlabel metal2 27496 2142 27496 2142 0 io_wbs_datwr[1]
rlabel metal2 40320 3528 40320 3528 0 io_wbs_datwr[20]
rlabel metal3 41272 4312 41272 4312 0 io_wbs_datwr[21]
rlabel metal2 41608 2058 41608 2058 0 io_wbs_datwr[22]
rlabel metal2 42280 2058 42280 2058 0 io_wbs_datwr[23]
rlabel metal3 43288 3528 43288 3528 0 io_wbs_datwr[24]
rlabel metal2 43568 3192 43568 3192 0 io_wbs_datwr[25]
rlabel metal2 44968 3864 44968 3864 0 io_wbs_datwr[26]
rlabel metal2 45024 2856 45024 2856 0 io_wbs_datwr[27]
rlabel metal2 45696 2744 45696 2744 0 io_wbs_datwr[28]
rlabel metal2 46200 2856 46200 2856 0 io_wbs_datwr[29]
rlabel metal2 28168 2086 28168 2086 0 io_wbs_datwr[2]
rlabel metal2 47992 3864 47992 3864 0 io_wbs_datwr[30]
rlabel metal2 47768 3080 47768 3080 0 io_wbs_datwr[31]
rlabel metal2 28728 4200 28728 4200 0 io_wbs_datwr[3]
rlabel metal2 29624 3136 29624 3136 0 io_wbs_datwr[4]
rlabel metal2 30072 4200 30072 4200 0 io_wbs_datwr[5]
rlabel metal2 30744 3416 30744 3416 0 io_wbs_datwr[6]
rlabel metal2 31528 2086 31528 2086 0 io_wbs_datwr[7]
rlabel metal2 31976 3528 31976 3528 0 io_wbs_datwr[8]
rlabel metal2 32424 3080 32424 3080 0 io_wbs_datwr[9]
rlabel metal2 77784 26600 77784 26600 0 io_wbs_datwr_0[0]
rlabel metal2 76104 33824 76104 33824 0 io_wbs_datwr_0[10]
rlabel metal2 76216 34496 76216 34496 0 io_wbs_datwr_0[11]
rlabel metal2 77784 34552 77784 34552 0 io_wbs_datwr_0[12]
rlabel metal3 77658 35560 77658 35560 0 io_wbs_datwr_0[13]
rlabel metal2 77784 36008 77784 36008 0 io_wbs_datwr_0[14]
rlabel metal2 76104 37072 76104 37072 0 io_wbs_datwr_0[15]
rlabel metal2 77784 37464 77784 37464 0 io_wbs_datwr_0[16]
rlabel metal2 76104 38472 76104 38472 0 io_wbs_datwr_0[17]
rlabel metal2 76216 39200 76216 39200 0 io_wbs_datwr_0[18]
rlabel metal2 77784 39256 77784 39256 0 io_wbs_datwr_0[19]
rlabel metal2 76104 27608 76104 27608 0 io_wbs_datwr_0[1]
rlabel metal3 75992 40320 75992 40320 0 io_wbs_datwr_0[20]
rlabel metal2 77784 40712 77784 40712 0 io_wbs_datwr_0[21]
rlabel metal2 76104 41720 76104 41720 0 io_wbs_datwr_0[22]
rlabel metal3 77840 41944 77840 41944 0 io_wbs_datwr_0[23]
rlabel metal2 77896 43176 77896 43176 0 io_wbs_datwr_0[24]
rlabel metal2 77896 44352 77896 44352 0 io_wbs_datwr_0[25]
rlabel metal2 76104 44632 76104 44632 0 io_wbs_datwr_0[26]
rlabel metal2 77784 45752 77784 45752 0 io_wbs_datwr_0[27]
rlabel metal2 76216 45696 76216 45696 0 io_wbs_datwr_0[28]
rlabel metal2 76104 46424 76104 46424 0 io_wbs_datwr_0[29]
rlabel metal2 77784 28056 77784 28056 0 io_wbs_datwr_0[2]
rlabel metal2 77896 47600 77896 47600 0 io_wbs_datwr_0[30]
rlabel metal2 76104 47880 76104 47880 0 io_wbs_datwr_0[31]
rlabel metal2 76104 29064 76104 29064 0 io_wbs_datwr_0[3]
rlabel metal2 76216 29792 76216 29792 0 io_wbs_datwr_0[4]
rlabel metal2 77784 29848 77784 29848 0 io_wbs_datwr_0[5]
rlabel metal3 77658 30856 77658 30856 0 io_wbs_datwr_0[6]
rlabel metal2 77784 31304 77784 31304 0 io_wbs_datwr_0[7]
rlabel metal2 76104 32312 76104 32312 0 io_wbs_datwr_0[8]
rlabel metal2 77784 32760 77784 32760 0 io_wbs_datwr_0[9]
rlabel metal3 1470 26824 1470 26824 0 io_wbs_datwr_1[0]
rlabel metal3 1414 33544 1414 33544 0 io_wbs_datwr_1[10]
rlabel metal3 1470 34216 1470 34216 0 io_wbs_datwr_1[11]
rlabel metal3 2310 34888 2310 34888 0 io_wbs_datwr_1[12]
rlabel metal2 2072 35280 2072 35280 0 io_wbs_datwr_1[13]
rlabel metal3 1470 36232 1470 36232 0 io_wbs_datwr_1[14]
rlabel metal2 2072 36736 2072 36736 0 io_wbs_datwr_1[15]
rlabel metal3 1470 37576 1470 37576 0 io_wbs_datwr_1[16]
rlabel metal3 1414 38248 1414 38248 0 io_wbs_datwr_1[17]
rlabel metal3 1470 38920 1470 38920 0 io_wbs_datwr_1[18]
rlabel metal3 1470 39592 1470 39592 0 io_wbs_datwr_1[19]
rlabel metal2 2072 27328 2072 27328 0 io_wbs_datwr_1[1]
rlabel metal3 1414 40264 1414 40264 0 io_wbs_datwr_1[20]
rlabel metal3 1470 40936 1470 40936 0 io_wbs_datwr_1[21]
rlabel metal3 1414 41608 1414 41608 0 io_wbs_datwr_1[22]
rlabel metal3 1470 42280 1470 42280 0 io_wbs_datwr_1[23]
rlabel metal3 1414 42952 1414 42952 0 io_wbs_datwr_1[24]
rlabel metal3 1470 43624 1470 43624 0 io_wbs_datwr_1[25]
rlabel metal3 1414 44296 1414 44296 0 io_wbs_datwr_1[26]
rlabel metal3 1470 44968 1470 44968 0 io_wbs_datwr_1[27]
rlabel metal3 1414 45640 1414 45640 0 io_wbs_datwr_1[28]
rlabel metal3 1470 46312 1470 46312 0 io_wbs_datwr_1[29]
rlabel metal3 1470 28168 1470 28168 0 io_wbs_datwr_1[2]
rlabel metal3 1414 46984 1414 46984 0 io_wbs_datwr_1[30]
rlabel metal3 1470 47656 1470 47656 0 io_wbs_datwr_1[31]
rlabel metal3 1414 28840 1414 28840 0 io_wbs_datwr_1[3]
rlabel metal3 1470 29512 1470 29512 0 io_wbs_datwr_1[4]
rlabel metal3 2310 30184 2310 30184 0 io_wbs_datwr_1[5]
rlabel metal2 2184 30520 2184 30520 0 io_wbs_datwr_1[6]
rlabel metal3 1470 31528 1470 31528 0 io_wbs_datwr_1[7]
rlabel metal3 1414 32200 1414 32200 0 io_wbs_datwr_1[8]
rlabel metal3 1470 32872 1470 32872 0 io_wbs_datwr_1[9]
rlabel metal3 71624 3416 71624 3416 0 io_wbs_sel[0]
rlabel metal3 71624 4312 71624 4312 0 io_wbs_sel[1]
rlabel metal2 71624 4088 71624 4088 0 io_wbs_sel[2]
rlabel metal2 73416 3640 73416 3640 0 io_wbs_sel[3]
rlabel metal2 77896 71120 77896 71120 0 io_wbs_sel_0[0]
rlabel metal2 76104 71400 76104 71400 0 io_wbs_sel_0[1]
rlabel metal2 77896 72520 77896 72520 0 io_wbs_sel_0[2]
rlabel metal2 76104 72856 76104 72856 0 io_wbs_sel_0[3]
rlabel metal3 1470 70504 1470 70504 0 io_wbs_sel_1[0]
rlabel metal3 1414 71176 1414 71176 0 io_wbs_sel_1[1]
rlabel metal3 1470 71848 1470 71848 0 io_wbs_sel_1[2]
rlabel metal3 1414 72520 1414 72520 0 io_wbs_sel_1[3]
rlabel metal3 74032 4312 74032 4312 0 io_wbs_stb
rlabel metal2 77896 74088 77896 74088 0 io_wbs_stb_0
rlabel metal3 1470 73192 1470 73192 0 io_wbs_stb_1
rlabel metal3 70336 4312 70336 4312 0 io_wbs_we
rlabel metal2 77896 69944 77896 69944 0 io_wbs_we_0
rlabel metal3 1414 69832 1414 69832 0 io_wbs_we_1
rlabel metal2 77672 73864 77672 73864 0 net1
rlabel metal2 16072 15568 16072 15568 0 net10
rlabel metal3 26824 25368 26824 25368 0 net100
rlabel metal2 33320 17612 33320 17612 0 net101
rlabel metal2 34552 5852 34552 5852 0 net102
rlabel metal2 35504 4536 35504 4536 0 net103
rlabel metal3 35616 3304 35616 3304 0 net104
rlabel metal2 36792 34272 36792 34272 0 net105
rlabel metal2 37464 18228 37464 18228 0 net106
rlabel metal3 36904 37128 36904 37128 0 net107
rlabel metal2 38640 37128 38640 37128 0 net108
rlabel metal2 39592 35364 39592 35364 0 net109
rlabel metal3 17080 15176 17080 15176 0 net11
rlabel metal3 39424 39480 39424 39480 0 net110
rlabel metal3 26880 26936 26880 26936 0 net111
rlabel metal2 39984 3304 39984 3304 0 net112
rlabel metal2 41384 35644 41384 35644 0 net113
rlabel metal3 42504 40936 42504 40936 0 net114
rlabel metal2 42896 41944 42896 41944 0 net115
rlabel metal2 44128 42504 44128 42504 0 net116
rlabel metal2 44240 43512 44240 43512 0 net117
rlabel metal3 44352 44184 44352 44184 0 net118
rlabel metal3 44296 45080 44296 45080 0 net119
rlabel metal2 18144 15176 18144 15176 0 net12
rlabel metal2 47208 44968 47208 44968 0 net120
rlabel metal3 46536 45752 46536 45752 0 net121
rlabel metal2 28560 27832 28560 27832 0 net122
rlabel metal2 47600 3304 47600 3304 0 net123
rlabel via2 47880 47320 47880 47320 0 net124
rlabel metal2 29344 4536 29344 4536 0 net125
rlabel metal2 29456 3304 29456 3304 0 net126
rlabel metal2 30688 4536 30688 4536 0 net127
rlabel metal2 31136 29288 31136 29288 0 net128
rlabel metal2 31192 5852 31192 5852 0 net129
rlabel metal2 18536 16576 18536 16576 0 net13
rlabel metal2 32816 4536 32816 4536 0 net130
rlabel metal2 32088 5852 32088 5852 0 net131
rlabel metal3 71568 3304 71568 3304 0 net132
rlabel metal2 71792 70952 71792 70952 0 net133
rlabel metal3 72576 71736 72576 71736 0 net134
rlabel metal3 73416 72520 73416 72520 0 net135
rlabel metal3 73920 4536 73920 4536 0 net136
rlabel metal3 70784 4536 70784 4536 0 net137
rlabel metal2 74424 5320 74424 5320 0 net138
rlabel metal2 74648 5320 74648 5320 0 net139
rlabel metal2 6384 5880 6384 5880 0 net14
rlabel metal2 74648 11648 74648 11648 0 net140
rlabel metal2 76888 12208 76888 12208 0 net141
rlabel metal3 74872 13720 74872 13720 0 net142
rlabel metal2 76888 13776 76888 13776 0 net143
rlabel metal2 75096 15232 75096 15232 0 net144
rlabel metal2 74760 15624 74760 15624 0 net145
rlabel metal2 76888 15568 76888 15568 0 net146
rlabel metal2 74592 17080 74592 17080 0 net147
rlabel metal2 76888 16912 76888 16912 0 net148
rlabel metal2 74648 18088 74648 18088 0 net149
rlabel metal2 20552 18144 20552 18144 0 net15
rlabel metal2 74760 6216 74760 6216 0 net150
rlabel metal2 21112 18088 21112 18088 0 net151
rlabel metal2 74648 19488 74648 19488 0 net152
rlabel metal2 74704 20552 74704 20552 0 net153
rlabel metal2 21224 20048 21224 20048 0 net154
rlabel metal2 74592 21448 74592 21448 0 net155
rlabel metal2 76888 21616 76888 21616 0 net156
rlabel metal2 74648 22568 74648 22568 0 net157
rlabel metal2 76888 23184 76888 23184 0 net158
rlabel metal2 74648 24192 74648 24192 0 net159
rlabel metal2 21616 18648 21616 18648 0 net16
rlabel metal2 74760 25032 74760 25032 0 net160
rlabel metal2 76888 6160 76888 6160 0 net161
rlabel metal2 76664 24360 76664 24360 0 net162
rlabel metal2 74648 25704 74648 25704 0 net163
rlabel metal2 74648 6944 74648 6944 0 net164
rlabel metal2 76888 7504 76888 7504 0 net165
rlabel metal2 74872 9016 74872 9016 0 net166
rlabel metal2 76776 9016 76776 9016 0 net167
rlabel metal2 74648 10024 74648 10024 0 net168
rlabel metal2 74760 10976 74760 10976 0 net169
rlabel metal2 21784 19376 21784 19376 0 net17
rlabel metal2 76888 10864 76888 10864 0 net170
rlabel metal3 3864 4984 3864 4984 0 net171
rlabel metal2 3080 11424 3080 11424 0 net172
rlabel metal2 3080 12208 3080 12208 0 net173
rlabel metal2 3080 12824 3080 12824 0 net174
rlabel metal2 3080 13664 3080 13664 0 net175
rlabel metal2 3080 14392 3080 14392 0 net176
rlabel metal2 3080 15232 3080 15232 0 net177
rlabel metal3 5152 16856 5152 16856 0 net178
rlabel metal2 3080 15960 3080 15960 0 net179
rlabel metal2 20272 17640 20272 17640 0 net18
rlabel metal2 3080 16912 3080 16912 0 net180
rlabel metal2 3080 17528 3080 17528 0 net181
rlabel metal2 3080 5936 3080 5936 0 net182
rlabel metal2 3080 18368 3080 18368 0 net183
rlabel metal2 3640 18928 3640 18928 0 net184
rlabel metal2 3080 19936 3080 19936 0 net185
rlabel metal2 4872 21504 4872 21504 0 net186
rlabel metal2 3080 20720 3080 20720 0 net187
rlabel metal2 2968 21056 2968 21056 0 net188
rlabel metal2 3080 22288 3080 22288 0 net189
rlabel metal2 22008 20412 22008 20412 0 net19
rlabel metal2 3080 23072 3080 23072 0 net190
rlabel metal2 3080 23800 3080 23800 0 net191
rlabel metal2 3080 24640 3080 24640 0 net192
rlabel metal3 5432 6552 5432 6552 0 net193
rlabel metal2 4872 26208 4872 26208 0 net194
rlabel metal2 3080 25424 3080 25424 0 net195
rlabel metal2 3080 6720 3080 6720 0 net196
rlabel metal2 3080 7504 3080 7504 0 net197
rlabel metal3 5544 8120 5544 8120 0 net198
rlabel metal2 3080 9072 3080 9072 0 net199
rlabel metal2 4088 73864 4088 73864 0 net2
rlabel metal3 22176 20552 22176 20552 0 net20
rlabel metal2 3080 9744 3080 9744 0 net200
rlabel metal2 3080 10640 3080 10640 0 net201
rlabel metal2 4872 11704 4872 11704 0 net202
rlabel metal2 73752 74200 73752 74200 0 net203
rlabel metal3 4480 74760 4480 74760 0 net204
rlabel metal2 69272 7084 69272 7084 0 net205
rlabel metal2 55160 6104 55160 6104 0 net206
rlabel metal3 54600 14224 54600 14224 0 net207
rlabel metal2 58184 6216 58184 6216 0 net208
rlabel metal2 58632 5096 58632 5096 0 net209
rlabel metal2 22456 21840 22456 21840 0 net21
rlabel metal3 58464 6104 58464 6104 0 net210
rlabel metal2 60312 6384 60312 6384 0 net211
rlabel metal3 60480 6104 60480 6104 0 net212
rlabel metal2 61656 6160 61656 6160 0 net213
rlabel metal2 62104 6216 62104 6216 0 net214
rlabel metal2 61320 5096 61320 5096 0 net215
rlabel metal2 49280 31920 49280 31920 0 net216
rlabel metal3 63168 4312 63168 4312 0 net217
rlabel metal2 64232 6160 64232 6160 0 net218
rlabel metal3 64064 5096 64064 5096 0 net219
rlabel metal2 23744 23128 23744 23128 0 net22
rlabel metal2 65800 6216 65800 6216 0 net220
rlabel metal2 66192 6104 66192 6104 0 net221
rlabel metal2 66808 6160 66808 6160 0 net222
rlabel metal2 67704 6384 67704 6384 0 net223
rlabel metal2 68152 4648 68152 4648 0 net224
rlabel metal2 67312 5768 67312 5768 0 net225
rlabel metal2 69496 6160 69496 6160 0 net226
rlabel metal2 50904 4368 50904 4368 0 net227
rlabel metal2 71288 3976 71288 3976 0 net228
rlabel metal3 68768 6104 68768 6104 0 net229
rlabel metal2 24024 23408 24024 23408 0 net23
rlabel metal2 51240 4312 51240 4312 0 net230
rlabel metal2 52752 3528 52752 3528 0 net231
rlabel metal2 52192 5208 52192 5208 0 net232
rlabel metal3 53480 6104 53480 6104 0 net233
rlabel metal2 53480 5320 53480 5320 0 net234
rlabel metal2 54432 14280 54432 14280 0 net235
rlabel metal2 54936 7252 54936 7252 0 net236
rlabel metal2 76888 26320 76888 26320 0 net237
rlabel metal2 74648 33544 74648 33544 0 net238
rlabel metal2 74760 34496 74760 34496 0 net239
rlabel metal2 25648 23016 25648 23016 0 net24
rlabel metal2 76888 34384 76888 34384 0 net240
rlabel metal2 74648 35168 74648 35168 0 net241
rlabel metal2 76888 35728 76888 35728 0 net242
rlabel metal2 74648 36680 74648 36680 0 net243
rlabel metal2 76888 37296 76888 37296 0 net244
rlabel metal2 74648 38248 74648 38248 0 net245
rlabel metal2 74760 39200 74760 39200 0 net246
rlabel metal2 76888 39088 76888 39088 0 net247
rlabel metal2 74648 27272 74648 27272 0 net248
rlabel metal2 74648 39928 74648 39928 0 net249
rlabel metal2 6888 5544 6888 5544 0 net25
rlabel metal2 76888 40432 76888 40432 0 net250
rlabel metal2 74648 41440 74648 41440 0 net251
rlabel metal2 76776 41944 76776 41944 0 net252
rlabel metal2 76440 42952 76440 42952 0 net253
rlabel metal2 76552 43904 76552 43904 0 net254
rlabel metal2 74648 44576 74648 44576 0 net255
rlabel metal2 77112 45360 77112 45360 0 net256
rlabel metal2 46536 45472 46536 45472 0 net257
rlabel metal2 74648 46144 74648 46144 0 net258
rlabel metal2 76888 27888 76888 27888 0 net259
rlabel metal2 25928 24080 25928 24080 0 net26
rlabel metal2 77000 47488 77000 47488 0 net260
rlabel metal2 74648 47656 74648 47656 0 net261
rlabel metal2 74648 28840 74648 28840 0 net262
rlabel metal2 74760 29792 74760 29792 0 net263
rlabel metal2 76888 29680 76888 29680 0 net264
rlabel metal2 74648 30464 74648 30464 0 net265
rlabel metal2 76888 31024 76888 31024 0 net266
rlabel metal2 74872 32536 74872 32536 0 net267
rlabel metal2 76776 32536 76776 32536 0 net268
rlabel metal2 2968 25760 2968 25760 0 net269
rlabel metal2 26600 24528 26600 24528 0 net27
rlabel metal2 3080 33208 3080 33208 0 net270
rlabel metal2 3640 33936 3640 33936 0 net271
rlabel metal2 4872 35616 4872 35616 0 net272
rlabel metal2 3080 34776 3080 34776 0 net273
rlabel metal2 3080 35728 3080 35728 0 net274
rlabel metal2 3080 36344 3080 36344 0 net275
rlabel metal2 3640 37072 3640 37072 0 net276
rlabel metal2 3080 37912 3080 37912 0 net277
rlabel metal3 3360 38808 3360 38808 0 net278
rlabel metal2 3080 39536 3080 39536 0 net279
rlabel metal2 6944 7448 6944 7448 0 net28
rlabel metal3 3360 27048 3360 27048 0 net280
rlabel metal3 3360 40376 3360 40376 0 net281
rlabel metal2 3080 41048 3080 41048 0 net282
rlabel metal2 3080 41888 3080 41888 0 net283
rlabel metal2 3080 42616 3080 42616 0 net284
rlabel metal2 3080 43456 3080 43456 0 net285
rlabel metal2 3080 44184 3080 44184 0 net286
rlabel metal2 3080 45024 3080 45024 0 net287
rlabel metal2 3528 45472 3528 45472 0 net288
rlabel metal2 3640 45864 3640 45864 0 net289
rlabel metal2 7672 6776 7672 6776 0 net29
rlabel metal2 3528 46536 3528 46536 0 net290
rlabel metal2 3080 27776 3080 27776 0 net291
rlabel metal2 3696 48104 3696 48104 0 net292
rlabel metal2 3528 48328 3528 48328 0 net293
rlabel metal3 3360 28616 3360 28616 0 net294
rlabel metal2 3640 29232 3640 29232 0 net295
rlabel metal2 4872 30912 4872 30912 0 net296
rlabel metal2 3080 30072 3080 30072 0 net297
rlabel metal2 3080 31024 3080 31024 0 net298
rlabel metal2 3080 31640 3080 31640 0 net299
rlabel metal3 5376 4984 5376 4984 0 net3
rlabel metal3 9464 8120 9464 8120 0 net30
rlabel metal2 3640 32368 3640 32368 0 net300
rlabel metal2 71288 70504 71288 70504 0 net301
rlabel metal3 73528 70840 73528 70840 0 net302
rlabel metal2 72520 72128 72520 72128 0 net303
rlabel metal2 73304 72856 73304 72856 0 net304
rlabel metal2 3528 70504 3528 70504 0 net305
rlabel metal2 3080 71680 3080 71680 0 net306
rlabel metal2 3528 72072 3528 72072 0 net307
rlabel metal2 3080 73248 3080 73248 0 net308
rlabel metal2 74088 73304 74088 73304 0 net309
rlabel metal2 8904 5852 8904 5852 0 net31
rlabel metal2 4368 73976 4368 73976 0 net310
rlabel metal3 73752 69272 73752 69272 0 net311
rlabel metal2 3080 70112 3080 70112 0 net312
rlabel metal2 9744 3304 9744 3304 0 net32
rlabel metal2 11088 10584 11088 10584 0 net33
rlabel metal2 11648 11256 11648 11256 0 net34
rlabel metal2 74200 71176 74200 71176 0 net35
rlabel metal2 77784 48608 77784 48608 0 net36
rlabel metal2 56280 55608 56280 55608 0 net37
rlabel metal2 77840 56616 77840 56616 0 net38
rlabel metal2 77672 56896 77672 56896 0 net39
rlabel metal2 11648 3304 11648 3304 0 net4
rlabel metal2 59808 56616 59808 56616 0 net40
rlabel metal2 77896 58464 77896 58464 0 net41
rlabel metal2 77672 59136 77672 59136 0 net42
rlabel metal2 76888 58856 76888 58856 0 net43
rlabel metal2 77784 60536 77784 60536 0 net44
rlabel metal2 77672 60704 77672 60704 0 net45
rlabel metal3 71568 62440 71568 62440 0 net46
rlabel metal2 50568 48832 50568 48832 0 net47
rlabel metal2 77896 62104 77896 62104 0 net48
rlabel metal2 77448 62776 77448 62776 0 net49
rlabel metal2 12824 5852 12824 5852 0 net5
rlabel metal3 73248 62552 73248 62552 0 net50
rlabel metal2 76888 64176 76888 64176 0 net51
rlabel metal2 77784 65128 77784 65128 0 net52
rlabel metal2 77784 65912 77784 65912 0 net53
rlabel metal2 77784 66696 77784 66696 0 net54
rlabel metal2 77840 67592 77840 67592 0 net55
rlabel metal2 77728 68712 77728 68712 0 net56
rlabel metal2 70056 67984 70056 67984 0 net57
rlabel metal2 50344 48944 50344 48944 0 net58
rlabel metal3 73192 67928 73192 67928 0 net59
rlabel metal3 12432 13720 12432 13720 0 net6
rlabel metal3 72464 68712 72464 68712 0 net60
rlabel metal2 52752 49672 52752 49672 0 net61
rlabel metal2 77672 51240 77672 51240 0 net62
rlabel metal2 77784 52584 77784 52584 0 net63
rlabel metal2 77672 52864 77672 52864 0 net64
rlabel metal2 56952 54152 56952 54152 0 net65
rlabel metal2 77672 54376 77672 54376 0 net66
rlabel metal2 53816 54656 53816 54656 0 net67
rlabel metal3 51688 49784 51688 49784 0 net68
rlabel metal2 2072 55076 2072 55076 0 net69
rlabel metal2 54376 13552 54376 13552 0 net7
rlabel metal2 2240 56616 2240 56616 0 net70
rlabel metal2 2072 56840 2072 56840 0 net71
rlabel metal2 2744 57456 2744 57456 0 net72
rlabel metal2 3304 58072 3304 58072 0 net73
rlabel metal2 2296 59136 2296 59136 0 net74
rlabel metal2 3080 58856 3080 58856 0 net75
rlabel metal2 2184 60424 2184 60424 0 net76
rlabel metal2 2296 60704 2296 60704 0 net77
rlabel metal2 2072 61544 2072 61544 0 net78
rlabel metal2 2296 49224 2296 49224 0 net79
rlabel metal2 55048 14448 55048 14448 0 net8
rlabel metal2 2296 62216 2296 62216 0 net80
rlabel metal2 2184 63560 2184 63560 0 net81
rlabel metal2 2408 63336 2408 63336 0 net82
rlabel metal2 3192 63448 3192 63448 0 net83
rlabel metal2 2072 64288 2072 64288 0 net84
rlabel metal2 2296 65352 2296 65352 0 net85
rlabel metal2 2072 66304 2072 66304 0 net86
rlabel metal2 2296 67592 2296 67592 0 net87
rlabel metal2 2184 67368 2184 67368 0 net88
rlabel metal2 2296 68488 2296 68488 0 net89
rlabel metal2 54824 15008 54824 15008 0 net9
rlabel metal2 3080 49840 3080 49840 0 net90
rlabel metal2 67760 67928 67760 67928 0 net91
rlabel metal2 3192 68824 3192 68824 0 net92
rlabel metal2 2968 50568 2968 50568 0 net93
rlabel metal2 49224 51296 49224 51296 0 net94
rlabel metal2 48776 52640 48776 52640 0 net95
rlabel metal2 46984 52920 46984 52920 0 net96
rlabel metal2 2296 53984 2296 53984 0 net97
rlabel metal2 2744 52920 2744 52920 0 net98
rlabel metal3 51912 54600 51912 54600 0 net99
<< properties >>
string FIXED_BBOX 0 0 80000 80000
<< end >>
