// This is the unpowered netlist.
module wb_memory (csb_mem0,
    csb_mem1,
    io_wbs_ack,
    io_wbs_clk,
    io_wbs_cyc,
    io_wbs_rst,
    io_wbs_stb,
    io_wbs_we,
    web_mem0,
    web_mem1,
    addr_mem0,
    addr_mem1,
    din_mem0,
    din_mem1,
    dout_mem0,
    dout_mem1,
    io_wbs_adr,
    io_wbs_datrd,
    io_wbs_datwr,
    io_wbs_sel,
    wmask_mem0,
    wmask_mem1);
 output csb_mem0;
 output csb_mem1;
 output io_wbs_ack;
 input io_wbs_clk;
 input io_wbs_cyc;
 input io_wbs_rst;
 input io_wbs_stb;
 input io_wbs_we;
 output web_mem0;
 output web_mem1;
 output [8:0] addr_mem0;
 output [8:0] addr_mem1;
 output [31:0] din_mem0;
 output [31:0] din_mem1;
 input [31:0] dout_mem0;
 input [31:0] dout_mem1;
 input [31:0] io_wbs_adr;
 output [31:0] io_wbs_datrd;
 input [31:0] io_wbs_datwr;
 input [3:0] io_wbs_sel;
 output [3:0] wmask_mem0;
 output [3:0] wmask_mem1;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire net241;
 wire clknet_0_io_wbs_clk;
 wire operation;
 wire web_mem;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire clknet_2_0__leaf_io_wbs_clk;
 wire clknet_2_1__leaf_io_wbs_clk;
 wire clknet_2_2__leaf_io_wbs_clk;
 wire clknet_2_3__leaf_io_wbs_clk;

 gf180mcu_fd_sc_mcu7t5v0__buf_1 _168_ (.I(net66),
    .Z(_069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _169_ (.I0(net25),
    .I1(net57),
    .S(_069_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _170_ (.I(operation),
    .Z(_071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _171_ (.I(_071_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _172_ (.I0(net222),
    .I1(_070_),
    .S(_072_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _173_ (.I(_073_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _174_ (.I0(net24),
    .I1(net56),
    .S(_069_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _175_ (.I0(net221),
    .I1(_074_),
    .S(_072_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _176_ (.I(_075_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _177_ (.I(net66),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _178_ (.I(_076_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _179_ (.I0(net22),
    .I1(net54),
    .S(_077_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _180_ (.I0(net219),
    .I1(_078_),
    .S(_072_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _181_ (.I(_079_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _182_ (.I0(net21),
    .I1(net53),
    .S(_077_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _183_ (.I0(net218),
    .I1(_080_),
    .S(_072_),
    .Z(_081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _184_ (.I(_081_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _185_ (.I0(net20),
    .I1(net52),
    .S(_077_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _186_ (.I(_071_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _187_ (.I0(net217),
    .I1(_082_),
    .S(_083_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _188_ (.I(_084_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _189_ (.I0(net19),
    .I1(net51),
    .S(_077_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _190_ (.I0(net216),
    .I1(_085_),
    .S(_083_),
    .Z(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _191_ (.I(_086_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _192_ (.I(_076_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _193_ (.I0(net18),
    .I1(net50),
    .S(_087_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _194_ (.I0(net215),
    .I1(_088_),
    .S(_083_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _195_ (.I(_089_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _196_ (.I0(net17),
    .I1(net49),
    .S(_087_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _197_ (.I0(net214),
    .I1(_090_),
    .S(_083_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _198_ (.I(_091_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _199_ (.I0(net16),
    .I1(net48),
    .S(_087_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _200_ (.I(_071_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _201_ (.I0(net213),
    .I1(_092_),
    .S(_093_),
    .Z(_094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _202_ (.I(_094_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _203_ (.I0(net15),
    .I1(net47),
    .S(_087_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _204_ (.I0(net212),
    .I1(_095_),
    .S(_093_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _205_ (.I(_096_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _206_ (.I(net66),
    .Z(_097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _207_ (.I(_097_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _208_ (.I0(net14),
    .I1(net46),
    .S(_098_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _209_ (.I0(net211),
    .I1(_099_),
    .S(_093_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _210_ (.I(_100_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _211_ (.I0(net13),
    .I1(net45),
    .S(_098_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _212_ (.I0(net210),
    .I1(_101_),
    .S(_093_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _213_ (.I(_102_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _214_ (.I0(net11),
    .I1(net43),
    .S(_098_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _215_ (.I(operation),
    .Z(_104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _216_ (.I(_104_),
    .Z(_105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _217_ (.I0(net208),
    .I1(_103_),
    .S(_105_),
    .Z(_106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _218_ (.I(_106_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _219_ (.I0(net10),
    .I1(net42),
    .S(_098_),
    .Z(_107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _220_ (.I0(net207),
    .I1(_107_),
    .S(_105_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _221_ (.I(_108_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _222_ (.I(_097_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _223_ (.I0(net9),
    .I1(net41),
    .S(_109_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _224_ (.I0(net206),
    .I1(_110_),
    .S(_105_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _225_ (.I(_111_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _226_ (.I0(net8),
    .I1(net40),
    .S(_109_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _227_ (.I0(net205),
    .I1(_112_),
    .S(_105_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _228_ (.I(_113_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _229_ (.I0(net7),
    .I1(net39),
    .S(_109_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _230_ (.I(_104_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _231_ (.I0(net204),
    .I1(_114_),
    .S(_115_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _232_ (.I(_116_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _233_ (.I0(net6),
    .I1(net38),
    .S(_109_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _234_ (.I0(net203),
    .I1(_117_),
    .S(_115_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _235_ (.I(_118_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _236_ (.I(_097_),
    .Z(_119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _237_ (.I0(net5),
    .I1(net37),
    .S(_119_),
    .Z(_120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _238_ (.I0(net202),
    .I1(_120_),
    .S(_115_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _239_ (.I(_121_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _240_ (.I0(net4),
    .I1(net36),
    .S(_119_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _241_ (.I0(net201),
    .I1(_122_),
    .S(_115_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _242_ (.I(_123_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _243_ (.I0(net3),
    .I1(net35),
    .S(_119_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _244_ (.I(_104_),
    .Z(_125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _245_ (.I0(net200),
    .I1(_124_),
    .S(_125_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _246_ (.I(_126_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _247_ (.I0(net2),
    .I1(net34),
    .S(_119_),
    .Z(_127_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _248_ (.I0(net199),
    .I1(_127_),
    .S(_125_),
    .Z(_128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _249_ (.I(_128_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _250_ (.I(_097_),
    .Z(_129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _251_ (.I0(net32),
    .I1(net64),
    .S(_129_),
    .Z(_130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _252_ (.I0(net229),
    .I1(_130_),
    .S(_125_),
    .Z(_131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _253_ (.I(_131_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _254_ (.I0(net31),
    .I1(net63),
    .S(_129_),
    .Z(_132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _255_ (.I0(net228),
    .I1(_132_),
    .S(_125_),
    .Z(_133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _256_ (.I(_133_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _257_ (.I0(net30),
    .I1(net62),
    .S(_129_),
    .Z(_134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _258_ (.I(_104_),
    .Z(_135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _259_ (.I0(net227),
    .I1(_134_),
    .S(_135_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _260_ (.I(_136_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _261_ (.I0(net29),
    .I1(net61),
    .S(_129_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _262_ (.I0(net226),
    .I1(_137_),
    .S(_135_),
    .Z(_138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _263_ (.I(_138_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _264_ (.I(net66),
    .Z(_139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _265_ (.I0(net28),
    .I1(net60),
    .S(_139_),
    .Z(_140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _266_ (.I0(net225),
    .I1(_140_),
    .S(_135_),
    .Z(_141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _267_ (.I(_141_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _268_ (.I0(net27),
    .I1(net59),
    .S(_139_),
    .Z(_142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _269_ (.I0(net224),
    .I1(_142_),
    .S(_135_),
    .Z(_143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _270_ (.I(_143_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _271_ (.I0(net26),
    .I1(net58),
    .S(_139_),
    .Z(_144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _272_ (.I(operation),
    .Z(_145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _273_ (.I0(net223),
    .I1(_144_),
    .S(_145_),
    .Z(_146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _274_ (.I(_146_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _275_ (.I0(net23),
    .I1(net55),
    .S(_139_),
    .Z(_147_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _276_ (.I0(net220),
    .I1(_147_),
    .S(_145_),
    .Z(_148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _277_ (.I(_148_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _278_ (.I0(net12),
    .I1(net44),
    .S(_076_),
    .Z(_149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _279_ (.I0(net209),
    .I1(_149_),
    .S(_145_),
    .Z(_150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _280_ (.I(_150_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _281_ (.I0(net1),
    .I1(net33),
    .S(_076_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _282_ (.I0(net198),
    .I1(_151_),
    .S(_145_),
    .Z(_152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _283_ (.I(_152_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _284_ (.A1(_071_),
    .A2(net197),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _285_ (.A1(net113),
    .A2(net75),
    .A3(_153_),
    .Z(_154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _286_ (.I(_154_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _287_ (.A1(net113),
    .A2(net75),
    .A3(net114),
    .A4(_153_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _288_ (.I(web_mem),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _289_ (.A1(_155_),
    .A2(_069_),
    .ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _290_ (.A1(web_mem),
    .A2(_069_),
    .Z(_156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _291_ (.I(_156_),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _292_ (.I(net108),
    .Z(_157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _293_ (.I(_157_),
    .Z(_158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _294_ (.I(_158_),
    .Z(_159_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _295_ (.I(_159_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _296_ (.I(_159_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _297_ (.I(_159_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _298_ (.I(_159_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _299_ (.I(net108),
    .Z(_160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _300_ (.I(_160_),
    .Z(_161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _301_ (.I(_161_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _302_ (.I(_161_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _303_ (.I(_161_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _304_ (.I(_161_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _305_ (.I(_160_),
    .Z(_162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _306_ (.I(_162_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _307_ (.I(_162_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _308_ (.I(_162_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _309_ (.I(_162_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _310_ (.I(_160_),
    .Z(_163_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _311_ (.I(_163_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _312_ (.I(_163_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _313_ (.I(_163_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _314_ (.I(_163_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _315_ (.I(_160_),
    .Z(_164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _316_ (.I(_164_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _317_ (.I(_164_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _318_ (.I(_164_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _319_ (.I(_164_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _320_ (.I(_157_),
    .Z(_165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _321_ (.I(_165_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _322_ (.I(_165_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _323_ (.I(_165_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _324_ (.I(_165_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _325_ (.I(_157_),
    .Z(_166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _326_ (.I(_166_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _327_ (.I(_166_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _328_ (.I(_166_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _329_ (.I(_166_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _330_ (.I(_157_),
    .Z(_167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _331_ (.I(_167_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _332_ (.I(_167_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _333_ (.I(_167_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _334_ (.I(_167_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _335_ (.I(_158_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _336_ (.I(_158_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _337_ (.I(_158_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _338_ (.D(_037_),
    .RN(_002_),
    .CLK(clknet_2_1__leaf_io_wbs_clk),
    .Q(net198));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _339_ (.D(_038_),
    .RN(_003_),
    .CLK(clknet_2_0__leaf_io_wbs_clk),
    .Q(net209));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _340_ (.D(_039_),
    .RN(_004_),
    .CLK(clknet_2_0__leaf_io_wbs_clk),
    .Q(net220));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _341_ (.D(_040_),
    .RN(_005_),
    .CLK(clknet_2_1__leaf_io_wbs_clk),
    .Q(net223));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _342_ (.D(_041_),
    .RN(_006_),
    .CLK(clknet_2_1__leaf_io_wbs_clk),
    .Q(net224));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _343_ (.D(_042_),
    .RN(_007_),
    .CLK(clknet_2_0__leaf_io_wbs_clk),
    .Q(net225));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _344_ (.D(_043_),
    .RN(_008_),
    .CLK(clknet_2_1__leaf_io_wbs_clk),
    .Q(net226));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _345_ (.D(_044_),
    .RN(_009_),
    .CLK(clknet_2_1__leaf_io_wbs_clk),
    .Q(net227));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _346_ (.D(_045_),
    .RN(_010_),
    .CLK(clknet_2_1__leaf_io_wbs_clk),
    .Q(net228));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _347_ (.D(_046_),
    .RN(_011_),
    .CLK(clknet_2_3__leaf_io_wbs_clk),
    .Q(net229));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _348_ (.D(_047_),
    .RN(_012_),
    .CLK(clknet_2_1__leaf_io_wbs_clk),
    .Q(net199));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _349_ (.D(_048_),
    .RN(_013_),
    .CLK(clknet_2_0__leaf_io_wbs_clk),
    .Q(net200));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _350_ (.D(_049_),
    .RN(_014_),
    .CLK(clknet_2_2__leaf_io_wbs_clk),
    .Q(net201));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _351_ (.D(_050_),
    .RN(_015_),
    .CLK(clknet_2_3__leaf_io_wbs_clk),
    .Q(net202));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _352_ (.D(_051_),
    .RN(_016_),
    .CLK(clknet_2_2__leaf_io_wbs_clk),
    .Q(net203));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _353_ (.D(_052_),
    .RN(_017_),
    .CLK(clknet_2_3__leaf_io_wbs_clk),
    .Q(net204));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _354_ (.D(_053_),
    .RN(_018_),
    .CLK(clknet_2_3__leaf_io_wbs_clk),
    .Q(net205));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _355_ (.D(_054_),
    .RN(_019_),
    .CLK(clknet_2_2__leaf_io_wbs_clk),
    .Q(net206));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _356_ (.D(_055_),
    .RN(_020_),
    .CLK(clknet_2_2__leaf_io_wbs_clk),
    .Q(net207));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _357_ (.D(_056_),
    .RN(_021_),
    .CLK(clknet_2_3__leaf_io_wbs_clk),
    .Q(net208));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _358_ (.D(_057_),
    .RN(_022_),
    .CLK(clknet_2_2__leaf_io_wbs_clk),
    .Q(net210));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _359_ (.D(_058_),
    .RN(_023_),
    .CLK(clknet_2_3__leaf_io_wbs_clk),
    .Q(net211));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _360_ (.D(_059_),
    .RN(_024_),
    .CLK(clknet_2_3__leaf_io_wbs_clk),
    .Q(net212));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _361_ (.D(_060_),
    .RN(_025_),
    .CLK(clknet_2_2__leaf_io_wbs_clk),
    .Q(net213));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _362_ (.D(_061_),
    .RN(_026_),
    .CLK(clknet_2_3__leaf_io_wbs_clk),
    .Q(net214));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _363_ (.D(_062_),
    .RN(_027_),
    .CLK(clknet_2_2__leaf_io_wbs_clk),
    .Q(net215));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _364_ (.D(_063_),
    .RN(_028_),
    .CLK(clknet_2_2__leaf_io_wbs_clk),
    .Q(net216));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _365_ (.D(_064_),
    .RN(_029_),
    .CLK(clknet_2_2__leaf_io_wbs_clk),
    .Q(net217));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _366_ (.D(_065_),
    .RN(_030_),
    .CLK(clknet_2_2__leaf_io_wbs_clk),
    .Q(net218));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _367_ (.D(_066_),
    .RN(_031_),
    .CLK(clknet_2_3__leaf_io_wbs_clk),
    .Q(net219));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _368_ (.D(_067_),
    .RN(_032_),
    .CLK(clknet_2_3__leaf_io_wbs_clk),
    .Q(net221));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _369_ (.D(_068_),
    .RN(_033_),
    .CLK(clknet_2_3__leaf_io_wbs_clk),
    .Q(net222));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _370_ (.D(operation),
    .RN(_034_),
    .CLK(clknet_2_0__leaf_io_wbs_clk),
    .Q(net197));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _371_ (.D(_001_),
    .SETN(_035_),
    .CLK(clknet_2_0__leaf_io_wbs_clk),
    .Q(web_mem));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _372_ (.D(_000_),
    .RN(_036_),
    .CLK(clknet_2_0__leaf_io_wbs_clk),
    .Q(operation));
 gf180mcu_fd_sc_mcu7t5v0__tiel wb_memory_241 (.ZN(net241));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_io_wbs_clk (.I(io_wbs_clk),
    .Z(clknet_0_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _375_ (.I(net67),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _376_ (.I(net68),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _377_ (.I(net69),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _378_ (.I(net70),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _379_ (.I(net71),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _380_ (.I(net72),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _381_ (.I(net73),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _382_ (.I(net74),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _383_ (.I(net65),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _384_ (.I(net67),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _385_ (.I(net68),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _386_ (.I(net69),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _387_ (.I(net70),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _388_ (.I(net71),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _389_ (.I(net72),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _390_ (.I(net73),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _391_ (.I(net74),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _392_ (.I(net65),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _393_ (.I(net76),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _394_ (.I(net87),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _395_ (.I(net98),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _396_ (.I(net101),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _397_ (.I(net102),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _398_ (.I(net103),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _399_ (.I(net104),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _400_ (.I(net105),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _401_ (.I(net106),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _402_ (.I(net107),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _403_ (.I(net77),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _404_ (.I(net78),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _405_ (.I(net79),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _406_ (.I(net80),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _407_ (.I(net81),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _408_ (.I(net82),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _409_ (.I(net83),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _410_ (.I(net84),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _411_ (.I(net85),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _412_ (.I(net86),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _413_ (.I(net88),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _414_ (.I(net89),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _415_ (.I(net90),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _416_ (.I(net91),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _417_ (.I(net92),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _418_ (.I(net93),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _419_ (.I(net94),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _420_ (.I(net95),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _421_ (.I(net96),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _422_ (.I(net97),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _423_ (.I(net99),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _424_ (.I(net100),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _425_ (.I(net76),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _426_ (.I(net87),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _427_ (.I(net98),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _428_ (.I(net101),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _429_ (.I(net102),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _430_ (.I(net103),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _431_ (.I(net104),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _432_ (.I(net105),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _433_ (.I(net106),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _434_ (.I(net107),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _435_ (.I(net77),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _436_ (.I(net78),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _437_ (.I(net79),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _438_ (.I(net80),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _439_ (.I(net81),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _440_ (.I(net82),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _441_ (.I(net83),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _442_ (.I(net84),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _443_ (.I(net85),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _444_ (.I(net86),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _445_ (.I(net88),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _446_ (.I(net89),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _447_ (.I(net90),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _448_ (.I(net91),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _449_ (.I(net92),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _450_ (.I(net93),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _451_ (.I(net94),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _452_ (.I(net95),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _453_ (.I(net96),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _454_ (.I(net97),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _455_ (.I(net99),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _456_ (.I(net100),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _457_ (.I(net109),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _458_ (.I(net110),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _459_ (.I(net111),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _460_ (.I(net112),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _461_ (.I(net109),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _462_ (.I(net110),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _463_ (.I(net111),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _464_ (.I(net112),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(dout_mem0[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(dout_mem0[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(dout_mem0[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(dout_mem0[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(dout_mem0[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(dout_mem0[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(dout_mem0[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(dout_mem0[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(dout_mem0[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(dout_mem0[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(dout_mem0[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(dout_mem0[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(dout_mem0[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(dout_mem0[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(dout_mem0[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(dout_mem0[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(dout_mem0[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(dout_mem0[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(dout_mem0[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(dout_mem0[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(dout_mem0[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(dout_mem0[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(dout_mem0[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(dout_mem0[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(dout_mem0[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(dout_mem0[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(dout_mem0[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(dout_mem0[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(dout_mem0[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(dout_mem0[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(dout_mem0[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(dout_mem0[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(dout_mem1[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(dout_mem1[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(dout_mem1[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(dout_mem1[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(dout_mem1[13]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(dout_mem1[14]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(dout_mem1[15]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(dout_mem1[16]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(dout_mem1[17]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(dout_mem1[18]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(dout_mem1[19]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(dout_mem1[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(dout_mem1[20]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input46 (.I(dout_mem1[21]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input47 (.I(dout_mem1[22]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input48 (.I(dout_mem1[23]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input49 (.I(dout_mem1[24]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input50 (.I(dout_mem1[25]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(dout_mem1[26]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(dout_mem1[27]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(dout_mem1[28]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(dout_mem1[29]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(dout_mem1[2]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(dout_mem1[30]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(dout_mem1[31]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(dout_mem1[3]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input59 (.I(dout_mem1[4]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input60 (.I(dout_mem1[5]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input61 (.I(dout_mem1[6]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input62 (.I(dout_mem1[7]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input63 (.I(dout_mem1[8]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input64 (.I(dout_mem1[9]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input65 (.I(io_wbs_adr[10]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input66 (.I(io_wbs_adr[11]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input67 (.I(io_wbs_adr[2]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(io_wbs_adr[3]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input69 (.I(io_wbs_adr[4]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input70 (.I(io_wbs_adr[5]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(io_wbs_adr[6]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input72 (.I(io_wbs_adr[7]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input73 (.I(io_wbs_adr[8]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input74 (.I(io_wbs_adr[9]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input75 (.I(io_wbs_cyc),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input76 (.I(io_wbs_datwr[0]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input77 (.I(io_wbs_datwr[10]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(io_wbs_datwr[11]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input79 (.I(io_wbs_datwr[12]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(io_wbs_datwr[13]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(io_wbs_datwr[14]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input82 (.I(io_wbs_datwr[15]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input83 (.I(io_wbs_datwr[16]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input84 (.I(io_wbs_datwr[17]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input85 (.I(io_wbs_datwr[18]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input86 (.I(io_wbs_datwr[19]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input87 (.I(io_wbs_datwr[1]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input88 (.I(io_wbs_datwr[20]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input89 (.I(io_wbs_datwr[21]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input90 (.I(io_wbs_datwr[22]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input91 (.I(io_wbs_datwr[23]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input92 (.I(io_wbs_datwr[24]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input93 (.I(io_wbs_datwr[25]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input94 (.I(io_wbs_datwr[26]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input95 (.I(io_wbs_datwr[27]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input96 (.I(io_wbs_datwr[28]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input97 (.I(io_wbs_datwr[29]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input98 (.I(io_wbs_datwr[2]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input99 (.I(io_wbs_datwr[30]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input100 (.I(io_wbs_datwr[31]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input101 (.I(io_wbs_datwr[3]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input102 (.I(io_wbs_datwr[4]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input103 (.I(io_wbs_datwr[5]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input104 (.I(io_wbs_datwr[6]),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input105 (.I(io_wbs_datwr[7]),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input106 (.I(io_wbs_datwr[8]),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input107 (.I(io_wbs_datwr[9]),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input108 (.I(io_wbs_rst),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input109 (.I(io_wbs_sel[0]),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input110 (.I(io_wbs_sel[1]),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input111 (.I(io_wbs_sel[2]),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input112 (.I(io_wbs_sel[3]),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input113 (.I(io_wbs_stb),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input114 (.I(io_wbs_we),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output115 (.I(net115),
    .Z(addr_mem0[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output116 (.I(net116),
    .Z(addr_mem0[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output117 (.I(net117),
    .Z(addr_mem0[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output118 (.I(net118),
    .Z(addr_mem0[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output119 (.I(net119),
    .Z(addr_mem0[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output120 (.I(net120),
    .Z(addr_mem0[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output121 (.I(net121),
    .Z(addr_mem0[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output122 (.I(net122),
    .Z(addr_mem0[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output123 (.I(net123),
    .Z(addr_mem0[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output124 (.I(net124),
    .Z(addr_mem1[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output125 (.I(net125),
    .Z(addr_mem1[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output126 (.I(net126),
    .Z(addr_mem1[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output127 (.I(net127),
    .Z(addr_mem1[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output128 (.I(net128),
    .Z(addr_mem1[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output129 (.I(net129),
    .Z(addr_mem1[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output130 (.I(net130),
    .Z(addr_mem1[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output131 (.I(net131),
    .Z(addr_mem1[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output132 (.I(net132),
    .Z(addr_mem1[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output133 (.I(net133),
    .Z(din_mem0[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output134 (.I(net134),
    .Z(din_mem0[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output135 (.I(net135),
    .Z(din_mem0[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output136 (.I(net136),
    .Z(din_mem0[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output137 (.I(net137),
    .Z(din_mem0[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output138 (.I(net138),
    .Z(din_mem0[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output139 (.I(net139),
    .Z(din_mem0[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output140 (.I(net140),
    .Z(din_mem0[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output141 (.I(net141),
    .Z(din_mem0[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output142 (.I(net142),
    .Z(din_mem0[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output143 (.I(net143),
    .Z(din_mem0[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output144 (.I(net144),
    .Z(din_mem0[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output145 (.I(net145),
    .Z(din_mem0[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output146 (.I(net146),
    .Z(din_mem0[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output147 (.I(net147),
    .Z(din_mem0[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output148 (.I(net148),
    .Z(din_mem0[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output149 (.I(net149),
    .Z(din_mem0[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output150 (.I(net150),
    .Z(din_mem0[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output151 (.I(net151),
    .Z(din_mem0[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output152 (.I(net152),
    .Z(din_mem0[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output153 (.I(net153),
    .Z(din_mem0[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output154 (.I(net154),
    .Z(din_mem0[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output155 (.I(net155),
    .Z(din_mem0[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output156 (.I(net156),
    .Z(din_mem0[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output157 (.I(net157),
    .Z(din_mem0[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output158 (.I(net158),
    .Z(din_mem0[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output159 (.I(net159),
    .Z(din_mem0[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output160 (.I(net160),
    .Z(din_mem0[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output161 (.I(net161),
    .Z(din_mem0[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output162 (.I(net162),
    .Z(din_mem0[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output163 (.I(net163),
    .Z(din_mem0[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output164 (.I(net164),
    .Z(din_mem0[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output165 (.I(net165),
    .Z(din_mem1[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output166 (.I(net166),
    .Z(din_mem1[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output167 (.I(net167),
    .Z(din_mem1[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output168 (.I(net168),
    .Z(din_mem1[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output169 (.I(net169),
    .Z(din_mem1[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output170 (.I(net170),
    .Z(din_mem1[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output171 (.I(net171),
    .Z(din_mem1[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output172 (.I(net172),
    .Z(din_mem1[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output173 (.I(net173),
    .Z(din_mem1[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output174 (.I(net174),
    .Z(din_mem1[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output175 (.I(net175),
    .Z(din_mem1[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output176 (.I(net176),
    .Z(din_mem1[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output177 (.I(net177),
    .Z(din_mem1[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output178 (.I(net178),
    .Z(din_mem1[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output179 (.I(net179),
    .Z(din_mem1[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output180 (.I(net180),
    .Z(din_mem1[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output181 (.I(net181),
    .Z(din_mem1[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output182 (.I(net182),
    .Z(din_mem1[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output183 (.I(net183),
    .Z(din_mem1[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output184 (.I(net184),
    .Z(din_mem1[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output185 (.I(net185),
    .Z(din_mem1[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output186 (.I(net186),
    .Z(din_mem1[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output187 (.I(net187),
    .Z(din_mem1[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output188 (.I(net188),
    .Z(din_mem1[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output189 (.I(net189),
    .Z(din_mem1[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output190 (.I(net190),
    .Z(din_mem1[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output191 (.I(net191),
    .Z(din_mem1[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output192 (.I(net192),
    .Z(din_mem1[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output193 (.I(net193),
    .Z(din_mem1[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output194 (.I(net194),
    .Z(din_mem1[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output195 (.I(net195),
    .Z(din_mem1[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output196 (.I(net196),
    .Z(din_mem1[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output197 (.I(net197),
    .Z(io_wbs_ack));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output198 (.I(net198),
    .Z(io_wbs_datrd[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output199 (.I(net199),
    .Z(io_wbs_datrd[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output200 (.I(net200),
    .Z(io_wbs_datrd[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output201 (.I(net201),
    .Z(io_wbs_datrd[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output202 (.I(net202),
    .Z(io_wbs_datrd[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output203 (.I(net203),
    .Z(io_wbs_datrd[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output204 (.I(net204),
    .Z(io_wbs_datrd[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output205 (.I(net205),
    .Z(io_wbs_datrd[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output206 (.I(net206),
    .Z(io_wbs_datrd[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output207 (.I(net207),
    .Z(io_wbs_datrd[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output208 (.I(net208),
    .Z(io_wbs_datrd[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output209 (.I(net209),
    .Z(io_wbs_datrd[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output210 (.I(net210),
    .Z(io_wbs_datrd[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output211 (.I(net211),
    .Z(io_wbs_datrd[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output212 (.I(net212),
    .Z(io_wbs_datrd[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output213 (.I(net213),
    .Z(io_wbs_datrd[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output214 (.I(net214),
    .Z(io_wbs_datrd[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output215 (.I(net215),
    .Z(io_wbs_datrd[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output216 (.I(net216),
    .Z(io_wbs_datrd[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output217 (.I(net217),
    .Z(io_wbs_datrd[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output218 (.I(net218),
    .Z(io_wbs_datrd[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output219 (.I(net219),
    .Z(io_wbs_datrd[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output220 (.I(net220),
    .Z(io_wbs_datrd[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output221 (.I(net221),
    .Z(io_wbs_datrd[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output222 (.I(net222),
    .Z(io_wbs_datrd[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output223 (.I(net223),
    .Z(io_wbs_datrd[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output224 (.I(net224),
    .Z(io_wbs_datrd[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output225 (.I(net225),
    .Z(io_wbs_datrd[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output226 (.I(net226),
    .Z(io_wbs_datrd[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output227 (.I(net227),
    .Z(io_wbs_datrd[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output228 (.I(net228),
    .Z(io_wbs_datrd[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output229 (.I(net229),
    .Z(io_wbs_datrd[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output230 (.I(net230),
    .Z(web_mem0));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output231 (.I(net231),
    .Z(web_mem1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output232 (.I(net232),
    .Z(wmask_mem0[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output233 (.I(net233),
    .Z(wmask_mem0[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output234 (.I(net234),
    .Z(wmask_mem0[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output235 (.I(net235),
    .Z(wmask_mem0[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output236 (.I(net236),
    .Z(wmask_mem1[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output237 (.I(net237),
    .Z(wmask_mem1[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output238 (.I(net238),
    .Z(wmask_mem1[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output239 (.I(net239),
    .Z(wmask_mem1[3]));
 gf180mcu_fd_sc_mcu7t5v0__tiel wb_memory_240 (.ZN(net240));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_io_wbs_clk (.I(clknet_0_io_wbs_clk),
    .Z(clknet_2_0__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_io_wbs_clk (.I(clknet_0_io_wbs_clk),
    .Z(clknet_2_1__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_io_wbs_clk (.I(clknet_0_io_wbs_clk),
    .Z(clknet_2_2__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_io_wbs_clk (.I(clknet_0_io_wbs_clk),
    .Z(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__D (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__D (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__D (.I(_066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__S (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__S (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__I1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__I (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__186__I (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__171__I (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__S (.I(_072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__S (.I(_072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__S (.I(_072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__S (.I(_072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__I1 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__S (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__S (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__192__I (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__I (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__189__S (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__S (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__S (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__S (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__I1 (.I(_078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__I1 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__187__I1 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__S (.I(_083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__194__S (.I(_083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__190__S (.I(_083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__187__S (.I(_083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__190__I1 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__194__I1 (.I(_088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__I1 (.I(_090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__201__I1 (.I(_092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__S (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__209__S (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__S (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__201__S (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__I1 (.I(_095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__250__I (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__236__I (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__222__I (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__207__I (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__S (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__S (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__211__S (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__208__S (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__209__I1 (.I(_099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__I1 (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__217__I1 (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__I (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__244__I (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__I (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__216__I (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__S (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__S (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__S (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__217__S (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__I1 (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__I1 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__I1 (.I(_112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__I1 (.I(_114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__S (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__S (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__S (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__S (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__I1 (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__S (.I(_119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__S (.I(_119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__240__S (.I(_119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__S (.I(_119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__I1 (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__I1 (.I(_122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__245__I1 (.I(_124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__248__I1 (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__S (.I(_129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__S (.I(_129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__S (.I(_129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__S (.I(_129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__I1 (.I(_130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__I1 (.I(_132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__I1 (.I(_134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__S (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__S (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__S (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__S (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__I1 (.I(_137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__S (.I(_139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__S (.I(_139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__S (.I(_139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__S (.I(_139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__I1 (.I(_140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__I1 (.I(_142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__273__I1 (.I(_144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__S (.I(_145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__S (.I(_145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__S (.I(_145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__273__S (.I(_145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__I1 (.I(_147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__I1 (.I(_149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__I1 (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A4 (.I(_153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__285__A3 (.I(_153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__330__I (.I(_157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__I (.I(_157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__I (.I(_157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__I (.I(_157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__I (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__I (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__I (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__I (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__I (.I(_159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__I (.I(_159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__I (.I(_159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__I (.I(_159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__I (.I(_160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__I (.I(_160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__I (.I(_160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__I (.I(_160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__I (.I(_163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__I (.I(_163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__I (.I(_163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__I (.I(_163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__I (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__318__I (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__I (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__I (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__324__I (.I(_165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__323__I (.I(_165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__I (.I(_165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__321__I (.I(_165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_io_wbs_clk_I (.I(clknet_0_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_io_wbs_clk_I (.I(clknet_0_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_io_wbs_clk_I (.I(clknet_0_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_io_wbs_clk_I (.I(clknet_0_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(dout_mem0[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(dout_mem0[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(dout_mem0[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(dout_mem0[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(dout_mem0[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(dout_mem0[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(dout_mem0[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(dout_mem0[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(dout_mem0[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(dout_mem0[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(dout_mem0[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(dout_mem0[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(dout_mem0[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(dout_mem0[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(dout_mem0[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(dout_mem0[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(dout_mem0[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(dout_mem0[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(dout_mem0[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(dout_mem0[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(dout_mem0[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(dout_mem0[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(dout_mem0[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(dout_mem0[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(dout_mem0[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(dout_mem0[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(dout_mem0[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(dout_mem0[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(dout_mem0[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(dout_mem0[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(dout_mem0[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(dout_mem0[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(dout_mem1[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(dout_mem1[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(dout_mem1[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(dout_mem1[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(dout_mem1[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(dout_mem1[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(dout_mem1[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(dout_mem1[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(dout_mem1[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(dout_mem1[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(dout_mem1[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(dout_mem1[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(dout_mem1[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(dout_mem1[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(dout_mem1[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(dout_mem1[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(dout_mem1[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(dout_mem1[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(dout_mem1[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(dout_mem1[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(dout_mem1[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(dout_mem1[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(dout_mem1[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(dout_mem1[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(dout_mem1[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(dout_mem1[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(dout_mem1[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(dout_mem1[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(dout_mem1[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(dout_mem1[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(dout_mem1[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(dout_mem1[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(io_wbs_adr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(io_wbs_adr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(io_wbs_adr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(io_wbs_adr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(io_wbs_adr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(io_wbs_adr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(io_wbs_adr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(io_wbs_adr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(io_wbs_adr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(io_wbs_adr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_io_wbs_clk_I (.I(io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(io_wbs_cyc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(io_wbs_datwr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(io_wbs_datwr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(io_wbs_datwr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(io_wbs_datwr[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(io_wbs_datwr[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(io_wbs_datwr[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(io_wbs_datwr[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(io_wbs_datwr[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(io_wbs_datwr[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(io_wbs_datwr[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(io_wbs_datwr[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(io_wbs_datwr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(io_wbs_datwr[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(io_wbs_datwr[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(io_wbs_datwr[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(io_wbs_datwr[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(io_wbs_datwr[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(io_wbs_datwr[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(io_wbs_datwr[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(io_wbs_datwr[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(io_wbs_datwr[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(io_wbs_datwr[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input98_I (.I(io_wbs_datwr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input99_I (.I(io_wbs_datwr[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input100_I (.I(io_wbs_datwr[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input101_I (.I(io_wbs_datwr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input102_I (.I(io_wbs_datwr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input103_I (.I(io_wbs_datwr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input104_I (.I(io_wbs_datwr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input105_I (.I(io_wbs_datwr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input106_I (.I(io_wbs_datwr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input107_I (.I(io_wbs_datwr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input108_I (.I(io_wbs_rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input109_I (.I(io_wbs_sel[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input110_I (.I(io_wbs_sel[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input111_I (.I(io_wbs_sel[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input112_I (.I(io_wbs_sel[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input113_I (.I(io_wbs_stb));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input114_I (.I(io_wbs_we));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__D (.I(operation));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__I (.I(operation));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__215__I (.I(operation));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__I (.I(operation));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A1 (.I(web_mem));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__288__I (.I(web_mem));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__I0 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__I0 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__I0 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__240__I0 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__I0 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__I0 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__I0 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__I0 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__223__I0 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__I0 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__I0 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__211__I0 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__208__I0 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I0 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__199__I0 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__I0 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__193__I0 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__189__I0 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__I0 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__I0 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__I0 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__I0 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__I0 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__I0 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__I0 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__I0 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__I0 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__I0 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__I0 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__I1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__I1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__I1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__240__I1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__I1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__I1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__I1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__I1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__223__I1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__I1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__I1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__I1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__211__I1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__208__I1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__199__I1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__I1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__I1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__I1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__I1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__I1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__I1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__I1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__I1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__I1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__I1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__392__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__383__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__177__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__385__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__376__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__386__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__377__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__387__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__378__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__379__I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__389__I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__380__I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__390__I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__381__I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__382__I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__425__I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__393__I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__435__I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__436__I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__437__I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__406__I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__439__I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__440__I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__409__I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__442__I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__443__I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__411__I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__444__I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__426__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__394__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__445__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__415__I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__416__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__449__I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__417__I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__450__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__418__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__452__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__453__I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__454__I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__422__I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__427__I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__395__I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__456__I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__424__I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__428__I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__429__I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__397__I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__430__I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__398__I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__431__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__399__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__432__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__400__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__433__I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__434__I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__461__I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__462__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__459__I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output128_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output129_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output130_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output131_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output132_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output138_I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output145_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output149_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output152_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output153_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output154_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output157_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output180_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output191_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output193_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output194_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output195_I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output196_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output197_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__A2 (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output201_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__I0 (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output202_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__I0 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output203_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__I0 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output204_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__I0 (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output205_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__I0 (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output206_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__I0 (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output207_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__I0 (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output208_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__217__I0 (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output210_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__I0 (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output212_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__I0 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output214_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__I0 (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output215_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__194__I0 (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output216_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__190__I0 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output217_I (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__187__I0 (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output218_I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__I0 (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output219_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__I0 (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output221_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__I0 (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output222_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__I0 (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output224_I (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__I0 (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output226_I (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__I0 (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output227_I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__I0 (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output228_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__I0 (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output229_I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__I0 (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output230_I (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output236_I (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output237_I (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output239_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__339__CLK (.I(clknet_2_0__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__CLK (.I(clknet_2_0__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__CLK (.I(clknet_2_0__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__CLK (.I(clknet_2_0__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__CLK (.I(clknet_2_0__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__CLK (.I(clknet_2_0__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__372__CLK (.I(clknet_2_0__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__CLK (.I(clknet_2_1__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__341__CLK (.I(clknet_2_1__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__CLK (.I(clknet_2_1__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__CLK (.I(clknet_2_1__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__CLK (.I(clknet_2_1__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__CLK (.I(clknet_2_1__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__CLK (.I(clknet_2_1__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__CLK (.I(clknet_2_2__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__CLK (.I(clknet_2_2__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__CLK (.I(clknet_2_2__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__CLK (.I(clknet_2_2__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__CLK (.I(clknet_2_2__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__CLK (.I(clknet_2_2__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__CLK (.I(clknet_2_2__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__CLK (.I(clknet_2_2__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__CLK (.I(clknet_2_2__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__CLK (.I(clknet_2_2__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__CLK (.I(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__CLK (.I(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__CLK (.I(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__CLK (.I(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__CLK (.I(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__359__CLK (.I(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__CLK (.I(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__CLK (.I(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__CLK (.I(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__CLK (.I(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__CLK (.I(clknet_2_3__leaf_io_wbs_clk));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1297 ();
 assign csb_mem0 = net240;
 assign csb_mem1 = net241;
endmodule

