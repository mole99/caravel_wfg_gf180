magic
tech gf180mcuC
magscale 1 5
timestamp 1670255127
<< obsm1 >>
rect 672 1538 39312 38446
<< metal2 >>
rect 2632 0 2688 400
rect 2968 0 3024 400
rect 3304 0 3360 400
rect 3640 0 3696 400
rect 3976 0 4032 400
rect 4312 0 4368 400
rect 4648 0 4704 400
rect 4984 0 5040 400
rect 5320 0 5376 400
rect 5656 0 5712 400
rect 5992 0 6048 400
rect 6328 0 6384 400
rect 6664 0 6720 400
rect 7000 0 7056 400
rect 7336 0 7392 400
rect 7672 0 7728 400
rect 8008 0 8064 400
rect 8344 0 8400 400
rect 8680 0 8736 400
rect 9016 0 9072 400
rect 9352 0 9408 400
rect 9688 0 9744 400
rect 10024 0 10080 400
rect 10360 0 10416 400
rect 10696 0 10752 400
rect 11032 0 11088 400
rect 11368 0 11424 400
rect 11704 0 11760 400
rect 12040 0 12096 400
rect 12376 0 12432 400
rect 12712 0 12768 400
rect 13048 0 13104 400
rect 13384 0 13440 400
rect 13720 0 13776 400
rect 14056 0 14112 400
rect 14392 0 14448 400
rect 14728 0 14784 400
rect 15064 0 15120 400
rect 15400 0 15456 400
rect 15736 0 15792 400
rect 16072 0 16128 400
rect 16408 0 16464 400
rect 16744 0 16800 400
rect 17080 0 17136 400
rect 17416 0 17472 400
rect 17752 0 17808 400
rect 18088 0 18144 400
rect 18424 0 18480 400
rect 18760 0 18816 400
rect 19096 0 19152 400
rect 19432 0 19488 400
rect 19768 0 19824 400
rect 20104 0 20160 400
rect 20440 0 20496 400
rect 20776 0 20832 400
rect 21112 0 21168 400
rect 21448 0 21504 400
rect 21784 0 21840 400
rect 22120 0 22176 400
rect 22456 0 22512 400
rect 22792 0 22848 400
rect 23128 0 23184 400
rect 23464 0 23520 400
rect 23800 0 23856 400
rect 24136 0 24192 400
rect 24472 0 24528 400
rect 24808 0 24864 400
rect 25144 0 25200 400
rect 25480 0 25536 400
rect 25816 0 25872 400
rect 26152 0 26208 400
rect 26488 0 26544 400
rect 26824 0 26880 400
rect 27160 0 27216 400
rect 27496 0 27552 400
rect 27832 0 27888 400
rect 28168 0 28224 400
rect 28504 0 28560 400
rect 28840 0 28896 400
rect 29176 0 29232 400
rect 29512 0 29568 400
rect 29848 0 29904 400
rect 30184 0 30240 400
rect 30520 0 30576 400
rect 30856 0 30912 400
rect 31192 0 31248 400
rect 31528 0 31584 400
rect 31864 0 31920 400
rect 32200 0 32256 400
rect 32536 0 32592 400
rect 32872 0 32928 400
rect 33208 0 33264 400
rect 33544 0 33600 400
rect 33880 0 33936 400
rect 34216 0 34272 400
rect 34552 0 34608 400
rect 34888 0 34944 400
rect 35224 0 35280 400
rect 35560 0 35616 400
rect 35896 0 35952 400
rect 36232 0 36288 400
rect 36568 0 36624 400
rect 36904 0 36960 400
rect 37240 0 37296 400
<< obsm2 >>
rect 854 430 38962 38435
rect 854 400 2602 430
rect 2718 400 2938 430
rect 3054 400 3274 430
rect 3390 400 3610 430
rect 3726 400 3946 430
rect 4062 400 4282 430
rect 4398 400 4618 430
rect 4734 400 4954 430
rect 5070 400 5290 430
rect 5406 400 5626 430
rect 5742 400 5962 430
rect 6078 400 6298 430
rect 6414 400 6634 430
rect 6750 400 6970 430
rect 7086 400 7306 430
rect 7422 400 7642 430
rect 7758 400 7978 430
rect 8094 400 8314 430
rect 8430 400 8650 430
rect 8766 400 8986 430
rect 9102 400 9322 430
rect 9438 400 9658 430
rect 9774 400 9994 430
rect 10110 400 10330 430
rect 10446 400 10666 430
rect 10782 400 11002 430
rect 11118 400 11338 430
rect 11454 400 11674 430
rect 11790 400 12010 430
rect 12126 400 12346 430
rect 12462 400 12682 430
rect 12798 400 13018 430
rect 13134 400 13354 430
rect 13470 400 13690 430
rect 13806 400 14026 430
rect 14142 400 14362 430
rect 14478 400 14698 430
rect 14814 400 15034 430
rect 15150 400 15370 430
rect 15486 400 15706 430
rect 15822 400 16042 430
rect 16158 400 16378 430
rect 16494 400 16714 430
rect 16830 400 17050 430
rect 17166 400 17386 430
rect 17502 400 17722 430
rect 17838 400 18058 430
rect 18174 400 18394 430
rect 18510 400 18730 430
rect 18846 400 19066 430
rect 19182 400 19402 430
rect 19518 400 19738 430
rect 19854 400 20074 430
rect 20190 400 20410 430
rect 20526 400 20746 430
rect 20862 400 21082 430
rect 21198 400 21418 430
rect 21534 400 21754 430
rect 21870 400 22090 430
rect 22206 400 22426 430
rect 22542 400 22762 430
rect 22878 400 23098 430
rect 23214 400 23434 430
rect 23550 400 23770 430
rect 23886 400 24106 430
rect 24222 400 24442 430
rect 24558 400 24778 430
rect 24894 400 25114 430
rect 25230 400 25450 430
rect 25566 400 25786 430
rect 25902 400 26122 430
rect 26238 400 26458 430
rect 26574 400 26794 430
rect 26910 400 27130 430
rect 27246 400 27466 430
rect 27582 400 27802 430
rect 27918 400 28138 430
rect 28254 400 28474 430
rect 28590 400 28810 430
rect 28926 400 29146 430
rect 29262 400 29482 430
rect 29598 400 29818 430
rect 29934 400 30154 430
rect 30270 400 30490 430
rect 30606 400 30826 430
rect 30942 400 31162 430
rect 31278 400 31498 430
rect 31614 400 31834 430
rect 31950 400 32170 430
rect 32286 400 32506 430
rect 32622 400 32842 430
rect 32958 400 33178 430
rect 33294 400 33514 430
rect 33630 400 33850 430
rect 33966 400 34186 430
rect 34302 400 34522 430
rect 34638 400 34858 430
rect 34974 400 35194 430
rect 35310 400 35530 430
rect 35646 400 35866 430
rect 35982 400 36202 430
rect 36318 400 36538 430
rect 36654 400 36874 430
rect 36990 400 37210 430
rect 37326 400 38962 430
<< metal3 >>
rect 0 37240 400 37296
rect 39600 37240 40000 37296
rect 0 36904 400 36960
rect 39600 36904 40000 36960
rect 0 36568 400 36624
rect 39600 36568 40000 36624
rect 0 36232 400 36288
rect 39600 36232 40000 36288
rect 0 35896 400 35952
rect 39600 35896 40000 35952
rect 0 35560 400 35616
rect 39600 35560 40000 35616
rect 0 35224 400 35280
rect 39600 35224 40000 35280
rect 0 34888 400 34944
rect 39600 34888 40000 34944
rect 0 34552 400 34608
rect 39600 34552 40000 34608
rect 0 34216 400 34272
rect 39600 34216 40000 34272
rect 0 33880 400 33936
rect 39600 33880 40000 33936
rect 0 33544 400 33600
rect 39600 33544 40000 33600
rect 0 33208 400 33264
rect 39600 33208 40000 33264
rect 0 32872 400 32928
rect 39600 32872 40000 32928
rect 0 32536 400 32592
rect 39600 32536 40000 32592
rect 0 32200 400 32256
rect 39600 32200 40000 32256
rect 0 31864 400 31920
rect 39600 31864 40000 31920
rect 0 31528 400 31584
rect 39600 31528 40000 31584
rect 0 31192 400 31248
rect 39600 31192 40000 31248
rect 0 30856 400 30912
rect 39600 30856 40000 30912
rect 0 30520 400 30576
rect 39600 30520 40000 30576
rect 0 30184 400 30240
rect 39600 30184 40000 30240
rect 0 29848 400 29904
rect 39600 29848 40000 29904
rect 0 29512 400 29568
rect 39600 29512 40000 29568
rect 0 29176 400 29232
rect 39600 29176 40000 29232
rect 0 28840 400 28896
rect 39600 28840 40000 28896
rect 0 28504 400 28560
rect 39600 28504 40000 28560
rect 0 28168 400 28224
rect 39600 28168 40000 28224
rect 0 27832 400 27888
rect 39600 27832 40000 27888
rect 0 27496 400 27552
rect 39600 27496 40000 27552
rect 0 27160 400 27216
rect 39600 27160 40000 27216
rect 0 26824 400 26880
rect 39600 26824 40000 26880
rect 0 26488 400 26544
rect 39600 26488 40000 26544
rect 0 26152 400 26208
rect 39600 26152 40000 26208
rect 0 25816 400 25872
rect 39600 25816 40000 25872
rect 0 25480 400 25536
rect 39600 25480 40000 25536
rect 0 25144 400 25200
rect 39600 25144 40000 25200
rect 0 24808 400 24864
rect 39600 24808 40000 24864
rect 0 24472 400 24528
rect 39600 24472 40000 24528
rect 0 24136 400 24192
rect 39600 24136 40000 24192
rect 0 23800 400 23856
rect 39600 23800 40000 23856
rect 0 23464 400 23520
rect 39600 23464 40000 23520
rect 0 23128 400 23184
rect 39600 23128 40000 23184
rect 0 22792 400 22848
rect 39600 22792 40000 22848
rect 0 22456 400 22512
rect 39600 22456 40000 22512
rect 0 22120 400 22176
rect 39600 22120 40000 22176
rect 0 21784 400 21840
rect 39600 21784 40000 21840
rect 0 21448 400 21504
rect 39600 21448 40000 21504
rect 0 21112 400 21168
rect 39600 21112 40000 21168
rect 0 20776 400 20832
rect 39600 20776 40000 20832
rect 0 20440 400 20496
rect 39600 20440 40000 20496
rect 0 20104 400 20160
rect 39600 20104 40000 20160
rect 0 19768 400 19824
rect 39600 19768 40000 19824
rect 0 19432 400 19488
rect 39600 19432 40000 19488
rect 0 19096 400 19152
rect 39600 19096 40000 19152
rect 0 18760 400 18816
rect 39600 18760 40000 18816
rect 0 18424 400 18480
rect 39600 18424 40000 18480
rect 0 18088 400 18144
rect 39600 18088 40000 18144
rect 0 17752 400 17808
rect 39600 17752 40000 17808
rect 0 17416 400 17472
rect 39600 17416 40000 17472
rect 0 17080 400 17136
rect 39600 17080 40000 17136
rect 0 16744 400 16800
rect 39600 16744 40000 16800
rect 0 16408 400 16464
rect 39600 16408 40000 16464
rect 0 16072 400 16128
rect 39600 16072 40000 16128
rect 0 15736 400 15792
rect 39600 15736 40000 15792
rect 0 15400 400 15456
rect 39600 15400 40000 15456
rect 0 15064 400 15120
rect 39600 15064 40000 15120
rect 0 14728 400 14784
rect 39600 14728 40000 14784
rect 0 14392 400 14448
rect 39600 14392 40000 14448
rect 0 14056 400 14112
rect 39600 14056 40000 14112
rect 0 13720 400 13776
rect 39600 13720 40000 13776
rect 0 13384 400 13440
rect 39600 13384 40000 13440
rect 0 13048 400 13104
rect 39600 13048 40000 13104
rect 0 12712 400 12768
rect 39600 12712 40000 12768
rect 0 12376 400 12432
rect 39600 12376 40000 12432
rect 0 12040 400 12096
rect 39600 12040 40000 12096
rect 0 11704 400 11760
rect 39600 11704 40000 11760
rect 0 11368 400 11424
rect 39600 11368 40000 11424
rect 0 11032 400 11088
rect 39600 11032 40000 11088
rect 0 10696 400 10752
rect 39600 10696 40000 10752
rect 0 10360 400 10416
rect 39600 10360 40000 10416
rect 0 10024 400 10080
rect 39600 10024 40000 10080
rect 0 9688 400 9744
rect 39600 9688 40000 9744
rect 0 9352 400 9408
rect 39600 9352 40000 9408
rect 0 9016 400 9072
rect 39600 9016 40000 9072
rect 0 8680 400 8736
rect 39600 8680 40000 8736
rect 0 8344 400 8400
rect 39600 8344 40000 8400
rect 0 8008 400 8064
rect 39600 8008 40000 8064
rect 0 7672 400 7728
rect 39600 7672 40000 7728
rect 0 7336 400 7392
rect 39600 7336 40000 7392
rect 0 7000 400 7056
rect 39600 7000 40000 7056
rect 0 6664 400 6720
rect 39600 6664 40000 6720
rect 0 6328 400 6384
rect 39600 6328 40000 6384
rect 0 5992 400 6048
rect 39600 5992 40000 6048
rect 0 5656 400 5712
rect 39600 5656 40000 5712
rect 0 5320 400 5376
rect 39600 5320 40000 5376
rect 0 4984 400 5040
rect 39600 4984 40000 5040
rect 0 4648 400 4704
rect 39600 4648 40000 4704
rect 0 4312 400 4368
rect 39600 4312 40000 4368
rect 0 3976 400 4032
rect 39600 3976 40000 4032
rect 0 3640 400 3696
rect 39600 3640 40000 3696
rect 0 3304 400 3360
rect 39600 3304 40000 3360
rect 0 2968 400 3024
rect 39600 2968 40000 3024
rect 0 2632 400 2688
rect 39600 2632 40000 2688
<< obsm3 >>
rect 400 37326 39634 38430
rect 430 37210 39570 37326
rect 400 36990 39634 37210
rect 430 36874 39570 36990
rect 400 36654 39634 36874
rect 430 36538 39570 36654
rect 400 36318 39634 36538
rect 430 36202 39570 36318
rect 400 35982 39634 36202
rect 430 35866 39570 35982
rect 400 35646 39634 35866
rect 430 35530 39570 35646
rect 400 35310 39634 35530
rect 430 35194 39570 35310
rect 400 34974 39634 35194
rect 430 34858 39570 34974
rect 400 34638 39634 34858
rect 430 34522 39570 34638
rect 400 34302 39634 34522
rect 430 34186 39570 34302
rect 400 33966 39634 34186
rect 430 33850 39570 33966
rect 400 33630 39634 33850
rect 430 33514 39570 33630
rect 400 33294 39634 33514
rect 430 33178 39570 33294
rect 400 32958 39634 33178
rect 430 32842 39570 32958
rect 400 32622 39634 32842
rect 430 32506 39570 32622
rect 400 32286 39634 32506
rect 430 32170 39570 32286
rect 400 31950 39634 32170
rect 430 31834 39570 31950
rect 400 31614 39634 31834
rect 430 31498 39570 31614
rect 400 31278 39634 31498
rect 430 31162 39570 31278
rect 400 30942 39634 31162
rect 430 30826 39570 30942
rect 400 30606 39634 30826
rect 430 30490 39570 30606
rect 400 30270 39634 30490
rect 430 30154 39570 30270
rect 400 29934 39634 30154
rect 430 29818 39570 29934
rect 400 29598 39634 29818
rect 430 29482 39570 29598
rect 400 29262 39634 29482
rect 430 29146 39570 29262
rect 400 28926 39634 29146
rect 430 28810 39570 28926
rect 400 28590 39634 28810
rect 430 28474 39570 28590
rect 400 28254 39634 28474
rect 430 28138 39570 28254
rect 400 27918 39634 28138
rect 430 27802 39570 27918
rect 400 27582 39634 27802
rect 430 27466 39570 27582
rect 400 27246 39634 27466
rect 430 27130 39570 27246
rect 400 26910 39634 27130
rect 430 26794 39570 26910
rect 400 26574 39634 26794
rect 430 26458 39570 26574
rect 400 26238 39634 26458
rect 430 26122 39570 26238
rect 400 25902 39634 26122
rect 430 25786 39570 25902
rect 400 25566 39634 25786
rect 430 25450 39570 25566
rect 400 25230 39634 25450
rect 430 25114 39570 25230
rect 400 24894 39634 25114
rect 430 24778 39570 24894
rect 400 24558 39634 24778
rect 430 24442 39570 24558
rect 400 24222 39634 24442
rect 430 24106 39570 24222
rect 400 23886 39634 24106
rect 430 23770 39570 23886
rect 400 23550 39634 23770
rect 430 23434 39570 23550
rect 400 23214 39634 23434
rect 430 23098 39570 23214
rect 400 22878 39634 23098
rect 430 22762 39570 22878
rect 400 22542 39634 22762
rect 430 22426 39570 22542
rect 400 22206 39634 22426
rect 430 22090 39570 22206
rect 400 21870 39634 22090
rect 430 21754 39570 21870
rect 400 21534 39634 21754
rect 430 21418 39570 21534
rect 400 21198 39634 21418
rect 430 21082 39570 21198
rect 400 20862 39634 21082
rect 430 20746 39570 20862
rect 400 20526 39634 20746
rect 430 20410 39570 20526
rect 400 20190 39634 20410
rect 430 20074 39570 20190
rect 400 19854 39634 20074
rect 430 19738 39570 19854
rect 400 19518 39634 19738
rect 430 19402 39570 19518
rect 400 19182 39634 19402
rect 430 19066 39570 19182
rect 400 18846 39634 19066
rect 430 18730 39570 18846
rect 400 18510 39634 18730
rect 430 18394 39570 18510
rect 400 18174 39634 18394
rect 430 18058 39570 18174
rect 400 17838 39634 18058
rect 430 17722 39570 17838
rect 400 17502 39634 17722
rect 430 17386 39570 17502
rect 400 17166 39634 17386
rect 430 17050 39570 17166
rect 400 16830 39634 17050
rect 430 16714 39570 16830
rect 400 16494 39634 16714
rect 430 16378 39570 16494
rect 400 16158 39634 16378
rect 430 16042 39570 16158
rect 400 15822 39634 16042
rect 430 15706 39570 15822
rect 400 15486 39634 15706
rect 430 15370 39570 15486
rect 400 15150 39634 15370
rect 430 15034 39570 15150
rect 400 14814 39634 15034
rect 430 14698 39570 14814
rect 400 14478 39634 14698
rect 430 14362 39570 14478
rect 400 14142 39634 14362
rect 430 14026 39570 14142
rect 400 13806 39634 14026
rect 430 13690 39570 13806
rect 400 13470 39634 13690
rect 430 13354 39570 13470
rect 400 13134 39634 13354
rect 430 13018 39570 13134
rect 400 12798 39634 13018
rect 430 12682 39570 12798
rect 400 12462 39634 12682
rect 430 12346 39570 12462
rect 400 12126 39634 12346
rect 430 12010 39570 12126
rect 400 11790 39634 12010
rect 430 11674 39570 11790
rect 400 11454 39634 11674
rect 430 11338 39570 11454
rect 400 11118 39634 11338
rect 430 11002 39570 11118
rect 400 10782 39634 11002
rect 430 10666 39570 10782
rect 400 10446 39634 10666
rect 430 10330 39570 10446
rect 400 10110 39634 10330
rect 430 9994 39570 10110
rect 400 9774 39634 9994
rect 430 9658 39570 9774
rect 400 9438 39634 9658
rect 430 9322 39570 9438
rect 400 9102 39634 9322
rect 430 8986 39570 9102
rect 400 8766 39634 8986
rect 430 8650 39570 8766
rect 400 8430 39634 8650
rect 430 8314 39570 8430
rect 400 8094 39634 8314
rect 430 7978 39570 8094
rect 400 7758 39634 7978
rect 430 7642 39570 7758
rect 400 7422 39634 7642
rect 430 7306 39570 7422
rect 400 7086 39634 7306
rect 430 6970 39570 7086
rect 400 6750 39634 6970
rect 430 6634 39570 6750
rect 400 6414 39634 6634
rect 430 6298 39570 6414
rect 400 6078 39634 6298
rect 430 5962 39570 6078
rect 400 5742 39634 5962
rect 430 5626 39570 5742
rect 400 5406 39634 5626
rect 430 5290 39570 5406
rect 400 5070 39634 5290
rect 430 4954 39570 5070
rect 400 4734 39634 4954
rect 430 4618 39570 4734
rect 400 4398 39634 4618
rect 430 4282 39570 4398
rect 400 4062 39634 4282
rect 430 3946 39570 4062
rect 400 3726 39634 3946
rect 430 3610 39570 3726
rect 400 3390 39634 3610
rect 430 3274 39570 3390
rect 400 3054 39634 3274
rect 430 2938 39570 3054
rect 400 2718 39634 2938
rect 430 2602 39570 2718
rect 400 1554 39634 2602
<< metal4 >>
rect 2224 1538 2384 38446
rect 9904 1538 10064 38446
rect 17584 1538 17744 38446
rect 25264 1538 25424 38446
rect 32944 1538 33104 38446
<< labels >>
rlabel metal2 s 36904 0 36960 400 6 io_wbs_ack
port 1 nsew signal output
rlabel metal3 s 39600 36904 40000 36960 6 io_wbs_ack_0
port 2 nsew signal input
rlabel metal3 s 0 36904 400 36960 6 io_wbs_ack_1
port 3 nsew signal input
rlabel metal2 s 2632 0 2688 400 6 io_wbs_adr[0]
port 4 nsew signal input
rlabel metal2 s 5992 0 6048 400 6 io_wbs_adr[10]
port 5 nsew signal input
rlabel metal2 s 6328 0 6384 400 6 io_wbs_adr[11]
port 6 nsew signal input
rlabel metal2 s 6664 0 6720 400 6 io_wbs_adr[12]
port 7 nsew signal input
rlabel metal2 s 7000 0 7056 400 6 io_wbs_adr[13]
port 8 nsew signal input
rlabel metal2 s 7336 0 7392 400 6 io_wbs_adr[14]
port 9 nsew signal input
rlabel metal2 s 7672 0 7728 400 6 io_wbs_adr[15]
port 10 nsew signal input
rlabel metal2 s 8008 0 8064 400 6 io_wbs_adr[16]
port 11 nsew signal input
rlabel metal2 s 8344 0 8400 400 6 io_wbs_adr[17]
port 12 nsew signal input
rlabel metal2 s 8680 0 8736 400 6 io_wbs_adr[18]
port 13 nsew signal input
rlabel metal2 s 9016 0 9072 400 6 io_wbs_adr[19]
port 14 nsew signal input
rlabel metal2 s 2968 0 3024 400 6 io_wbs_adr[1]
port 15 nsew signal input
rlabel metal2 s 9352 0 9408 400 6 io_wbs_adr[20]
port 16 nsew signal input
rlabel metal2 s 9688 0 9744 400 6 io_wbs_adr[21]
port 17 nsew signal input
rlabel metal2 s 10024 0 10080 400 6 io_wbs_adr[22]
port 18 nsew signal input
rlabel metal2 s 10360 0 10416 400 6 io_wbs_adr[23]
port 19 nsew signal input
rlabel metal2 s 10696 0 10752 400 6 io_wbs_adr[24]
port 20 nsew signal input
rlabel metal2 s 11032 0 11088 400 6 io_wbs_adr[25]
port 21 nsew signal input
rlabel metal2 s 11368 0 11424 400 6 io_wbs_adr[26]
port 22 nsew signal input
rlabel metal2 s 11704 0 11760 400 6 io_wbs_adr[27]
port 23 nsew signal input
rlabel metal2 s 12040 0 12096 400 6 io_wbs_adr[28]
port 24 nsew signal input
rlabel metal2 s 12376 0 12432 400 6 io_wbs_adr[29]
port 25 nsew signal input
rlabel metal2 s 3304 0 3360 400 6 io_wbs_adr[2]
port 26 nsew signal input
rlabel metal2 s 12712 0 12768 400 6 io_wbs_adr[30]
port 27 nsew signal input
rlabel metal2 s 13048 0 13104 400 6 io_wbs_adr[31]
port 28 nsew signal input
rlabel metal2 s 3640 0 3696 400 6 io_wbs_adr[3]
port 29 nsew signal input
rlabel metal2 s 3976 0 4032 400 6 io_wbs_adr[4]
port 30 nsew signal input
rlabel metal2 s 4312 0 4368 400 6 io_wbs_adr[5]
port 31 nsew signal input
rlabel metal2 s 4648 0 4704 400 6 io_wbs_adr[6]
port 32 nsew signal input
rlabel metal2 s 4984 0 5040 400 6 io_wbs_adr[7]
port 33 nsew signal input
rlabel metal2 s 5320 0 5376 400 6 io_wbs_adr[8]
port 34 nsew signal input
rlabel metal2 s 5656 0 5712 400 6 io_wbs_adr[9]
port 35 nsew signal input
rlabel metal3 s 39600 2632 40000 2688 6 io_wbs_adr_0[0]
port 36 nsew signal output
rlabel metal3 s 39600 5992 40000 6048 6 io_wbs_adr_0[10]
port 37 nsew signal output
rlabel metal3 s 39600 6328 40000 6384 6 io_wbs_adr_0[11]
port 38 nsew signal output
rlabel metal3 s 39600 6664 40000 6720 6 io_wbs_adr_0[12]
port 39 nsew signal output
rlabel metal3 s 39600 7000 40000 7056 6 io_wbs_adr_0[13]
port 40 nsew signal output
rlabel metal3 s 39600 7336 40000 7392 6 io_wbs_adr_0[14]
port 41 nsew signal output
rlabel metal3 s 39600 7672 40000 7728 6 io_wbs_adr_0[15]
port 42 nsew signal output
rlabel metal3 s 39600 8008 40000 8064 6 io_wbs_adr_0[16]
port 43 nsew signal output
rlabel metal3 s 39600 8344 40000 8400 6 io_wbs_adr_0[17]
port 44 nsew signal output
rlabel metal3 s 39600 8680 40000 8736 6 io_wbs_adr_0[18]
port 45 nsew signal output
rlabel metal3 s 39600 9016 40000 9072 6 io_wbs_adr_0[19]
port 46 nsew signal output
rlabel metal3 s 39600 2968 40000 3024 6 io_wbs_adr_0[1]
port 47 nsew signal output
rlabel metal3 s 39600 9352 40000 9408 6 io_wbs_adr_0[20]
port 48 nsew signal output
rlabel metal3 s 39600 9688 40000 9744 6 io_wbs_adr_0[21]
port 49 nsew signal output
rlabel metal3 s 39600 10024 40000 10080 6 io_wbs_adr_0[22]
port 50 nsew signal output
rlabel metal3 s 39600 10360 40000 10416 6 io_wbs_adr_0[23]
port 51 nsew signal output
rlabel metal3 s 39600 10696 40000 10752 6 io_wbs_adr_0[24]
port 52 nsew signal output
rlabel metal3 s 39600 11032 40000 11088 6 io_wbs_adr_0[25]
port 53 nsew signal output
rlabel metal3 s 39600 11368 40000 11424 6 io_wbs_adr_0[26]
port 54 nsew signal output
rlabel metal3 s 39600 11704 40000 11760 6 io_wbs_adr_0[27]
port 55 nsew signal output
rlabel metal3 s 39600 12040 40000 12096 6 io_wbs_adr_0[28]
port 56 nsew signal output
rlabel metal3 s 39600 12376 40000 12432 6 io_wbs_adr_0[29]
port 57 nsew signal output
rlabel metal3 s 39600 3304 40000 3360 6 io_wbs_adr_0[2]
port 58 nsew signal output
rlabel metal3 s 39600 12712 40000 12768 6 io_wbs_adr_0[30]
port 59 nsew signal output
rlabel metal3 s 39600 13048 40000 13104 6 io_wbs_adr_0[31]
port 60 nsew signal output
rlabel metal3 s 39600 3640 40000 3696 6 io_wbs_adr_0[3]
port 61 nsew signal output
rlabel metal3 s 39600 3976 40000 4032 6 io_wbs_adr_0[4]
port 62 nsew signal output
rlabel metal3 s 39600 4312 40000 4368 6 io_wbs_adr_0[5]
port 63 nsew signal output
rlabel metal3 s 39600 4648 40000 4704 6 io_wbs_adr_0[6]
port 64 nsew signal output
rlabel metal3 s 39600 4984 40000 5040 6 io_wbs_adr_0[7]
port 65 nsew signal output
rlabel metal3 s 39600 5320 40000 5376 6 io_wbs_adr_0[8]
port 66 nsew signal output
rlabel metal3 s 39600 5656 40000 5712 6 io_wbs_adr_0[9]
port 67 nsew signal output
rlabel metal3 s 0 2632 400 2688 6 io_wbs_adr_1[0]
port 68 nsew signal output
rlabel metal3 s 0 5992 400 6048 6 io_wbs_adr_1[10]
port 69 nsew signal output
rlabel metal3 s 0 6328 400 6384 6 io_wbs_adr_1[11]
port 70 nsew signal output
rlabel metal3 s 0 6664 400 6720 6 io_wbs_adr_1[12]
port 71 nsew signal output
rlabel metal3 s 0 7000 400 7056 6 io_wbs_adr_1[13]
port 72 nsew signal output
rlabel metal3 s 0 7336 400 7392 6 io_wbs_adr_1[14]
port 73 nsew signal output
rlabel metal3 s 0 7672 400 7728 6 io_wbs_adr_1[15]
port 74 nsew signal output
rlabel metal3 s 0 8008 400 8064 6 io_wbs_adr_1[16]
port 75 nsew signal output
rlabel metal3 s 0 8344 400 8400 6 io_wbs_adr_1[17]
port 76 nsew signal output
rlabel metal3 s 0 8680 400 8736 6 io_wbs_adr_1[18]
port 77 nsew signal output
rlabel metal3 s 0 9016 400 9072 6 io_wbs_adr_1[19]
port 78 nsew signal output
rlabel metal3 s 0 2968 400 3024 6 io_wbs_adr_1[1]
port 79 nsew signal output
rlabel metal3 s 0 9352 400 9408 6 io_wbs_adr_1[20]
port 80 nsew signal output
rlabel metal3 s 0 9688 400 9744 6 io_wbs_adr_1[21]
port 81 nsew signal output
rlabel metal3 s 0 10024 400 10080 6 io_wbs_adr_1[22]
port 82 nsew signal output
rlabel metal3 s 0 10360 400 10416 6 io_wbs_adr_1[23]
port 83 nsew signal output
rlabel metal3 s 0 10696 400 10752 6 io_wbs_adr_1[24]
port 84 nsew signal output
rlabel metal3 s 0 11032 400 11088 6 io_wbs_adr_1[25]
port 85 nsew signal output
rlabel metal3 s 0 11368 400 11424 6 io_wbs_adr_1[26]
port 86 nsew signal output
rlabel metal3 s 0 11704 400 11760 6 io_wbs_adr_1[27]
port 87 nsew signal output
rlabel metal3 s 0 12040 400 12096 6 io_wbs_adr_1[28]
port 88 nsew signal output
rlabel metal3 s 0 12376 400 12432 6 io_wbs_adr_1[29]
port 89 nsew signal output
rlabel metal3 s 0 3304 400 3360 6 io_wbs_adr_1[2]
port 90 nsew signal output
rlabel metal3 s 0 12712 400 12768 6 io_wbs_adr_1[30]
port 91 nsew signal output
rlabel metal3 s 0 13048 400 13104 6 io_wbs_adr_1[31]
port 92 nsew signal output
rlabel metal3 s 0 3640 400 3696 6 io_wbs_adr_1[3]
port 93 nsew signal output
rlabel metal3 s 0 3976 400 4032 6 io_wbs_adr_1[4]
port 94 nsew signal output
rlabel metal3 s 0 4312 400 4368 6 io_wbs_adr_1[5]
port 95 nsew signal output
rlabel metal3 s 0 4648 400 4704 6 io_wbs_adr_1[6]
port 96 nsew signal output
rlabel metal3 s 0 4984 400 5040 6 io_wbs_adr_1[7]
port 97 nsew signal output
rlabel metal3 s 0 5320 400 5376 6 io_wbs_adr_1[8]
port 98 nsew signal output
rlabel metal3 s 0 5656 400 5712 6 io_wbs_adr_1[9]
port 99 nsew signal output
rlabel metal2 s 37240 0 37296 400 6 io_wbs_cyc
port 100 nsew signal input
rlabel metal3 s 39600 37240 40000 37296 6 io_wbs_cyc_0
port 101 nsew signal output
rlabel metal3 s 0 37240 400 37296 6 io_wbs_cyc_1
port 102 nsew signal output
rlabel metal2 s 24136 0 24192 400 6 io_wbs_datrd[0]
port 103 nsew signal output
rlabel metal2 s 27496 0 27552 400 6 io_wbs_datrd[10]
port 104 nsew signal output
rlabel metal2 s 27832 0 27888 400 6 io_wbs_datrd[11]
port 105 nsew signal output
rlabel metal2 s 28168 0 28224 400 6 io_wbs_datrd[12]
port 106 nsew signal output
rlabel metal2 s 28504 0 28560 400 6 io_wbs_datrd[13]
port 107 nsew signal output
rlabel metal2 s 28840 0 28896 400 6 io_wbs_datrd[14]
port 108 nsew signal output
rlabel metal2 s 29176 0 29232 400 6 io_wbs_datrd[15]
port 109 nsew signal output
rlabel metal2 s 29512 0 29568 400 6 io_wbs_datrd[16]
port 110 nsew signal output
rlabel metal2 s 29848 0 29904 400 6 io_wbs_datrd[17]
port 111 nsew signal output
rlabel metal2 s 30184 0 30240 400 6 io_wbs_datrd[18]
port 112 nsew signal output
rlabel metal2 s 30520 0 30576 400 6 io_wbs_datrd[19]
port 113 nsew signal output
rlabel metal2 s 24472 0 24528 400 6 io_wbs_datrd[1]
port 114 nsew signal output
rlabel metal2 s 30856 0 30912 400 6 io_wbs_datrd[20]
port 115 nsew signal output
rlabel metal2 s 31192 0 31248 400 6 io_wbs_datrd[21]
port 116 nsew signal output
rlabel metal2 s 31528 0 31584 400 6 io_wbs_datrd[22]
port 117 nsew signal output
rlabel metal2 s 31864 0 31920 400 6 io_wbs_datrd[23]
port 118 nsew signal output
rlabel metal2 s 32200 0 32256 400 6 io_wbs_datrd[24]
port 119 nsew signal output
rlabel metal2 s 32536 0 32592 400 6 io_wbs_datrd[25]
port 120 nsew signal output
rlabel metal2 s 32872 0 32928 400 6 io_wbs_datrd[26]
port 121 nsew signal output
rlabel metal2 s 33208 0 33264 400 6 io_wbs_datrd[27]
port 122 nsew signal output
rlabel metal2 s 33544 0 33600 400 6 io_wbs_datrd[28]
port 123 nsew signal output
rlabel metal2 s 33880 0 33936 400 6 io_wbs_datrd[29]
port 124 nsew signal output
rlabel metal2 s 24808 0 24864 400 6 io_wbs_datrd[2]
port 125 nsew signal output
rlabel metal2 s 34216 0 34272 400 6 io_wbs_datrd[30]
port 126 nsew signal output
rlabel metal2 s 34552 0 34608 400 6 io_wbs_datrd[31]
port 127 nsew signal output
rlabel metal2 s 25144 0 25200 400 6 io_wbs_datrd[3]
port 128 nsew signal output
rlabel metal2 s 25480 0 25536 400 6 io_wbs_datrd[4]
port 129 nsew signal output
rlabel metal2 s 25816 0 25872 400 6 io_wbs_datrd[5]
port 130 nsew signal output
rlabel metal2 s 26152 0 26208 400 6 io_wbs_datrd[6]
port 131 nsew signal output
rlabel metal2 s 26488 0 26544 400 6 io_wbs_datrd[7]
port 132 nsew signal output
rlabel metal2 s 26824 0 26880 400 6 io_wbs_datrd[8]
port 133 nsew signal output
rlabel metal2 s 27160 0 27216 400 6 io_wbs_datrd[9]
port 134 nsew signal output
rlabel metal3 s 39600 24136 40000 24192 6 io_wbs_datrd_0[0]
port 135 nsew signal input
rlabel metal3 s 39600 27496 40000 27552 6 io_wbs_datrd_0[10]
port 136 nsew signal input
rlabel metal3 s 39600 27832 40000 27888 6 io_wbs_datrd_0[11]
port 137 nsew signal input
rlabel metal3 s 39600 28168 40000 28224 6 io_wbs_datrd_0[12]
port 138 nsew signal input
rlabel metal3 s 39600 28504 40000 28560 6 io_wbs_datrd_0[13]
port 139 nsew signal input
rlabel metal3 s 39600 28840 40000 28896 6 io_wbs_datrd_0[14]
port 140 nsew signal input
rlabel metal3 s 39600 29176 40000 29232 6 io_wbs_datrd_0[15]
port 141 nsew signal input
rlabel metal3 s 39600 29512 40000 29568 6 io_wbs_datrd_0[16]
port 142 nsew signal input
rlabel metal3 s 39600 29848 40000 29904 6 io_wbs_datrd_0[17]
port 143 nsew signal input
rlabel metal3 s 39600 30184 40000 30240 6 io_wbs_datrd_0[18]
port 144 nsew signal input
rlabel metal3 s 39600 30520 40000 30576 6 io_wbs_datrd_0[19]
port 145 nsew signal input
rlabel metal3 s 39600 24472 40000 24528 6 io_wbs_datrd_0[1]
port 146 nsew signal input
rlabel metal3 s 39600 30856 40000 30912 6 io_wbs_datrd_0[20]
port 147 nsew signal input
rlabel metal3 s 39600 31192 40000 31248 6 io_wbs_datrd_0[21]
port 148 nsew signal input
rlabel metal3 s 39600 31528 40000 31584 6 io_wbs_datrd_0[22]
port 149 nsew signal input
rlabel metal3 s 39600 31864 40000 31920 6 io_wbs_datrd_0[23]
port 150 nsew signal input
rlabel metal3 s 39600 32200 40000 32256 6 io_wbs_datrd_0[24]
port 151 nsew signal input
rlabel metal3 s 39600 32536 40000 32592 6 io_wbs_datrd_0[25]
port 152 nsew signal input
rlabel metal3 s 39600 32872 40000 32928 6 io_wbs_datrd_0[26]
port 153 nsew signal input
rlabel metal3 s 39600 33208 40000 33264 6 io_wbs_datrd_0[27]
port 154 nsew signal input
rlabel metal3 s 39600 33544 40000 33600 6 io_wbs_datrd_0[28]
port 155 nsew signal input
rlabel metal3 s 39600 33880 40000 33936 6 io_wbs_datrd_0[29]
port 156 nsew signal input
rlabel metal3 s 39600 24808 40000 24864 6 io_wbs_datrd_0[2]
port 157 nsew signal input
rlabel metal3 s 39600 34216 40000 34272 6 io_wbs_datrd_0[30]
port 158 nsew signal input
rlabel metal3 s 39600 34552 40000 34608 6 io_wbs_datrd_0[31]
port 159 nsew signal input
rlabel metal3 s 39600 25144 40000 25200 6 io_wbs_datrd_0[3]
port 160 nsew signal input
rlabel metal3 s 39600 25480 40000 25536 6 io_wbs_datrd_0[4]
port 161 nsew signal input
rlabel metal3 s 39600 25816 40000 25872 6 io_wbs_datrd_0[5]
port 162 nsew signal input
rlabel metal3 s 39600 26152 40000 26208 6 io_wbs_datrd_0[6]
port 163 nsew signal input
rlabel metal3 s 39600 26488 40000 26544 6 io_wbs_datrd_0[7]
port 164 nsew signal input
rlabel metal3 s 39600 26824 40000 26880 6 io_wbs_datrd_0[8]
port 165 nsew signal input
rlabel metal3 s 39600 27160 40000 27216 6 io_wbs_datrd_0[9]
port 166 nsew signal input
rlabel metal3 s 0 24136 400 24192 6 io_wbs_datrd_1[0]
port 167 nsew signal input
rlabel metal3 s 0 27496 400 27552 6 io_wbs_datrd_1[10]
port 168 nsew signal input
rlabel metal3 s 0 27832 400 27888 6 io_wbs_datrd_1[11]
port 169 nsew signal input
rlabel metal3 s 0 28168 400 28224 6 io_wbs_datrd_1[12]
port 170 nsew signal input
rlabel metal3 s 0 28504 400 28560 6 io_wbs_datrd_1[13]
port 171 nsew signal input
rlabel metal3 s 0 28840 400 28896 6 io_wbs_datrd_1[14]
port 172 nsew signal input
rlabel metal3 s 0 29176 400 29232 6 io_wbs_datrd_1[15]
port 173 nsew signal input
rlabel metal3 s 0 29512 400 29568 6 io_wbs_datrd_1[16]
port 174 nsew signal input
rlabel metal3 s 0 29848 400 29904 6 io_wbs_datrd_1[17]
port 175 nsew signal input
rlabel metal3 s 0 30184 400 30240 6 io_wbs_datrd_1[18]
port 176 nsew signal input
rlabel metal3 s 0 30520 400 30576 6 io_wbs_datrd_1[19]
port 177 nsew signal input
rlabel metal3 s 0 24472 400 24528 6 io_wbs_datrd_1[1]
port 178 nsew signal input
rlabel metal3 s 0 30856 400 30912 6 io_wbs_datrd_1[20]
port 179 nsew signal input
rlabel metal3 s 0 31192 400 31248 6 io_wbs_datrd_1[21]
port 180 nsew signal input
rlabel metal3 s 0 31528 400 31584 6 io_wbs_datrd_1[22]
port 181 nsew signal input
rlabel metal3 s 0 31864 400 31920 6 io_wbs_datrd_1[23]
port 182 nsew signal input
rlabel metal3 s 0 32200 400 32256 6 io_wbs_datrd_1[24]
port 183 nsew signal input
rlabel metal3 s 0 32536 400 32592 6 io_wbs_datrd_1[25]
port 184 nsew signal input
rlabel metal3 s 0 32872 400 32928 6 io_wbs_datrd_1[26]
port 185 nsew signal input
rlabel metal3 s 0 33208 400 33264 6 io_wbs_datrd_1[27]
port 186 nsew signal input
rlabel metal3 s 0 33544 400 33600 6 io_wbs_datrd_1[28]
port 187 nsew signal input
rlabel metal3 s 0 33880 400 33936 6 io_wbs_datrd_1[29]
port 188 nsew signal input
rlabel metal3 s 0 24808 400 24864 6 io_wbs_datrd_1[2]
port 189 nsew signal input
rlabel metal3 s 0 34216 400 34272 6 io_wbs_datrd_1[30]
port 190 nsew signal input
rlabel metal3 s 0 34552 400 34608 6 io_wbs_datrd_1[31]
port 191 nsew signal input
rlabel metal3 s 0 25144 400 25200 6 io_wbs_datrd_1[3]
port 192 nsew signal input
rlabel metal3 s 0 25480 400 25536 6 io_wbs_datrd_1[4]
port 193 nsew signal input
rlabel metal3 s 0 25816 400 25872 6 io_wbs_datrd_1[5]
port 194 nsew signal input
rlabel metal3 s 0 26152 400 26208 6 io_wbs_datrd_1[6]
port 195 nsew signal input
rlabel metal3 s 0 26488 400 26544 6 io_wbs_datrd_1[7]
port 196 nsew signal input
rlabel metal3 s 0 26824 400 26880 6 io_wbs_datrd_1[8]
port 197 nsew signal input
rlabel metal3 s 0 27160 400 27216 6 io_wbs_datrd_1[9]
port 198 nsew signal input
rlabel metal2 s 13384 0 13440 400 6 io_wbs_datwr[0]
port 199 nsew signal input
rlabel metal2 s 16744 0 16800 400 6 io_wbs_datwr[10]
port 200 nsew signal input
rlabel metal2 s 17080 0 17136 400 6 io_wbs_datwr[11]
port 201 nsew signal input
rlabel metal2 s 17416 0 17472 400 6 io_wbs_datwr[12]
port 202 nsew signal input
rlabel metal2 s 17752 0 17808 400 6 io_wbs_datwr[13]
port 203 nsew signal input
rlabel metal2 s 18088 0 18144 400 6 io_wbs_datwr[14]
port 204 nsew signal input
rlabel metal2 s 18424 0 18480 400 6 io_wbs_datwr[15]
port 205 nsew signal input
rlabel metal2 s 18760 0 18816 400 6 io_wbs_datwr[16]
port 206 nsew signal input
rlabel metal2 s 19096 0 19152 400 6 io_wbs_datwr[17]
port 207 nsew signal input
rlabel metal2 s 19432 0 19488 400 6 io_wbs_datwr[18]
port 208 nsew signal input
rlabel metal2 s 19768 0 19824 400 6 io_wbs_datwr[19]
port 209 nsew signal input
rlabel metal2 s 13720 0 13776 400 6 io_wbs_datwr[1]
port 210 nsew signal input
rlabel metal2 s 20104 0 20160 400 6 io_wbs_datwr[20]
port 211 nsew signal input
rlabel metal2 s 20440 0 20496 400 6 io_wbs_datwr[21]
port 212 nsew signal input
rlabel metal2 s 20776 0 20832 400 6 io_wbs_datwr[22]
port 213 nsew signal input
rlabel metal2 s 21112 0 21168 400 6 io_wbs_datwr[23]
port 214 nsew signal input
rlabel metal2 s 21448 0 21504 400 6 io_wbs_datwr[24]
port 215 nsew signal input
rlabel metal2 s 21784 0 21840 400 6 io_wbs_datwr[25]
port 216 nsew signal input
rlabel metal2 s 22120 0 22176 400 6 io_wbs_datwr[26]
port 217 nsew signal input
rlabel metal2 s 22456 0 22512 400 6 io_wbs_datwr[27]
port 218 nsew signal input
rlabel metal2 s 22792 0 22848 400 6 io_wbs_datwr[28]
port 219 nsew signal input
rlabel metal2 s 23128 0 23184 400 6 io_wbs_datwr[29]
port 220 nsew signal input
rlabel metal2 s 14056 0 14112 400 6 io_wbs_datwr[2]
port 221 nsew signal input
rlabel metal2 s 23464 0 23520 400 6 io_wbs_datwr[30]
port 222 nsew signal input
rlabel metal2 s 23800 0 23856 400 6 io_wbs_datwr[31]
port 223 nsew signal input
rlabel metal2 s 14392 0 14448 400 6 io_wbs_datwr[3]
port 224 nsew signal input
rlabel metal2 s 14728 0 14784 400 6 io_wbs_datwr[4]
port 225 nsew signal input
rlabel metal2 s 15064 0 15120 400 6 io_wbs_datwr[5]
port 226 nsew signal input
rlabel metal2 s 15400 0 15456 400 6 io_wbs_datwr[6]
port 227 nsew signal input
rlabel metal2 s 15736 0 15792 400 6 io_wbs_datwr[7]
port 228 nsew signal input
rlabel metal2 s 16072 0 16128 400 6 io_wbs_datwr[8]
port 229 nsew signal input
rlabel metal2 s 16408 0 16464 400 6 io_wbs_datwr[9]
port 230 nsew signal input
rlabel metal3 s 39600 13384 40000 13440 6 io_wbs_datwr_0[0]
port 231 nsew signal output
rlabel metal3 s 39600 16744 40000 16800 6 io_wbs_datwr_0[10]
port 232 nsew signal output
rlabel metal3 s 39600 17080 40000 17136 6 io_wbs_datwr_0[11]
port 233 nsew signal output
rlabel metal3 s 39600 17416 40000 17472 6 io_wbs_datwr_0[12]
port 234 nsew signal output
rlabel metal3 s 39600 17752 40000 17808 6 io_wbs_datwr_0[13]
port 235 nsew signal output
rlabel metal3 s 39600 18088 40000 18144 6 io_wbs_datwr_0[14]
port 236 nsew signal output
rlabel metal3 s 39600 18424 40000 18480 6 io_wbs_datwr_0[15]
port 237 nsew signal output
rlabel metal3 s 39600 18760 40000 18816 6 io_wbs_datwr_0[16]
port 238 nsew signal output
rlabel metal3 s 39600 19096 40000 19152 6 io_wbs_datwr_0[17]
port 239 nsew signal output
rlabel metal3 s 39600 19432 40000 19488 6 io_wbs_datwr_0[18]
port 240 nsew signal output
rlabel metal3 s 39600 19768 40000 19824 6 io_wbs_datwr_0[19]
port 241 nsew signal output
rlabel metal3 s 39600 13720 40000 13776 6 io_wbs_datwr_0[1]
port 242 nsew signal output
rlabel metal3 s 39600 20104 40000 20160 6 io_wbs_datwr_0[20]
port 243 nsew signal output
rlabel metal3 s 39600 20440 40000 20496 6 io_wbs_datwr_0[21]
port 244 nsew signal output
rlabel metal3 s 39600 20776 40000 20832 6 io_wbs_datwr_0[22]
port 245 nsew signal output
rlabel metal3 s 39600 21112 40000 21168 6 io_wbs_datwr_0[23]
port 246 nsew signal output
rlabel metal3 s 39600 21448 40000 21504 6 io_wbs_datwr_0[24]
port 247 nsew signal output
rlabel metal3 s 39600 21784 40000 21840 6 io_wbs_datwr_0[25]
port 248 nsew signal output
rlabel metal3 s 39600 22120 40000 22176 6 io_wbs_datwr_0[26]
port 249 nsew signal output
rlabel metal3 s 39600 22456 40000 22512 6 io_wbs_datwr_0[27]
port 250 nsew signal output
rlabel metal3 s 39600 22792 40000 22848 6 io_wbs_datwr_0[28]
port 251 nsew signal output
rlabel metal3 s 39600 23128 40000 23184 6 io_wbs_datwr_0[29]
port 252 nsew signal output
rlabel metal3 s 39600 14056 40000 14112 6 io_wbs_datwr_0[2]
port 253 nsew signal output
rlabel metal3 s 39600 23464 40000 23520 6 io_wbs_datwr_0[30]
port 254 nsew signal output
rlabel metal3 s 39600 23800 40000 23856 6 io_wbs_datwr_0[31]
port 255 nsew signal output
rlabel metal3 s 39600 14392 40000 14448 6 io_wbs_datwr_0[3]
port 256 nsew signal output
rlabel metal3 s 39600 14728 40000 14784 6 io_wbs_datwr_0[4]
port 257 nsew signal output
rlabel metal3 s 39600 15064 40000 15120 6 io_wbs_datwr_0[5]
port 258 nsew signal output
rlabel metal3 s 39600 15400 40000 15456 6 io_wbs_datwr_0[6]
port 259 nsew signal output
rlabel metal3 s 39600 15736 40000 15792 6 io_wbs_datwr_0[7]
port 260 nsew signal output
rlabel metal3 s 39600 16072 40000 16128 6 io_wbs_datwr_0[8]
port 261 nsew signal output
rlabel metal3 s 39600 16408 40000 16464 6 io_wbs_datwr_0[9]
port 262 nsew signal output
rlabel metal3 s 0 13384 400 13440 6 io_wbs_datwr_1[0]
port 263 nsew signal output
rlabel metal3 s 0 16744 400 16800 6 io_wbs_datwr_1[10]
port 264 nsew signal output
rlabel metal3 s 0 17080 400 17136 6 io_wbs_datwr_1[11]
port 265 nsew signal output
rlabel metal3 s 0 17416 400 17472 6 io_wbs_datwr_1[12]
port 266 nsew signal output
rlabel metal3 s 0 17752 400 17808 6 io_wbs_datwr_1[13]
port 267 nsew signal output
rlabel metal3 s 0 18088 400 18144 6 io_wbs_datwr_1[14]
port 268 nsew signal output
rlabel metal3 s 0 18424 400 18480 6 io_wbs_datwr_1[15]
port 269 nsew signal output
rlabel metal3 s 0 18760 400 18816 6 io_wbs_datwr_1[16]
port 270 nsew signal output
rlabel metal3 s 0 19096 400 19152 6 io_wbs_datwr_1[17]
port 271 nsew signal output
rlabel metal3 s 0 19432 400 19488 6 io_wbs_datwr_1[18]
port 272 nsew signal output
rlabel metal3 s 0 19768 400 19824 6 io_wbs_datwr_1[19]
port 273 nsew signal output
rlabel metal3 s 0 13720 400 13776 6 io_wbs_datwr_1[1]
port 274 nsew signal output
rlabel metal3 s 0 20104 400 20160 6 io_wbs_datwr_1[20]
port 275 nsew signal output
rlabel metal3 s 0 20440 400 20496 6 io_wbs_datwr_1[21]
port 276 nsew signal output
rlabel metal3 s 0 20776 400 20832 6 io_wbs_datwr_1[22]
port 277 nsew signal output
rlabel metal3 s 0 21112 400 21168 6 io_wbs_datwr_1[23]
port 278 nsew signal output
rlabel metal3 s 0 21448 400 21504 6 io_wbs_datwr_1[24]
port 279 nsew signal output
rlabel metal3 s 0 21784 400 21840 6 io_wbs_datwr_1[25]
port 280 nsew signal output
rlabel metal3 s 0 22120 400 22176 6 io_wbs_datwr_1[26]
port 281 nsew signal output
rlabel metal3 s 0 22456 400 22512 6 io_wbs_datwr_1[27]
port 282 nsew signal output
rlabel metal3 s 0 22792 400 22848 6 io_wbs_datwr_1[28]
port 283 nsew signal output
rlabel metal3 s 0 23128 400 23184 6 io_wbs_datwr_1[29]
port 284 nsew signal output
rlabel metal3 s 0 14056 400 14112 6 io_wbs_datwr_1[2]
port 285 nsew signal output
rlabel metal3 s 0 23464 400 23520 6 io_wbs_datwr_1[30]
port 286 nsew signal output
rlabel metal3 s 0 23800 400 23856 6 io_wbs_datwr_1[31]
port 287 nsew signal output
rlabel metal3 s 0 14392 400 14448 6 io_wbs_datwr_1[3]
port 288 nsew signal output
rlabel metal3 s 0 14728 400 14784 6 io_wbs_datwr_1[4]
port 289 nsew signal output
rlabel metal3 s 0 15064 400 15120 6 io_wbs_datwr_1[5]
port 290 nsew signal output
rlabel metal3 s 0 15400 400 15456 6 io_wbs_datwr_1[6]
port 291 nsew signal output
rlabel metal3 s 0 15736 400 15792 6 io_wbs_datwr_1[7]
port 292 nsew signal output
rlabel metal3 s 0 16072 400 16128 6 io_wbs_datwr_1[8]
port 293 nsew signal output
rlabel metal3 s 0 16408 400 16464 6 io_wbs_datwr_1[9]
port 294 nsew signal output
rlabel metal2 s 35224 0 35280 400 6 io_wbs_sel[0]
port 295 nsew signal input
rlabel metal2 s 35560 0 35616 400 6 io_wbs_sel[1]
port 296 nsew signal input
rlabel metal2 s 35896 0 35952 400 6 io_wbs_sel[2]
port 297 nsew signal input
rlabel metal2 s 36232 0 36288 400 6 io_wbs_sel[3]
port 298 nsew signal input
rlabel metal3 s 39600 35224 40000 35280 6 io_wbs_sel_0[0]
port 299 nsew signal output
rlabel metal3 s 39600 35560 40000 35616 6 io_wbs_sel_0[1]
port 300 nsew signal output
rlabel metal3 s 39600 35896 40000 35952 6 io_wbs_sel_0[2]
port 301 nsew signal output
rlabel metal3 s 39600 36232 40000 36288 6 io_wbs_sel_0[3]
port 302 nsew signal output
rlabel metal3 s 0 35224 400 35280 6 io_wbs_sel_1[0]
port 303 nsew signal output
rlabel metal3 s 0 35560 400 35616 6 io_wbs_sel_1[1]
port 304 nsew signal output
rlabel metal3 s 0 35896 400 35952 6 io_wbs_sel_1[2]
port 305 nsew signal output
rlabel metal3 s 0 36232 400 36288 6 io_wbs_sel_1[3]
port 306 nsew signal output
rlabel metal2 s 36568 0 36624 400 6 io_wbs_stb
port 307 nsew signal input
rlabel metal3 s 39600 36568 40000 36624 6 io_wbs_stb_0
port 308 nsew signal output
rlabel metal3 s 0 36568 400 36624 6 io_wbs_stb_1
port 309 nsew signal output
rlabel metal2 s 34888 0 34944 400 6 io_wbs_we
port 310 nsew signal input
rlabel metal3 s 39600 34888 40000 34944 6 io_wbs_we_0
port 311 nsew signal output
rlabel metal3 s 0 34888 400 34944 6 io_wbs_we_1
port 312 nsew signal output
rlabel metal4 s 2224 1538 2384 38446 6 vdd
port 313 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 38446 6 vdd
port 313 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 38446 6 vdd
port 313 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 38446 6 vss
port 314 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 38446 6 vss
port 314 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1534642
string GDS_FILE /home/leo/Dokumente/the-final-workspace/caravel_user_project/openlane/wb_mux/runs/22_12_05_16_44/results/signoff/wb_mux.magic.gds
string GDS_START 87178
<< end >>

