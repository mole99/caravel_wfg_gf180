VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO merge_memory
  CLASS BLOCK ;
  FOREIGN merge_memory ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 200.000 ;
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 10.080 750.000 10.640 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 14.560 750.000 15.120 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 19.040 750.000 19.600 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 23.520 750.000 24.080 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 28.000 750.000 28.560 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 32.480 750.000 33.040 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 36.960 750.000 37.520 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 41.440 750.000 42.000 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 45.920 750.000 46.480 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 50.400 750.000 50.960 ;
    END
  END addr[9]
  PIN addr_mem0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.160 0.000 34.720 4.000 ;
    END
  END addr_mem0[0]
  PIN addr_mem0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 0.000 43.120 4.000 ;
    END
  END addr_mem0[1]
  PIN addr_mem0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.960 0.000 51.520 4.000 ;
    END
  END addr_mem0[2]
  PIN addr_mem0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.920 4.000 ;
    END
  END addr_mem0[3]
  PIN addr_mem0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.760 0.000 68.320 4.000 ;
    END
  END addr_mem0[4]
  PIN addr_mem0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 0.000 76.720 4.000 ;
    END
  END addr_mem0[5]
  PIN addr_mem0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.560 0.000 85.120 4.000 ;
    END
  END addr_mem0[6]
  PIN addr_mem0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 0.000 93.520 4.000 ;
    END
  END addr_mem0[7]
  PIN addr_mem0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.360 0.000 101.920 4.000 ;
    END
  END addr_mem0[8]
  PIN addr_mem1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.960 0.000 387.520 4.000 ;
    END
  END addr_mem1[0]
  PIN addr_mem1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 395.360 0.000 395.920 4.000 ;
    END
  END addr_mem1[1]
  PIN addr_mem1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.760 0.000 404.320 4.000 ;
    END
  END addr_mem1[2]
  PIN addr_mem1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 412.160 0.000 412.720 4.000 ;
    END
  END addr_mem1[3]
  PIN addr_mem1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.560 0.000 421.120 4.000 ;
    END
  END addr_mem1[4]
  PIN addr_mem1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 428.960 0.000 429.520 4.000 ;
    END
  END addr_mem1[5]
  PIN addr_mem1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.360 0.000 437.920 4.000 ;
    END
  END addr_mem1[6]
  PIN addr_mem1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 0.000 446.320 4.000 ;
    END
  END addr_mem1[7]
  PIN addr_mem1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 454.160 0.000 454.720 4.000 ;
    END
  END addr_mem1[8]
  PIN csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 5.600 750.000 6.160 ;
    END
  END csb
  PIN csb_mem0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END csb_mem0
  PIN csb_mem1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 0.000 379.120 4.000 ;
    END
  END csb_mem1
  PIN dout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 54.880 750.000 55.440 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 99.680 750.000 100.240 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 104.160 750.000 104.720 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 108.640 750.000 109.200 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 113.120 750.000 113.680 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 117.600 750.000 118.160 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 122.080 750.000 122.640 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 126.560 750.000 127.120 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 131.040 750.000 131.600 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 135.520 750.000 136.080 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 140.000 750.000 140.560 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 59.360 750.000 59.920 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 144.480 750.000 145.040 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 148.960 750.000 149.520 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 153.440 750.000 154.000 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 157.920 750.000 158.480 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 162.400 750.000 162.960 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 166.880 750.000 167.440 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 171.360 750.000 171.920 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 175.840 750.000 176.400 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 180.320 750.000 180.880 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 184.800 750.000 185.360 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 63.840 750.000 64.400 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 189.280 750.000 189.840 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 193.760 750.000 194.320 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 68.320 750.000 68.880 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 72.800 750.000 73.360 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 77.280 750.000 77.840 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 81.760 750.000 82.320 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 86.240 750.000 86.800 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 90.720 750.000 91.280 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 746.000 95.200 750.000 95.760 ;
    END
  END dout[9]
  PIN dout_mem0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 0.000 110.320 4.000 ;
    END
  END dout_mem0[0]
  PIN dout_mem0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 0.000 194.320 4.000 ;
    END
  END dout_mem0[10]
  PIN dout_mem0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 202.160 0.000 202.720 4.000 ;
    END
  END dout_mem0[11]
  PIN dout_mem0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 0.000 211.120 4.000 ;
    END
  END dout_mem0[12]
  PIN dout_mem0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.960 0.000 219.520 4.000 ;
    END
  END dout_mem0[13]
  PIN dout_mem0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 0.000 227.920 4.000 ;
    END
  END dout_mem0[14]
  PIN dout_mem0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.760 0.000 236.320 4.000 ;
    END
  END dout_mem0[15]
  PIN dout_mem0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 0.000 244.720 4.000 ;
    END
  END dout_mem0[16]
  PIN dout_mem0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.560 0.000 253.120 4.000 ;
    END
  END dout_mem0[17]
  PIN dout_mem0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 0.000 261.520 4.000 ;
    END
  END dout_mem0[18]
  PIN dout_mem0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.360 0.000 269.920 4.000 ;
    END
  END dout_mem0[19]
  PIN dout_mem0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 118.160 0.000 118.720 4.000 ;
    END
  END dout_mem0[1]
  PIN dout_mem0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 0.000 278.320 4.000 ;
    END
  END dout_mem0[20]
  PIN dout_mem0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 286.160 0.000 286.720 4.000 ;
    END
  END dout_mem0[21]
  PIN dout_mem0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 294.560 0.000 295.120 4.000 ;
    END
  END dout_mem0[22]
  PIN dout_mem0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.960 0.000 303.520 4.000 ;
    END
  END dout_mem0[23]
  PIN dout_mem0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 0.000 311.920 4.000 ;
    END
  END dout_mem0[24]
  PIN dout_mem0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.760 0.000 320.320 4.000 ;
    END
  END dout_mem0[25]
  PIN dout_mem0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 0.000 328.720 4.000 ;
    END
  END dout_mem0[26]
  PIN dout_mem0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.560 0.000 337.120 4.000 ;
    END
  END dout_mem0[27]
  PIN dout_mem0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 344.960 0.000 345.520 4.000 ;
    END
  END dout_mem0[28]
  PIN dout_mem0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 353.360 0.000 353.920 4.000 ;
    END
  END dout_mem0[29]
  PIN dout_mem0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 4.000 ;
    END
  END dout_mem0[2]
  PIN dout_mem0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 361.760 0.000 362.320 4.000 ;
    END
  END dout_mem0[30]
  PIN dout_mem0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 370.160 0.000 370.720 4.000 ;
    END
  END dout_mem0[31]
  PIN dout_mem0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.960 0.000 135.520 4.000 ;
    END
  END dout_mem0[3]
  PIN dout_mem0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 0.000 143.920 4.000 ;
    END
  END dout_mem0[4]
  PIN dout_mem0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.760 0.000 152.320 4.000 ;
    END
  END dout_mem0[5]
  PIN dout_mem0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 0.000 160.720 4.000 ;
    END
  END dout_mem0[6]
  PIN dout_mem0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.560 0.000 169.120 4.000 ;
    END
  END dout_mem0[7]
  PIN dout_mem0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 0.000 177.520 4.000 ;
    END
  END dout_mem0[8]
  PIN dout_mem0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 185.360 0.000 185.920 4.000 ;
    END
  END dout_mem0[9]
  PIN dout_mem1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 462.560 0.000 463.120 4.000 ;
    END
  END dout_mem1[0]
  PIN dout_mem1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 546.560 0.000 547.120 4.000 ;
    END
  END dout_mem1[10]
  PIN dout_mem1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.960 0.000 555.520 4.000 ;
    END
  END dout_mem1[11]
  PIN dout_mem1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 563.360 0.000 563.920 4.000 ;
    END
  END dout_mem1[12]
  PIN dout_mem1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.760 0.000 572.320 4.000 ;
    END
  END dout_mem1[13]
  PIN dout_mem1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 0.000 580.720 4.000 ;
    END
  END dout_mem1[14]
  PIN dout_mem1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.560 0.000 589.120 4.000 ;
    END
  END dout_mem1[15]
  PIN dout_mem1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 596.960 0.000 597.520 4.000 ;
    END
  END dout_mem1[16]
  PIN dout_mem1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 605.360 0.000 605.920 4.000 ;
    END
  END dout_mem1[17]
  PIN dout_mem1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 613.760 0.000 614.320 4.000 ;
    END
  END dout_mem1[18]
  PIN dout_mem1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 622.160 0.000 622.720 4.000 ;
    END
  END dout_mem1[19]
  PIN dout_mem1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.960 0.000 471.520 4.000 ;
    END
  END dout_mem1[1]
  PIN dout_mem1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 630.560 0.000 631.120 4.000 ;
    END
  END dout_mem1[20]
  PIN dout_mem1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 638.960 0.000 639.520 4.000 ;
    END
  END dout_mem1[21]
  PIN dout_mem1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 647.360 0.000 647.920 4.000 ;
    END
  END dout_mem1[22]
  PIN dout_mem1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 655.760 0.000 656.320 4.000 ;
    END
  END dout_mem1[23]
  PIN dout_mem1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 664.160 0.000 664.720 4.000 ;
    END
  END dout_mem1[24]
  PIN dout_mem1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.560 0.000 673.120 4.000 ;
    END
  END dout_mem1[25]
  PIN dout_mem1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 680.960 0.000 681.520 4.000 ;
    END
  END dout_mem1[26]
  PIN dout_mem1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 689.360 0.000 689.920 4.000 ;
    END
  END dout_mem1[27]
  PIN dout_mem1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 697.760 0.000 698.320 4.000 ;
    END
  END dout_mem1[28]
  PIN dout_mem1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 706.160 0.000 706.720 4.000 ;
    END
  END dout_mem1[29]
  PIN dout_mem1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 479.360 0.000 479.920 4.000 ;
    END
  END dout_mem1[2]
  PIN dout_mem1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 714.560 0.000 715.120 4.000 ;
    END
  END dout_mem1[30]
  PIN dout_mem1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 722.960 0.000 723.520 4.000 ;
    END
  END dout_mem1[31]
  PIN dout_mem1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.760 0.000 488.320 4.000 ;
    END
  END dout_mem1[3]
  PIN dout_mem1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 496.160 0.000 496.720 4.000 ;
    END
  END dout_mem1[4]
  PIN dout_mem1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.560 0.000 505.120 4.000 ;
    END
  END dout_mem1[5]
  PIN dout_mem1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 512.960 0.000 513.520 4.000 ;
    END
  END dout_mem1[6]
  PIN dout_mem1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 521.360 0.000 521.920 4.000 ;
    END
  END dout_mem1[7]
  PIN dout_mem1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 0.000 530.320 4.000 ;
    END
  END dout_mem1[8]
  PIN dout_mem1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 538.160 0.000 538.720 4.000 ;
    END
  END dout_mem1[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 97.970 15.380 99.570 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 282.070 15.380 283.670 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 466.170 15.380 467.770 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 650.270 15.380 651.870 184.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 190.020 15.380 191.620 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.120 15.380 375.720 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 558.220 15.380 559.820 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 742.320 15.380 743.920 184.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 743.920 184.540 ;
      LAYER Metal2 ;
        RECT 25.900 4.300 743.780 194.230 ;
        RECT 26.620 3.500 33.860 4.300 ;
        RECT 35.020 3.500 42.260 4.300 ;
        RECT 43.420 3.500 50.660 4.300 ;
        RECT 51.820 3.500 59.060 4.300 ;
        RECT 60.220 3.500 67.460 4.300 ;
        RECT 68.620 3.500 75.860 4.300 ;
        RECT 77.020 3.500 84.260 4.300 ;
        RECT 85.420 3.500 92.660 4.300 ;
        RECT 93.820 3.500 101.060 4.300 ;
        RECT 102.220 3.500 109.460 4.300 ;
        RECT 110.620 3.500 117.860 4.300 ;
        RECT 119.020 3.500 126.260 4.300 ;
        RECT 127.420 3.500 134.660 4.300 ;
        RECT 135.820 3.500 143.060 4.300 ;
        RECT 144.220 3.500 151.460 4.300 ;
        RECT 152.620 3.500 159.860 4.300 ;
        RECT 161.020 3.500 168.260 4.300 ;
        RECT 169.420 3.500 176.660 4.300 ;
        RECT 177.820 3.500 185.060 4.300 ;
        RECT 186.220 3.500 193.460 4.300 ;
        RECT 194.620 3.500 201.860 4.300 ;
        RECT 203.020 3.500 210.260 4.300 ;
        RECT 211.420 3.500 218.660 4.300 ;
        RECT 219.820 3.500 227.060 4.300 ;
        RECT 228.220 3.500 235.460 4.300 ;
        RECT 236.620 3.500 243.860 4.300 ;
        RECT 245.020 3.500 252.260 4.300 ;
        RECT 253.420 3.500 260.660 4.300 ;
        RECT 261.820 3.500 269.060 4.300 ;
        RECT 270.220 3.500 277.460 4.300 ;
        RECT 278.620 3.500 285.860 4.300 ;
        RECT 287.020 3.500 294.260 4.300 ;
        RECT 295.420 3.500 302.660 4.300 ;
        RECT 303.820 3.500 311.060 4.300 ;
        RECT 312.220 3.500 319.460 4.300 ;
        RECT 320.620 3.500 327.860 4.300 ;
        RECT 329.020 3.500 336.260 4.300 ;
        RECT 337.420 3.500 344.660 4.300 ;
        RECT 345.820 3.500 353.060 4.300 ;
        RECT 354.220 3.500 361.460 4.300 ;
        RECT 362.620 3.500 369.860 4.300 ;
        RECT 371.020 3.500 378.260 4.300 ;
        RECT 379.420 3.500 386.660 4.300 ;
        RECT 387.820 3.500 395.060 4.300 ;
        RECT 396.220 3.500 403.460 4.300 ;
        RECT 404.620 3.500 411.860 4.300 ;
        RECT 413.020 3.500 420.260 4.300 ;
        RECT 421.420 3.500 428.660 4.300 ;
        RECT 429.820 3.500 437.060 4.300 ;
        RECT 438.220 3.500 445.460 4.300 ;
        RECT 446.620 3.500 453.860 4.300 ;
        RECT 455.020 3.500 462.260 4.300 ;
        RECT 463.420 3.500 470.660 4.300 ;
        RECT 471.820 3.500 479.060 4.300 ;
        RECT 480.220 3.500 487.460 4.300 ;
        RECT 488.620 3.500 495.860 4.300 ;
        RECT 497.020 3.500 504.260 4.300 ;
        RECT 505.420 3.500 512.660 4.300 ;
        RECT 513.820 3.500 521.060 4.300 ;
        RECT 522.220 3.500 529.460 4.300 ;
        RECT 530.620 3.500 537.860 4.300 ;
        RECT 539.020 3.500 546.260 4.300 ;
        RECT 547.420 3.500 554.660 4.300 ;
        RECT 555.820 3.500 563.060 4.300 ;
        RECT 564.220 3.500 571.460 4.300 ;
        RECT 572.620 3.500 579.860 4.300 ;
        RECT 581.020 3.500 588.260 4.300 ;
        RECT 589.420 3.500 596.660 4.300 ;
        RECT 597.820 3.500 605.060 4.300 ;
        RECT 606.220 3.500 613.460 4.300 ;
        RECT 614.620 3.500 621.860 4.300 ;
        RECT 623.020 3.500 630.260 4.300 ;
        RECT 631.420 3.500 638.660 4.300 ;
        RECT 639.820 3.500 647.060 4.300 ;
        RECT 648.220 3.500 655.460 4.300 ;
        RECT 656.620 3.500 663.860 4.300 ;
        RECT 665.020 3.500 672.260 4.300 ;
        RECT 673.420 3.500 680.660 4.300 ;
        RECT 681.820 3.500 689.060 4.300 ;
        RECT 690.220 3.500 697.460 4.300 ;
        RECT 698.620 3.500 705.860 4.300 ;
        RECT 707.020 3.500 714.260 4.300 ;
        RECT 715.420 3.500 722.660 4.300 ;
        RECT 723.820 3.500 743.780 4.300 ;
      LAYER Metal3 ;
        RECT 25.850 193.460 745.700 194.180 ;
        RECT 25.850 190.140 746.000 193.460 ;
        RECT 25.850 188.980 745.700 190.140 ;
        RECT 25.850 185.660 746.000 188.980 ;
        RECT 25.850 184.500 745.700 185.660 ;
        RECT 25.850 181.180 746.000 184.500 ;
        RECT 25.850 180.020 745.700 181.180 ;
        RECT 25.850 176.700 746.000 180.020 ;
        RECT 25.850 175.540 745.700 176.700 ;
        RECT 25.850 172.220 746.000 175.540 ;
        RECT 25.850 171.060 745.700 172.220 ;
        RECT 25.850 167.740 746.000 171.060 ;
        RECT 25.850 166.580 745.700 167.740 ;
        RECT 25.850 163.260 746.000 166.580 ;
        RECT 25.850 162.100 745.700 163.260 ;
        RECT 25.850 158.780 746.000 162.100 ;
        RECT 25.850 157.620 745.700 158.780 ;
        RECT 25.850 154.300 746.000 157.620 ;
        RECT 25.850 153.140 745.700 154.300 ;
        RECT 25.850 149.820 746.000 153.140 ;
        RECT 25.850 148.660 745.700 149.820 ;
        RECT 25.850 145.340 746.000 148.660 ;
        RECT 25.850 144.180 745.700 145.340 ;
        RECT 25.850 140.860 746.000 144.180 ;
        RECT 25.850 139.700 745.700 140.860 ;
        RECT 25.850 136.380 746.000 139.700 ;
        RECT 25.850 135.220 745.700 136.380 ;
        RECT 25.850 131.900 746.000 135.220 ;
        RECT 25.850 130.740 745.700 131.900 ;
        RECT 25.850 127.420 746.000 130.740 ;
        RECT 25.850 126.260 745.700 127.420 ;
        RECT 25.850 122.940 746.000 126.260 ;
        RECT 25.850 121.780 745.700 122.940 ;
        RECT 25.850 118.460 746.000 121.780 ;
        RECT 25.850 117.300 745.700 118.460 ;
        RECT 25.850 113.980 746.000 117.300 ;
        RECT 25.850 112.820 745.700 113.980 ;
        RECT 25.850 109.500 746.000 112.820 ;
        RECT 25.850 108.340 745.700 109.500 ;
        RECT 25.850 105.020 746.000 108.340 ;
        RECT 25.850 103.860 745.700 105.020 ;
        RECT 25.850 100.540 746.000 103.860 ;
        RECT 25.850 99.380 745.700 100.540 ;
        RECT 25.850 96.060 746.000 99.380 ;
        RECT 25.850 94.900 745.700 96.060 ;
        RECT 25.850 91.580 746.000 94.900 ;
        RECT 25.850 90.420 745.700 91.580 ;
        RECT 25.850 87.100 746.000 90.420 ;
        RECT 25.850 85.940 745.700 87.100 ;
        RECT 25.850 82.620 746.000 85.940 ;
        RECT 25.850 81.460 745.700 82.620 ;
        RECT 25.850 78.140 746.000 81.460 ;
        RECT 25.850 76.980 745.700 78.140 ;
        RECT 25.850 73.660 746.000 76.980 ;
        RECT 25.850 72.500 745.700 73.660 ;
        RECT 25.850 69.180 746.000 72.500 ;
        RECT 25.850 68.020 745.700 69.180 ;
        RECT 25.850 64.700 746.000 68.020 ;
        RECT 25.850 63.540 745.700 64.700 ;
        RECT 25.850 60.220 746.000 63.540 ;
        RECT 25.850 59.060 745.700 60.220 ;
        RECT 25.850 55.740 746.000 59.060 ;
        RECT 25.850 54.580 745.700 55.740 ;
        RECT 25.850 51.260 746.000 54.580 ;
        RECT 25.850 50.100 745.700 51.260 ;
        RECT 25.850 46.780 746.000 50.100 ;
        RECT 25.850 45.620 745.700 46.780 ;
        RECT 25.850 42.300 746.000 45.620 ;
        RECT 25.850 41.140 745.700 42.300 ;
        RECT 25.850 37.820 746.000 41.140 ;
        RECT 25.850 36.660 745.700 37.820 ;
        RECT 25.850 33.340 746.000 36.660 ;
        RECT 25.850 32.180 745.700 33.340 ;
        RECT 25.850 28.860 746.000 32.180 ;
        RECT 25.850 27.700 745.700 28.860 ;
        RECT 25.850 24.380 746.000 27.700 ;
        RECT 25.850 23.220 745.700 24.380 ;
        RECT 25.850 19.900 746.000 23.220 ;
        RECT 25.850 18.740 745.700 19.900 ;
        RECT 25.850 15.420 746.000 18.740 ;
        RECT 25.850 14.260 745.700 15.420 ;
        RECT 25.850 10.940 746.000 14.260 ;
        RECT 25.850 9.780 745.700 10.940 ;
        RECT 25.850 6.460 746.000 9.780 ;
        RECT 25.850 5.300 745.700 6.460 ;
        RECT 25.850 4.060 746.000 5.300 ;
      LAYER Metal4 ;
        RECT 152.460 16.890 189.720 30.150 ;
        RECT 191.920 16.890 281.770 30.150 ;
        RECT 283.970 16.890 373.820 30.150 ;
        RECT 376.020 16.890 465.870 30.150 ;
        RECT 468.070 16.890 557.920 30.150 ;
        RECT 560.120 16.890 649.970 30.150 ;
        RECT 652.170 16.890 655.060 30.150 ;
  END
END merge_memory
END LIBRARY

