* NGSPICE file created from wb_mux.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

.subckt wb_mux io_wbs_ack io_wbs_ack_0 io_wbs_ack_1 io_wbs_adr[0] io_wbs_adr[10] io_wbs_adr[11]
+ io_wbs_adr[12] io_wbs_adr[13] io_wbs_adr[14] io_wbs_adr[15] io_wbs_adr[16] io_wbs_adr[17]
+ io_wbs_adr[18] io_wbs_adr[19] io_wbs_adr[1] io_wbs_adr[20] io_wbs_adr[21] io_wbs_adr[22]
+ io_wbs_adr[23] io_wbs_adr[24] io_wbs_adr[25] io_wbs_adr[26] io_wbs_adr[27] io_wbs_adr[28]
+ io_wbs_adr[29] io_wbs_adr[2] io_wbs_adr[30] io_wbs_adr[31] io_wbs_adr[3] io_wbs_adr[4]
+ io_wbs_adr[5] io_wbs_adr[6] io_wbs_adr[7] io_wbs_adr[8] io_wbs_adr[9] io_wbs_adr_0[0]
+ io_wbs_adr_0[10] io_wbs_adr_0[11] io_wbs_adr_0[12] io_wbs_adr_0[13] io_wbs_adr_0[14]
+ io_wbs_adr_0[15] io_wbs_adr_0[16] io_wbs_adr_0[17] io_wbs_adr_0[18] io_wbs_adr_0[19]
+ io_wbs_adr_0[1] io_wbs_adr_0[20] io_wbs_adr_0[21] io_wbs_adr_0[22] io_wbs_adr_0[23]
+ io_wbs_adr_0[24] io_wbs_adr_0[25] io_wbs_adr_0[26] io_wbs_adr_0[27] io_wbs_adr_0[28]
+ io_wbs_adr_0[29] io_wbs_adr_0[2] io_wbs_adr_0[30] io_wbs_adr_0[31] io_wbs_adr_0[3]
+ io_wbs_adr_0[4] io_wbs_adr_0[5] io_wbs_adr_0[6] io_wbs_adr_0[7] io_wbs_adr_0[8]
+ io_wbs_adr_0[9] io_wbs_adr_1[0] io_wbs_adr_1[10] io_wbs_adr_1[11] io_wbs_adr_1[12]
+ io_wbs_adr_1[13] io_wbs_adr_1[14] io_wbs_adr_1[15] io_wbs_adr_1[16] io_wbs_adr_1[17]
+ io_wbs_adr_1[18] io_wbs_adr_1[19] io_wbs_adr_1[1] io_wbs_adr_1[20] io_wbs_adr_1[21]
+ io_wbs_adr_1[22] io_wbs_adr_1[23] io_wbs_adr_1[24] io_wbs_adr_1[25] io_wbs_adr_1[26]
+ io_wbs_adr_1[27] io_wbs_adr_1[28] io_wbs_adr_1[29] io_wbs_adr_1[2] io_wbs_adr_1[30]
+ io_wbs_adr_1[31] io_wbs_adr_1[3] io_wbs_adr_1[4] io_wbs_adr_1[5] io_wbs_adr_1[6]
+ io_wbs_adr_1[7] io_wbs_adr_1[8] io_wbs_adr_1[9] io_wbs_cyc io_wbs_cyc_0 io_wbs_cyc_1
+ io_wbs_datrd[0] io_wbs_datrd[10] io_wbs_datrd[11] io_wbs_datrd[12] io_wbs_datrd[13]
+ io_wbs_datrd[14] io_wbs_datrd[15] io_wbs_datrd[16] io_wbs_datrd[17] io_wbs_datrd[18]
+ io_wbs_datrd[19] io_wbs_datrd[1] io_wbs_datrd[20] io_wbs_datrd[21] io_wbs_datrd[22]
+ io_wbs_datrd[23] io_wbs_datrd[24] io_wbs_datrd[25] io_wbs_datrd[26] io_wbs_datrd[27]
+ io_wbs_datrd[28] io_wbs_datrd[29] io_wbs_datrd[2] io_wbs_datrd[30] io_wbs_datrd[31]
+ io_wbs_datrd[3] io_wbs_datrd[4] io_wbs_datrd[5] io_wbs_datrd[6] io_wbs_datrd[7]
+ io_wbs_datrd[8] io_wbs_datrd[9] io_wbs_datrd_0[0] io_wbs_datrd_0[10] io_wbs_datrd_0[11]
+ io_wbs_datrd_0[12] io_wbs_datrd_0[13] io_wbs_datrd_0[14] io_wbs_datrd_0[15] io_wbs_datrd_0[16]
+ io_wbs_datrd_0[17] io_wbs_datrd_0[18] io_wbs_datrd_0[19] io_wbs_datrd_0[1] io_wbs_datrd_0[20]
+ io_wbs_datrd_0[21] io_wbs_datrd_0[22] io_wbs_datrd_0[23] io_wbs_datrd_0[24] io_wbs_datrd_0[25]
+ io_wbs_datrd_0[26] io_wbs_datrd_0[27] io_wbs_datrd_0[28] io_wbs_datrd_0[29] io_wbs_datrd_0[2]
+ io_wbs_datrd_0[30] io_wbs_datrd_0[31] io_wbs_datrd_0[3] io_wbs_datrd_0[4] io_wbs_datrd_0[5]
+ io_wbs_datrd_0[6] io_wbs_datrd_0[7] io_wbs_datrd_0[8] io_wbs_datrd_0[9] io_wbs_datrd_1[0]
+ io_wbs_datrd_1[10] io_wbs_datrd_1[11] io_wbs_datrd_1[12] io_wbs_datrd_1[13] io_wbs_datrd_1[14]
+ io_wbs_datrd_1[15] io_wbs_datrd_1[16] io_wbs_datrd_1[17] io_wbs_datrd_1[18] io_wbs_datrd_1[19]
+ io_wbs_datrd_1[1] io_wbs_datrd_1[20] io_wbs_datrd_1[21] io_wbs_datrd_1[22] io_wbs_datrd_1[23]
+ io_wbs_datrd_1[24] io_wbs_datrd_1[25] io_wbs_datrd_1[26] io_wbs_datrd_1[27] io_wbs_datrd_1[28]
+ io_wbs_datrd_1[29] io_wbs_datrd_1[2] io_wbs_datrd_1[30] io_wbs_datrd_1[31] io_wbs_datrd_1[3]
+ io_wbs_datrd_1[4] io_wbs_datrd_1[5] io_wbs_datrd_1[6] io_wbs_datrd_1[7] io_wbs_datrd_1[8]
+ io_wbs_datrd_1[9] io_wbs_datwr[0] io_wbs_datwr[10] io_wbs_datwr[11] io_wbs_datwr[12]
+ io_wbs_datwr[13] io_wbs_datwr[14] io_wbs_datwr[15] io_wbs_datwr[16] io_wbs_datwr[17]
+ io_wbs_datwr[18] io_wbs_datwr[19] io_wbs_datwr[1] io_wbs_datwr[20] io_wbs_datwr[21]
+ io_wbs_datwr[22] io_wbs_datwr[23] io_wbs_datwr[24] io_wbs_datwr[25] io_wbs_datwr[26]
+ io_wbs_datwr[27] io_wbs_datwr[28] io_wbs_datwr[29] io_wbs_datwr[2] io_wbs_datwr[30]
+ io_wbs_datwr[31] io_wbs_datwr[3] io_wbs_datwr[4] io_wbs_datwr[5] io_wbs_datwr[6]
+ io_wbs_datwr[7] io_wbs_datwr[8] io_wbs_datwr[9] io_wbs_datwr_0[0] io_wbs_datwr_0[10]
+ io_wbs_datwr_0[11] io_wbs_datwr_0[12] io_wbs_datwr_0[13] io_wbs_datwr_0[14] io_wbs_datwr_0[15]
+ io_wbs_datwr_0[16] io_wbs_datwr_0[17] io_wbs_datwr_0[18] io_wbs_datwr_0[19] io_wbs_datwr_0[1]
+ io_wbs_datwr_0[20] io_wbs_datwr_0[21] io_wbs_datwr_0[22] io_wbs_datwr_0[23] io_wbs_datwr_0[24]
+ io_wbs_datwr_0[25] io_wbs_datwr_0[26] io_wbs_datwr_0[27] io_wbs_datwr_0[28] io_wbs_datwr_0[29]
+ io_wbs_datwr_0[2] io_wbs_datwr_0[30] io_wbs_datwr_0[31] io_wbs_datwr_0[3] io_wbs_datwr_0[4]
+ io_wbs_datwr_0[5] io_wbs_datwr_0[6] io_wbs_datwr_0[7] io_wbs_datwr_0[8] io_wbs_datwr_0[9]
+ io_wbs_datwr_1[0] io_wbs_datwr_1[10] io_wbs_datwr_1[11] io_wbs_datwr_1[12] io_wbs_datwr_1[13]
+ io_wbs_datwr_1[14] io_wbs_datwr_1[15] io_wbs_datwr_1[16] io_wbs_datwr_1[17] io_wbs_datwr_1[18]
+ io_wbs_datwr_1[19] io_wbs_datwr_1[1] io_wbs_datwr_1[20] io_wbs_datwr_1[21] io_wbs_datwr_1[22]
+ io_wbs_datwr_1[23] io_wbs_datwr_1[24] io_wbs_datwr_1[25] io_wbs_datwr_1[26] io_wbs_datwr_1[27]
+ io_wbs_datwr_1[28] io_wbs_datwr_1[29] io_wbs_datwr_1[2] io_wbs_datwr_1[30] io_wbs_datwr_1[31]
+ io_wbs_datwr_1[3] io_wbs_datwr_1[4] io_wbs_datwr_1[5] io_wbs_datwr_1[6] io_wbs_datwr_1[7]
+ io_wbs_datwr_1[8] io_wbs_datwr_1[9] io_wbs_sel[0] io_wbs_sel[1] io_wbs_sel[2] io_wbs_sel[3]
+ io_wbs_sel_0[0] io_wbs_sel_0[1] io_wbs_sel_0[2] io_wbs_sel_0[3] io_wbs_sel_1[0]
+ io_wbs_sel_1[1] io_wbs_sel_1[2] io_wbs_sel_1[3] io_wbs_stb io_wbs_stb_0 io_wbs_stb_1
+ io_wbs_we io_wbs_we_0 io_wbs_we_1 vdd vss
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input108_I io_wbs_datwr[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__254__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input73_I io_wbs_datrd_1[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__105__A4 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_363_ net123 net292 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_294_ net20 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__164__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__339__I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__249__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output277_I net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_346_ net104 net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_277_ net33 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput220 net220 io_wbs_datrd[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput231 net231 io_wbs_datrd[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput242 net242 io_wbs_datwr_0[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput253 net253 io_wbs_datwr_0[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput264 net264 io_wbs_datwr_0[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput275 net275 io_wbs_datwr_1[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput286 net286 io_wbs_datwr_1[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput297 net297 io_wbs_datwr_1[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input36_I io_wbs_datrd_0[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_200_ net50 _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_131_ _026_ _022_ _024_ _027_ net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_3_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_329_ net120 net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__352__I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__262__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output142_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_114_ _013_ _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__172__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__347__I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__257__I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__108__A2 _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput120 io_wbs_datwr[28] net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput131 io_wbs_datwr[9] net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__360__I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input66_I io_wbs_datrd_0[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output222_I net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_362_ net121 net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_293_ net19 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__180__I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__355__I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input120_I io_wbs_datwr[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__265__I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output172_I net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__175__I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_345_ net103 net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_276_ net32 net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput210 net210 io_wbs_datrd[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput232 net232 io_wbs_datrd[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput221 net221 io_wbs_datrd[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput243 net243 io_wbs_datwr_0[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput265 net265 io_wbs_datwr_0[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput276 net276 io_wbs_datwr_1[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput254 net254 io_wbs_datwr_0[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput298 net298 io_wbs_datwr_1[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput287 net287 io_wbs_datwr_1[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input29_I io_wbs_adr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_130_ net58 _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_328_ net119 net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_259_ net17 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_113_ _012_ _003_ _006_ _007_ _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__363__I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input96_I io_wbs_datrd_1[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output252_I net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__183__I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__358__I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I io_wbs_adr[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__268__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__108__A3 _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput110 io_wbs_datwr[19] net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput132 io_wbs_sel[0] net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput121 io_wbs_datwr[29] net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__178__I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input3_I io_wbs_adr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input59_I io_wbs_datrd_0[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output215_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_361_ net120 net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_292_ net18 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__371__I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input113_I io_wbs_datwr[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__281__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output165_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_344_ net102 net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_275_ net31 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__191__I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__366__I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput200 net200 io_wbs_adr_1[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput222 net222 io_wbs_datrd[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput233 net233 io_wbs_datrd[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput211 net211 io_wbs_datrd[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput244 net244 io_wbs_datwr_0[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput266 net266 io_wbs_datwr_0[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput277 net277 io_wbs_datwr_1[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput255 net255 io_wbs_datwr_0[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_58_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput299 net299 io_wbs_datwr_1[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput288 net288 io_wbs_datwr_1[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output282_I net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__186__I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_327_ net118 net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_258_ net16 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_189_ net46 _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input41_I io_wbs_datrd_0[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_112_ net6 _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input89_I io_wbs_datrd_1[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output245_I net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__374__I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__284__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output195_I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput100 io_wbs_datwr[0] net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput111 io_wbs_datwr[1] net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput133 io_wbs_sel[1] net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput122 io_wbs_datwr[2] net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__194__I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__369__I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__279__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output208_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_360_ net119 net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_291_ net17 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__189__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input106_I io_wbs_datwr[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input71_I io_wbs_datrd_1[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output158_I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_343_ net101 net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_274_ net30 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput201 net201 io_wbs_adr_1[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput212 net212 io_wbs_datrd[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput223 net223 io_wbs_datrd[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput234 net234 io_wbs_datrd[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput267 net267 io_wbs_datwr_0[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput245 net245 io_wbs_datwr_0[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput256 net256 io_wbs_datwr_0[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput278 net278 io_wbs_datwr_1[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput289 net289 io_wbs_datwr_1[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_74_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__292__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output275_I net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_326_ net117 net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_257_ net15 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_188_ net78 _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input34_I io_wbs_adr[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__287__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_111_ _010_ _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__197__I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_309_ net130 net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output140_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output238_I net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input136_I io_wbs_stb vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output188_I net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput101 io_wbs_datwr[10] net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput123 io_wbs_datwr[30] net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput134 io_wbs_sel[2] net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput112 io_wbs_datwr[20] net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__295__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_290_ net16 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input64_I io_wbs_datrd_0[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output220_I net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_342_ net131 net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_273_ net29 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput202 net202 io_wbs_adr_1[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput224 net224 io_wbs_datrd[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput235 net235 io_wbs_datrd[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput213 net213 io_wbs_datrd[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput268 net268 io_wbs_datwr_0[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput246 net246 io_wbs_datwr_0[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput257 net257 io_wbs_datwr_0[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput279 net279 io_wbs_datwr_1[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output170_I net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output268_I net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_325_ net116 net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_256_ net13 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_187_ _066_ _063_ _064_ _067_ net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input27_I io_wbs_adr[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_110_ _009_ _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_308_ net129 net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_239_ net25 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__298__I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output300_I net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input129_I io_wbs_datwr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input94_I io_wbs_datrd_1[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output250_I net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput102 io_wbs_datwr[11] net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput113 io_wbs_datwr[21] net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput124 io_wbs_datwr[31] net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput135 io_wbs_sel[3] net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_56_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output298_I net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input1_I io_wbs_ack_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input57_I io_wbs_datrd_0[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__101__A1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output213_I net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_341_ net130 net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_272_ net28 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput203 net203 io_wbs_cyc_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput225 net225 io_wbs_datrd[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput214 net214 io_wbs_datrd[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput236 net236 io_wbs_datrd[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput247 net247 io_wbs_datwr_0[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput258 net258 io_wbs_datwr_0[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput269 net269 io_wbs_datwr_1[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input111_I io_wbs_datwr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output163_I net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_324_ net115 net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_255_ net12 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_186_ net45 _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output280_I net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_307_ net128 net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_238_ net14 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_169_ net40 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input87_I io_wbs_datrd_1[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput103 io_wbs_datwr[12] net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput136 io_wbs_stb net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput125 io_wbs_datwr[3] net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput114 io_wbs_datwr[22] net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_output243_I net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__101__A2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output206_I net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_340_ net129 net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_271_ net25 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput204 net204 io_wbs_cyc_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput226 net226 io_wbs_datrd[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput215 net215 io_wbs_datrd[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput248 net248 io_wbs_datwr_0[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput237 net237 io_wbs_datwr_0[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput259 net259 io_wbs_datwr_0[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__200__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input104_I io_wbs_datwr[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output156_I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__110__I _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_323_ net114 net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_254_ net11 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_185_ net77 _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output273_I net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_306_ net127 net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_237_ net3 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_168_ _023_ _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input32_I io_wbs_adr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput126 io_wbs_datwr[4] net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput104 io_wbs_datwr[13] net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput115 io_wbs_datwr[23] net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_output236_I net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput137 io_wbs_we net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__203__I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input134_I io_wbs_sel[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output186_I net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__101__A3 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_270_ net14 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput216 net216 io_wbs_datrd[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput205 net205 io_wbs_datrd[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput227 net227 io_wbs_datrd[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput238 net238 io_wbs_datwr_0[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput249 net249 io_wbs_datwr_0[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input62_I io_wbs_datrd_0[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output149_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_322_ net113 net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_253_ net10 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_184_ _062_ _063_ _064_ _065_ net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__301__I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__211__I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output266_I net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_305_ net126 net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_236_ _099_ _011_ net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_167_ _021_ _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__206__I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input25_I io_wbs_adr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_219_ net88 _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput127 io_wbs_datwr[5] net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput105 io_wbs_datwr[14] net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput116 io_wbs_datwr[24] net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output229_I net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input127_I io_wbs_datwr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input92_I io_wbs_datrd_1[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output179_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__104__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__304__I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__214__I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__101__A4 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output296_I net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput217 net217 io_wbs_datrd[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput206 net206 io_wbs_datrd[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput228 net228 io_wbs_datrd[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput239 net239 io_wbs_datwr_0[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_4_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__209__I _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input55_I io_wbs_datrd_0[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output211_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_321_ net112 net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__119__I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_252_ net9 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_183_ net44 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output161_I net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output259_I net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_304_ net125 net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_235_ _098_ _011_ net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_166_ net72 _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__312__I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__222__I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input18_I io_wbs_adr[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__132__I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__307__I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_218_ _088_ _083_ _084_ _089_ net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_149_ net98 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__217__I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput106 io_wbs_datwr[15] net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput117 io_wbs_datwr[25] net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput128 io_wbs_datwr[6] net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__127__I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__113__A2 _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input85_I io_wbs_datrd_1[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__104__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output241_I net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__320__I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output191_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output289_I net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__140__I _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__315__I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput207 net207 io_wbs_datrd[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput229 net229 io_wbs_datrd[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput218 net218 io_wbs_datrd[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__225__I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input48_I io_wbs_datrd_0[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output204_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_320_ net110 net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_251_ net8 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_182_ _014_ _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__135__I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input102_I io_wbs_datwr[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output154_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_303_ net122 net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_234_ _099_ _016_ net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_165_ _050_ _043_ _044_ _051_ net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_2_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output271_I net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_217_ net55 _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_148_ _038_ _033_ _034_ _039_ net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__323__I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__233__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput107 io_wbs_datwr[16] net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput118 io_wbs_datwr[26] net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput129 io_wbs_datwr[7] net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input30_I io_wbs_adr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__143__I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__318__I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__113__A3 _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__228__I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input78_I io_wbs_datrd_1[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__104__A3 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output234_I net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__138__I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input132_I io_wbs_sel[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output184_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput208 net208 io_wbs_datrd[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput219 net219 io_wbs_datrd[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__331__I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_250_ net7 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_181_ _009_ _063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__234__A2 _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__326__I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input60_I io_wbs_datrd_0[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output147_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_302_ net111 net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_233_ net35 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__146__I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_164_ net39 _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output264_I net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_216_ net87 _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_147_ net65 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput108 io_wbs_datwr[17] net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput119 io_wbs_datwr[27] net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input23_I io_wbs_adr[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__107__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__334__I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput90 io_wbs_datrd_1[2] net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__104__A4 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output227_I net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__154__I _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__329__I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input125_I io_wbs_datwr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input90_I io_wbs_datrd_1[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output177_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__149__I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput209 net209 io_wbs_datrd[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_4_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output294_I net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_180_ net76 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__342__I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__252__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input53_I io_wbs_datrd_0[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output307_I net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_301_ net100 net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_232_ _098_ _016_ net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_163_ net71 _050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__337__I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__247__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output257_I net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__157__I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_215_ _086_ _083_ _084_ _087_ net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_146_ net97 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput109 io_wbs_datwr[18] net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_69_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input16_I io_wbs_adr[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__107__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_129_ net90 _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__350__I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I io_wbs_adr[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput80 io_wbs_datrd_1[20] net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput91 io_wbs_datrd_1[30] net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__260__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__345__I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input118_I io_wbs_datwr[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__255__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input83_I io_wbs_datrd_1[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output287_I net287 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input46_I io_wbs_datrd_0[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_300_ net27 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_231_ net136 _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_162_ _048_ _043_ _044_ _049_ net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__353__I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 io_wbs_ack_0 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input100_I io_wbs_datwr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__263__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output152_I net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_214_ net54 _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_145_ _036_ _033_ _034_ _037_ net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__348__I net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__258__I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__107__A3 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput190 net190 io_wbs_adr_1[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__168__I _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_128_ _020_ _022_ _024_ _025_ net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput70 io_wbs_datrd_1[11] net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput81 io_wbs_datrd_1[21] net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput92 io_wbs_datrd_1[31] net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__361__I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input76_I io_wbs_datrd_1[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output232_I net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__181__I _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__356__I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input130_I io_wbs_datwr[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__266__I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input39_I io_wbs_datrd_0[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_230_ _096_ _010_ _015_ _097_ net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_50_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_161_ net38 _049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_359_ net118 net287 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 io_wbs_ack_1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output145_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output312_I net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_213_ net86 _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_144_ net64 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__364__I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output262_I net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput180 net180 io_wbs_adr_1[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput191 net191 io_wbs_adr_1[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_127_ net47 _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__359__I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput71 io_wbs_datrd_1[12] net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput82 io_wbs_datrd_1[22] net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput60 io_wbs_datrd_0[31] net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput93 io_wbs_datrd_1[3] net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input21_I io_wbs_adr[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input69_I io_wbs_datrd_1[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output225_I net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__372__I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input123_I io_wbs_datwr[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__282__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output175_I net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__192__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__367__I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output292_I net292 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_160_ net70 _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_358_ net117 net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_289_ net15 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput3 io_wbs_adr[0] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input51_I io_wbs_datrd_0[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output138_I net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output305_I net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_212_ _082_ _083_ _084_ _085_ net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_51_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_143_ net96 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input99_I io_wbs_datrd_1[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__290__I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput170 net170 io_wbs_adr_0[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output255_I net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput181 net181 io_wbs_adr_1[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput192 net192 io_wbs_adr_1[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_126_ _023_ _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput61 io_wbs_datrd_0[3] net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput72 io_wbs_datrd_1[13] net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput50 io_wbs_datrd_0[22] net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput94 io_wbs_datrd_1[4] net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput83 io_wbs_datrd_1[23] net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input14_I io_wbs_adr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__285__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__195__I _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_109_ _008_ _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_wbs_adr[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output218_I net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input116_I io_wbs_datwr[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input81_I io_wbs_datrd_1[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output168_I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_374_ net137 net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__293__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output285_I net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_357_ net116 net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_288_ net13 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_wbs_adr[10] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input44_I io_wbs_datrd_0[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__288__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_211_ net53 _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_142_ _032_ _033_ _034_ _035_ net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_2_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput160 net160 io_wbs_adr_0[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput193 net193 io_wbs_adr_1[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output150_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput182 net182 io_wbs_adr_1[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput171 net171 io_wbs_adr_1[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output248_I net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_125_ _013_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput40 io_wbs_datrd_0[13] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput62 io_wbs_datrd_0[4] net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput73 io_wbs_datrd_1[14] net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput51 io_wbs_datrd_0[23] net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput95 io_wbs_datrd_1[5] net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput84 io_wbs_datrd_1[24] net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_108_ net6 _003_ _006_ _007_ _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__296__I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input109_I io_wbs_datwr[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input74_I io_wbs_datrd_1[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output230_I net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_373_ net137 net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output180_I net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output278_I net278 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_356_ net115 net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_287_ net12 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 io_wbs_adr[11] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input37_I io_wbs_datrd_0[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_210_ _014_ _084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_141_ net63 _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_339_ net128 net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput161 net161 io_wbs_adr_0[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput150 net150 io_wbs_adr_0[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput172 net172 io_wbs_adr_1[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput183 net183 io_wbs_adr_1[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput194 net194 io_wbs_adr_1[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__299__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output143_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output310_I net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_124_ _021_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput30 io_wbs_adr[5] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_30_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput63 io_wbs_datrd_0[5] net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput41 io_wbs_datrd_0[14] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput52 io_wbs_datrd_0[24] net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput96 io_wbs_datrd_1[6] net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput74 io_wbs_datrd_1[15] net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput85 io_wbs_datrd_1[25] net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output260_I net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_107_ net9 net8 net7 _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input67_I io_wbs_datrd_0[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output223_I net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__100__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_372_ net135 net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input121_I io_wbs_datwr[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output173_I net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_355_ net114 net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_286_ net11 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput6 io_wbs_adr[12] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput310 net310 io_wbs_stb_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_140_ _023_ _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output290_I net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_338_ net127 net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_269_ net3 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput140 net140 io_wbs_adr_0[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput151 net151 io_wbs_adr_0[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput173 net173 io_wbs_adr_1[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput184 net184 io_wbs_adr_1[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput195 net195 io_wbs_adr_1[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput162 net162 io_wbs_adr_0[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_123_ _008_ _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__121__B1 _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput20 io_wbs_adr[25] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput31 io_wbs_adr[6] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput64 io_wbs_datrd_0[6] net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput42 io_wbs_datrd_0[15] net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput53 io_wbs_datrd_0[25] net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput97 io_wbs_datrd_1[7] net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput75 io_wbs_datrd_1[16] net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput86 io_wbs_datrd_1[26] net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input97_I io_wbs_datrd_1[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output253_I net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_106_ _004_ _005_ _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I io_wbs_adr[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I io_wbs_adr[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output216_I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_371_ net134 net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input114_I io_wbs_datwr[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output166_I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_354_ net113 net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_285_ net10 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput7 io_wbs_adr[13] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput300 net300 io_wbs_datwr_1[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput311 net311 io_wbs_we_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output283_I net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_337_ net126 net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_268_ net27 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_199_ net82 _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput141 net141 io_wbs_adr_0[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput152 net152 io_wbs_adr_0[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput174 net174 io_wbs_adr_1[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput185 net185 io_wbs_adr_1[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput163 net163 io_wbs_adr_0[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input42_I io_wbs_datrd_0[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput196 net196 io_wbs_adr_1[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_122_ net79 _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput21 io_wbs_adr[26] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput10 io_wbs_adr[16] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput32 io_wbs_adr[7] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput43 io_wbs_datrd_0[16] net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput54 io_wbs_datrd_0[26] net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput65 io_wbs_datrd_0[7] net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput98 io_wbs_datrd_1[8] net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput76 io_wbs_datrd_1[17] net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput87 io_wbs_datrd_1[27] net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__103__A1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output246_I net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_105_ net20 net19 net22 net21 _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__114__I _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output209_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_370_ net133 net306 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__109__I _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input107_I io_wbs_datwr[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input72_I io_wbs_datrd_1[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output159_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_353_ net112 net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_284_ net9 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__302__I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput8 io_wbs_adr[14] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput301 net301 io_wbs_sel_0[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput312 net312 io_wbs_we_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_28_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output276_I net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__122__I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_336_ net125 net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_267_ net26 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_198_ _072_ _073_ _074_ _075_ net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_2_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput142 net142 io_wbs_adr_0[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput175 net175 io_wbs_adr_1[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput164 net164 io_wbs_adr_0[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput153 net153 io_wbs_adr_0[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput186 net186 io_wbs_adr_1[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput197 net197 io_wbs_adr_1[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input35_I io_wbs_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_121_ _018_ _011_ _016_ _019_ net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__117__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__121__A2 _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 io_wbs_adr[17] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput22 io_wbs_adr[27] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_319_ net109 net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput33 io_wbs_adr[8] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput44 io_wbs_datrd_0[17] net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput55 io_wbs_datrd_0[27] net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput66 io_wbs_datrd_0[8] net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput77 io_wbs_datrd_1[18] net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput88 io_wbs_datrd_1[28] net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput99 io_wbs_datrd_1[9] net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__103__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output141_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output239_I net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_104_ net11 net10 net13 net12 _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_3_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__310__I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__220__I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input137_I io_wbs_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output189_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__130__I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__305__I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__125__I _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input65_I io_wbs_datrd_0[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output221_I net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_352_ net110 net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_283_ net8 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 io_wbs_adr[15] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput302 net302 io_wbs_sel_0[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_19_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output269_I net269 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_335_ net122 net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_266_ net24 net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_197_ net49 _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__313__I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput143 net143 io_wbs_adr_0[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput176 net176 io_wbs_adr_1[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput165 net165 io_wbs_adr_0[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput154 net154 io_wbs_adr_0[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput198 net198 io_wbs_adr_1[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput187 net187 io_wbs_adr_1[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input28_I io_wbs_adr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_120_ net36 _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__133__I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__308__I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput12 io_wbs_adr[18] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_318_ net108 net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_249_ net6 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput34 io_wbs_adr[9] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput23 io_wbs_adr[28] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput45 io_wbs_datrd_0[18] net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput67 io_wbs_datrd_0[9] net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput78 io_wbs_datrd_1[19] net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput56 io_wbs_datrd_0[28] net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput89 io_wbs_datrd_1[29] net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_103_ net24 net23 _001_ _002_ _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input95_I io_wbs_datrd_1[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output251_I net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__321__I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__231__I net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input10_I io_wbs_adr[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output299_I net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__141__I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__316__I net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I io_wbs_ack_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input58_I io_wbs_datrd_0[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output214_I net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_351_ net109 net278 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_282_ net7 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__136__I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput303 net303 io_wbs_sel_0[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input112_I io_wbs_datwr[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output164_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_334_ net111 net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_265_ net23 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_196_ _014_ _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput144 net144 io_wbs_adr_0[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput177 net177 io_wbs_adr_1[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput166 net166 io_wbs_adr_0[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput155 net155 io_wbs_adr_0[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput199 net199 io_wbs_adr_1[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput188 net188 io_wbs_adr_1[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_83_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output281_I net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_317_ net107 net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput13 io_wbs_adr[19] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_248_ net5 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput24 io_wbs_adr[29] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput35 io_wbs_cyc net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__324__I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput46 io_wbs_datrd_0[19] net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput68 io_wbs_datrd_1[0] net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput79 io_wbs_datrd_1[1] net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_179_ _060_ _053_ _054_ _061_ net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xinput57 io_wbs_datrd_0[29] net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input40_I io_wbs_datrd_0[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_102_ net27 net26 _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__144__I net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__319__I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input88_I io_wbs_datrd_1[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output244_I net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output194_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__332__I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output207_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_350_ net108 net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_281_ net6 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__152__I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__327__I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput304 net304 io_wbs_sel_0[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input105_I io_wbs_datwr[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input70_I io_wbs_datrd_1[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output157_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__147__I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_333_ net100 net269 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_264_ net22 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_195_ _009_ _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput145 net145 io_wbs_adr_0[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput167 net167 io_wbs_adr_0[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput156 net156 io_wbs_adr_0[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput178 net178 io_wbs_adr_1[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput189 net189 io_wbs_adr_1[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_46_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output274_I net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_316_ net106 net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_247_ net4 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 io_wbs_adr[2] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput14 io_wbs_adr[1] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput36 io_wbs_datrd_0[0] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput47 io_wbs_datrd_0[1] net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput58 io_wbs_datrd_0[2] net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput69 io_wbs_datrd_1[10] net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_178_ net43 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__340__I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__250__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input33_I io_wbs_adr[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_101_ net16 net15 net18 net17 _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_3_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__160__I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__335__I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output237_I net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__155__I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input135_I io_wbs_sel[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output187_I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_280_ net5 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__343__I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput305 net305 io_wbs_sel_1[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_55_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__253__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__118__B1 _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input63_I io_wbs_datrd_0[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_332_ net124 net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_263_ net21 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__163__I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_194_ net81 _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__338__I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput146 net146 io_wbs_adr_0[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput168 net168 io_wbs_adr_0[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput157 net157 io_wbs_adr_0[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput179 net179 io_wbs_adr_1[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_46_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__248__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output267_I net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__158__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_315_ net105 net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_246_ net34 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 io_wbs_adr[30] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput15 io_wbs_adr[20] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput37 io_wbs_datrd_0[10] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_177_ net75 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput48 io_wbs_datrd_0[20] net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput59 io_wbs_datrd_0[30] net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_65_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input26_I io_wbs_adr[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_100_ net2 _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_229_ net60 _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__351__I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__261__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__171__I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__236__A2 _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__346__I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input128_I io_wbs_datwr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__256__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input93_I io_wbs_datrd_1[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__166__I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output297_I net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput306 net306 io_wbs_sel_1[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input56_I io_wbs_datrd_0[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output212_I net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_331_ net123 net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_262_ net20 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_193_ _070_ _063_ _064_ _071_ net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_1_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__354__I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput147 net147 io_wbs_adr_0[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput158 net158 io_wbs_adr_0[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput169 net169 io_wbs_adr_0[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input110_I io_wbs_datwr[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__264__I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output162_I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_314_ net104 net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_245_ net33 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__174__I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput16 io_wbs_adr[21] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput27 io_wbs_adr[31] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_176_ _058_ _053_ _054_ _059_ net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xinput38 io_wbs_datrd_0[11] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput49 io_wbs_datrd_0[21] net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__349__I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__259__I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input19_I io_wbs_adr[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__169__I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_228_ net92 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_159_ _046_ _043_ _044_ _047_ net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__362__I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input86_I io_wbs_datrd_1[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output242_I net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__182__I _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__357__I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__267__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output192_I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__177__I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput307 net307 io_wbs_sel_1[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__118__A2 _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I io_wbs_datrd_0[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output205_I net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_330_ net121 net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_261_ net19 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_192_ net48 _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__370__I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput148 net148 io_wbs_adr_0[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput159 net159 io_wbs_adr_0[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input103_I io_wbs_datwr[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__280__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output155_I net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_313_ net103 net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_244_ net32 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput28 io_wbs_adr[3] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput17 io_wbs_adr[22] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_175_ net42 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput39 io_wbs_datrd_0[12] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__365__I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output272_I net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__185__I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_227_ _094_ _010_ _015_ _095_ net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_158_ net37 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input31_I io_wbs_adr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input79_I io_wbs_datrd_1[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output235_I net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__373__I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input133_I io_wbs_sel[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__283__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output185_I net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput308 net308 io_wbs_sel_1[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__368__I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_260_ net18 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_191_ net80 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__188__I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput138 net138 io_wbs_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput149 net149 io_wbs_adr_0[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input61_I io_wbs_datrd_0[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output148_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_312_ net102 net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_243_ net31 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput18 io_wbs_adr[23] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 io_wbs_adr[4] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_174_ net74 _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__291__I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output265_I net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_226_ net59 _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_157_ net69 _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input24_I io_wbs_adr[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__286__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__196__I _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_209_ _009_ _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output228_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input126_I io_wbs_datwr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input91_I io_wbs_datrd_1[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output178_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput309 net309 io_wbs_stb_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_4_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__294__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output295_I net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_190_ _068_ _063_ _064_ _069_ net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput139 net139 io_wbs_adr_0[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input54_I io_wbs_datrd_0[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__289__I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output210_I net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output308_I net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_311_ net101 net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_242_ net30 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 io_wbs_adr[24] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_173_ _056_ _053_ _054_ _057_ net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_2_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__199__I net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output160_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output258_I net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_225_ net91 _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_156_ _042_ _043_ _044_ _045_ net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input17_I io_wbs_adr[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_208_ net85 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_139_ _021_ _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I io_wbs_adr[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__297__I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input119_I io_wbs_datwr[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input84_I io_wbs_datrd_1[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output240_I net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output190_I net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output288_I net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input47_I io_wbs_datrd_0[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_310_ net131 net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_241_ net29 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_172_ net41 _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input101_I io_wbs_datwr[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output153_I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_224_ _092_ _010_ _015_ _093_ net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_155_ net67 _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output270_I net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput290 net290 io_wbs_datwr_1[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_75_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_207_ _080_ _073_ _074_ _081_ net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_138_ net95 _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input77_I io_wbs_datrd_1[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output233_I net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input131_I io_wbs_datwr[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output183_I net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_240_ net28 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_171_ net73 _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_369_ net132 net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__102__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output146_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_223_ net57 _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_154_ _023_ _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output263_I net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput280 net280 io_wbs_datwr_1[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput291 net291 io_wbs_datwr_1[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_206_ net52 _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_137_ _030_ _022_ _024_ _031_ net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input22_I io_wbs_adr[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output226_I net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__202__I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input124_I io_wbs_datwr[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output176_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__112__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output293_I net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_170_ _052_ _053_ _054_ _055_ net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_368_ net135 net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_299_ net26 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input52_I io_wbs_datrd_0[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__102__A2 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output139_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output306_I net306 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_222_ net89 _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_153_ _021_ _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__300__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__210__I _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput270 net270 io_wbs_datwr_1[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output256_I net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput281 net281 io_wbs_datwr_1[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput292 net292 io_wbs_datwr_1[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_58_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_205_ net84 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_136_ net62 _031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__205__I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input15_I io_wbs_adr[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__115__I _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_119_ net68 _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input7_I io_wbs_adr[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output219_I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input117_I io_wbs_datwr[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input82_I io_wbs_datrd_1[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output169_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__303__I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__213__I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output286_I net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__123__I _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_367_ net134 net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_298_ net24 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__208__I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input45_I io_wbs_datrd_0[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_221_ _090_ _083_ _084_ _091_ net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_152_ net99 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput271 net271 io_wbs_datwr_1[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput260 net260 io_wbs_datwr_0[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output151_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output249_I net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput282 net282 io_wbs_datwr_1[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput293 net293 io_wbs_datwr_1[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_75_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_204_ _078_ _073_ _074_ _079_ net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_135_ net94 _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__311__I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__232__A2 _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__306__I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_118_ _000_ _011_ _016_ _017_ net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__216__I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__126__I _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input75_I io_wbs_datrd_1[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output231_I net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output181_I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output279_I net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__105__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_366_ net133 net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_297_ net23 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__314__I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input38_I io_wbs_datrd_0[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_220_ net56 _091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_151_ _040_ _033_ _034_ _041_ net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_7_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__309__I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_349_ net107 net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__219__I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput250 net250 io_wbs_datwr_0[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput261 net261 io_wbs_datwr_0[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput294 net294 io_wbs_datwr_1[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput272 net272 io_wbs_datwr_1[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput283 net283 io_wbs_datwr_1[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output144_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__129__I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_203_ net51 _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_134_ _028_ _022_ _024_ _029_ net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output261_I net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_117_ net1 _017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__322__I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input20_I io_wbs_adr[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__317__I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input68_I io_wbs_datrd_1[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output224_I net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input122_I io_wbs_datwr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__105__A2 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output174_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_365_ net132 net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_296_ net22 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__330__I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output291_I net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_150_ net66 _041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__150__I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_348_ net106 net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__325__I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_279_ net4 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput262 net262 io_wbs_datwr_0[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput240 net240 io_wbs_datwr_0[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput251 net251 io_wbs_datwr_0[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input50_I io_wbs_datrd_0[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput295 net295 io_wbs_datwr_1[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput273 net273 io_wbs_datwr_1[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput284 net284 io_wbs_datwr_1[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_202_ net83 _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_133_ net61 _029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input98_I io_wbs_datrd_1[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output254_I net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_116_ _015_ _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input13_I io_wbs_adr[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__333__I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input5_I io_wbs_adr[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output217_I net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__328__I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input115_I io_wbs_datwr[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input80_I io_wbs_datrd_1[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__105__A3 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output167_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_364_ net124 net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_295_ net21 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output284_I net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_347_ net105 net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_278_ net34 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__341__I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__251__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput230 net230 io_wbs_datrd[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput241 net241 io_wbs_datwr_0[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput252 net252 io_wbs_datwr_0[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput263 net263 io_wbs_datwr_0[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput274 net274 io_wbs_datwr_1[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput285 net285 io_wbs_datwr_1[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_58_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input43_I io_wbs_datrd_0[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput296 net296 io_wbs_datwr_1[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_201_ _076_ _073_ _074_ _077_ net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_132_ net93 _028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__161__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__235__A2 _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__336__I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output247_I net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_115_ _014_ _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__108__A1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput130 io_wbs_datwr[8] net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__344__I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
.ends

