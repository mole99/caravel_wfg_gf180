magic
tech gf180mcuC
magscale 1 10
timestamp 1669806015
<< metal1 >>
rect 1344 36874 148624 36908
rect 1344 36822 19624 36874
rect 19676 36822 19728 36874
rect 19780 36822 19832 36874
rect 19884 36822 56444 36874
rect 56496 36822 56548 36874
rect 56600 36822 56652 36874
rect 56704 36822 93264 36874
rect 93316 36822 93368 36874
rect 93420 36822 93472 36874
rect 93524 36822 130084 36874
rect 130136 36822 130188 36874
rect 130240 36822 130292 36874
rect 130344 36822 148624 36874
rect 1344 36788 148624 36822
rect 30158 36706 30210 36718
rect 75070 36706 75122 36718
rect 35970 36654 35982 36706
rect 36034 36703 36046 36706
rect 36530 36703 36542 36706
rect 36034 36657 36542 36703
rect 36034 36654 36046 36657
rect 36530 36654 36542 36657
rect 36594 36654 36606 36706
rect 30158 36642 30210 36654
rect 75070 36642 75122 36654
rect 132414 36706 132466 36718
rect 132414 36642 132466 36654
rect 36094 36594 36146 36606
rect 64542 36594 64594 36606
rect 5954 36542 5966 36594
rect 6018 36542 6030 36594
rect 8194 36542 8206 36594
rect 8258 36542 8270 36594
rect 10434 36542 10446 36594
rect 10498 36542 10510 36594
rect 12114 36542 12126 36594
rect 12178 36542 12190 36594
rect 14466 36542 14478 36594
rect 14530 36542 14542 36594
rect 16034 36542 16046 36594
rect 16098 36542 16110 36594
rect 22194 36542 22206 36594
rect 22258 36542 22270 36594
rect 23874 36542 23886 36594
rect 23938 36542 23950 36594
rect 26002 36542 26014 36594
rect 26066 36542 26078 36594
rect 27794 36542 27806 36594
rect 27858 36542 27870 36594
rect 31490 36542 31502 36594
rect 31554 36542 31566 36594
rect 34626 36542 34638 36594
rect 34690 36542 34702 36594
rect 37762 36542 37774 36594
rect 37826 36542 37838 36594
rect 39554 36542 39566 36594
rect 39618 36542 39630 36594
rect 41346 36542 41358 36594
rect 41410 36542 41422 36594
rect 43138 36542 43150 36594
rect 43202 36542 43214 36594
rect 49522 36542 49534 36594
rect 49586 36542 49598 36594
rect 51314 36542 51326 36594
rect 51378 36542 51390 36594
rect 54898 36542 54910 36594
rect 54962 36542 54974 36594
rect 57922 36542 57934 36594
rect 57986 36542 57998 36594
rect 61058 36542 61070 36594
rect 61122 36542 61134 36594
rect 68898 36542 68910 36594
rect 68962 36542 68974 36594
rect 70578 36542 70590 36594
rect 70642 36542 70654 36594
rect 73378 36542 73390 36594
rect 73442 36542 73454 36594
rect 80882 36542 80894 36594
rect 80946 36542 80958 36594
rect 82674 36542 82686 36594
rect 82738 36542 82750 36594
rect 84802 36542 84814 36594
rect 84866 36542 84878 36594
rect 86146 36542 86158 36594
rect 86210 36542 86222 36594
rect 96562 36542 96574 36594
rect 96626 36542 96638 36594
rect 98354 36542 98366 36594
rect 98418 36542 98430 36594
rect 100034 36542 100046 36594
rect 100098 36542 100110 36594
rect 102386 36542 102398 36594
rect 102450 36542 102462 36594
rect 104402 36542 104414 36594
rect 104466 36542 104478 36594
rect 112242 36542 112254 36594
rect 112306 36542 112318 36594
rect 114034 36542 114046 36594
rect 114098 36542 114110 36594
rect 116610 36542 116622 36594
rect 116674 36542 116686 36594
rect 120194 36542 120206 36594
rect 120258 36542 120270 36594
rect 121986 36542 121998 36594
rect 122050 36542 122062 36594
rect 126018 36542 126030 36594
rect 126082 36542 126094 36594
rect 127922 36542 127934 36594
rect 127986 36542 127998 36594
rect 129714 36542 129726 36594
rect 129778 36542 129790 36594
rect 133746 36542 133758 36594
rect 133810 36542 133822 36594
rect 141586 36542 141598 36594
rect 141650 36542 141662 36594
rect 143602 36542 143614 36594
rect 143666 36542 143678 36594
rect 145394 36542 145406 36594
rect 145458 36542 145470 36594
rect 36094 36530 36146 36542
rect 64542 36530 64594 36542
rect 19742 36482 19794 36494
rect 33518 36482 33570 36494
rect 45726 36482 45778 36494
rect 6962 36430 6974 36482
rect 7026 36430 7038 36482
rect 7634 36430 7646 36482
rect 7698 36430 7710 36482
rect 9762 36430 9774 36482
rect 9826 36430 9838 36482
rect 12562 36430 12574 36482
rect 12626 36430 12638 36482
rect 13906 36430 13918 36482
rect 13970 36430 13982 36482
rect 16706 36430 16718 36482
rect 16770 36430 16782 36482
rect 18050 36430 18062 36482
rect 18114 36430 18126 36482
rect 21746 36430 21758 36482
rect 21810 36430 21822 36482
rect 24434 36430 24446 36482
rect 24498 36430 24510 36482
rect 26450 36430 26462 36482
rect 26514 36430 26526 36482
rect 28466 36430 28478 36482
rect 28530 36430 28542 36482
rect 32162 36430 32174 36482
rect 32226 36430 32238 36482
rect 35522 36430 35534 36482
rect 35586 36430 35598 36482
rect 38434 36430 38446 36482
rect 38498 36430 38510 36482
rect 40226 36430 40238 36482
rect 40290 36430 40302 36482
rect 42354 36430 42366 36482
rect 42418 36430 42430 36482
rect 44146 36430 44158 36482
rect 44210 36430 44222 36482
rect 19742 36418 19794 36430
rect 33518 36418 33570 36430
rect 45726 36418 45778 36430
rect 47518 36482 47570 36494
rect 53678 36482 53730 36494
rect 63310 36482 63362 36494
rect 48962 36430 48974 36482
rect 49026 36430 49038 36482
rect 51986 36430 51998 36482
rect 52050 36430 52062 36482
rect 52994 36430 53006 36482
rect 53058 36430 53070 36482
rect 55906 36430 55918 36482
rect 55970 36430 55982 36482
rect 58818 36430 58830 36482
rect 58882 36430 58894 36482
rect 61730 36430 61742 36482
rect 61794 36430 61806 36482
rect 62738 36430 62750 36482
rect 62802 36430 62814 36482
rect 47518 36418 47570 36430
rect 53678 36418 53730 36430
rect 63310 36418 63362 36430
rect 64990 36482 65042 36494
rect 66782 36482 66834 36494
rect 77422 36482 77474 36494
rect 87950 36482 88002 36494
rect 66098 36430 66110 36482
rect 66162 36430 66174 36482
rect 69682 36430 69694 36482
rect 69746 36430 69758 36482
rect 71474 36430 71486 36482
rect 71538 36430 71550 36482
rect 72370 36430 72382 36482
rect 72434 36430 72446 36482
rect 74386 36430 74398 36482
rect 74450 36430 74462 36482
rect 76738 36430 76750 36482
rect 76802 36430 76814 36482
rect 80434 36430 80446 36482
rect 80498 36430 80510 36482
rect 82002 36430 82014 36482
rect 82066 36430 82078 36482
rect 84130 36430 84142 36482
rect 84194 36430 84206 36482
rect 86930 36430 86942 36482
rect 86994 36430 87006 36482
rect 64990 36418 65042 36430
rect 66782 36418 66834 36430
rect 77422 36418 77474 36430
rect 87950 36418 88002 36430
rect 88958 36482 89010 36494
rect 94334 36482 94386 36494
rect 106430 36482 106482 36494
rect 109342 36482 109394 36494
rect 123790 36482 123842 36494
rect 132078 36482 132130 36494
rect 136558 36482 136610 36494
rect 139918 36482 139970 36494
rect 89730 36430 89742 36482
rect 89794 36430 89806 36482
rect 92194 36430 92206 36482
rect 92258 36430 92270 36482
rect 93650 36430 93662 36482
rect 93714 36430 93726 36482
rect 96114 36430 96126 36482
rect 96178 36430 96190 36482
rect 97906 36430 97918 36482
rect 97970 36430 97982 36482
rect 100818 36430 100830 36482
rect 100882 36430 100894 36482
rect 101602 36430 101614 36482
rect 101666 36430 101678 36482
rect 103730 36430 103742 36482
rect 103794 36430 103806 36482
rect 108658 36430 108670 36482
rect 108722 36430 108734 36482
rect 111570 36430 111582 36482
rect 111634 36430 111646 36482
rect 113362 36430 113374 36482
rect 113426 36430 113438 36482
rect 115938 36430 115950 36482
rect 116002 36430 116014 36482
rect 117842 36430 117854 36482
rect 117906 36430 117918 36482
rect 119522 36430 119534 36482
rect 119586 36430 119598 36482
rect 121314 36430 121326 36482
rect 121378 36430 121390 36482
rect 124562 36430 124574 36482
rect 124626 36430 124638 36482
rect 125234 36430 125246 36482
rect 125298 36430 125310 36482
rect 127250 36430 127262 36482
rect 127314 36430 127326 36482
rect 129266 36430 129278 36482
rect 129330 36430 129342 36482
rect 131394 36430 131406 36482
rect 131458 36430 131470 36482
rect 133074 36430 133086 36482
rect 133138 36430 133150 36482
rect 137778 36430 137790 36482
rect 137842 36430 137854 36482
rect 139234 36430 139246 36482
rect 139298 36430 139310 36482
rect 141026 36430 141038 36482
rect 141090 36430 141102 36482
rect 142930 36430 142942 36482
rect 142994 36430 143006 36482
rect 144946 36430 144958 36482
rect 145010 36430 145022 36482
rect 88958 36418 89010 36430
rect 94334 36418 94386 36430
rect 106430 36418 106482 36430
rect 109342 36418 109394 36430
rect 123790 36418 123842 36430
rect 132078 36418 132130 36430
rect 136558 36418 136610 36430
rect 139918 36418 139970 36430
rect 4846 36370 4898 36382
rect 4846 36306 4898 36318
rect 17502 36370 17554 36382
rect 33854 36370 33906 36382
rect 56814 36370 56866 36382
rect 18946 36318 18958 36370
rect 19010 36318 19022 36370
rect 19506 36318 19518 36370
rect 19570 36318 19582 36370
rect 29474 36318 29486 36370
rect 29538 36318 29550 36370
rect 29810 36318 29822 36370
rect 29874 36318 29886 36370
rect 46834 36318 46846 36370
rect 46898 36318 46910 36370
rect 47170 36318 47182 36370
rect 47234 36318 47246 36370
rect 52882 36318 52894 36370
rect 52946 36318 52958 36370
rect 17502 36306 17554 36318
rect 33854 36306 33906 36318
rect 56814 36306 56866 36318
rect 57150 36370 57202 36382
rect 57150 36306 57202 36318
rect 59502 36370 59554 36382
rect 65326 36370 65378 36382
rect 67790 36370 67842 36382
rect 78766 36370 78818 36382
rect 90750 36370 90802 36382
rect 62514 36318 62526 36370
rect 62578 36318 62590 36370
rect 65986 36318 65998 36370
rect 66050 36318 66062 36370
rect 74274 36318 74286 36370
rect 74338 36318 74350 36370
rect 76626 36318 76638 36370
rect 76690 36318 76702 36370
rect 89506 36318 89518 36370
rect 89570 36318 89582 36370
rect 59502 36306 59554 36318
rect 65326 36306 65378 36318
rect 67790 36306 67842 36318
rect 78766 36306 78818 36318
rect 90750 36306 90802 36318
rect 91198 36370 91250 36382
rect 91198 36306 91250 36318
rect 91982 36370 92034 36382
rect 110350 36370 110402 36382
rect 93762 36318 93774 36370
rect 93826 36318 93838 36370
rect 105634 36318 105646 36370
rect 105698 36318 105710 36370
rect 106194 36318 106206 36370
rect 106258 36318 106270 36370
rect 108546 36318 108558 36370
rect 108610 36318 108622 36370
rect 91982 36306 92034 36318
rect 110350 36306 110402 36318
rect 110686 36370 110738 36382
rect 110686 36306 110738 36318
rect 118078 36370 118130 36382
rect 124338 36318 124350 36370
rect 124402 36318 124414 36370
rect 131282 36318 131294 36370
rect 131346 36318 131358 36370
rect 135762 36318 135774 36370
rect 135826 36318 135838 36370
rect 136210 36318 136222 36370
rect 136274 36318 136286 36370
rect 139122 36318 139134 36370
rect 139186 36318 139198 36370
rect 118078 36306 118130 36318
rect 18286 36258 18338 36270
rect 18286 36194 18338 36206
rect 20078 36258 20130 36270
rect 20078 36194 20130 36206
rect 20750 36258 20802 36270
rect 20750 36194 20802 36206
rect 30494 36258 30546 36270
rect 30494 36194 30546 36206
rect 45278 36258 45330 36270
rect 45278 36194 45330 36206
rect 46062 36258 46114 36270
rect 46062 36194 46114 36206
rect 47854 36258 47906 36270
rect 47854 36194 47906 36206
rect 54014 36258 54066 36270
rect 54014 36194 54066 36206
rect 59838 36258 59890 36270
rect 59838 36194 59890 36206
rect 63646 36258 63698 36270
rect 63646 36194 63698 36206
rect 67118 36258 67170 36270
rect 67118 36194 67170 36206
rect 75406 36258 75458 36270
rect 75406 36194 75458 36206
rect 77758 36258 77810 36270
rect 77758 36194 77810 36206
rect 78430 36258 78482 36270
rect 78430 36194 78482 36206
rect 79214 36258 79266 36270
rect 79214 36194 79266 36206
rect 88622 36258 88674 36270
rect 88622 36194 88674 36206
rect 90414 36258 90466 36270
rect 90414 36194 90466 36206
rect 92766 36258 92818 36270
rect 92766 36194 92818 36206
rect 94670 36258 94722 36270
rect 94670 36194 94722 36206
rect 106766 36258 106818 36270
rect 106766 36194 106818 36206
rect 107550 36258 107602 36270
rect 107550 36194 107602 36206
rect 109678 36258 109730 36270
rect 109678 36194 109730 36206
rect 115502 36258 115554 36270
rect 115502 36194 115554 36206
rect 118526 36258 118578 36270
rect 118526 36194 118578 36206
rect 123454 36258 123506 36270
rect 123454 36194 123506 36206
rect 134990 36258 135042 36270
rect 134990 36194 135042 36206
rect 136894 36258 136946 36270
rect 136894 36194 136946 36206
rect 137566 36258 137618 36270
rect 137566 36194 137618 36206
rect 140254 36258 140306 36270
rect 140254 36194 140306 36206
rect 1344 36090 148784 36124
rect 1344 36038 38034 36090
rect 38086 36038 38138 36090
rect 38190 36038 38242 36090
rect 38294 36038 74854 36090
rect 74906 36038 74958 36090
rect 75010 36038 75062 36090
rect 75114 36038 111674 36090
rect 111726 36038 111778 36090
rect 111830 36038 111882 36090
rect 111934 36038 148494 36090
rect 148546 36038 148598 36090
rect 148650 36038 148702 36090
rect 148754 36038 148784 36090
rect 1344 36004 148784 36038
rect 6078 35922 6130 35934
rect 6078 35858 6130 35870
rect 8990 35922 9042 35934
rect 8990 35858 9042 35870
rect 19518 35922 19570 35934
rect 19518 35858 19570 35870
rect 23102 35922 23154 35934
rect 23102 35858 23154 35870
rect 26574 35922 26626 35934
rect 26574 35858 26626 35870
rect 39006 35922 39058 35934
rect 39006 35858 39058 35870
rect 41806 35922 41858 35934
rect 41806 35858 41858 35870
rect 42366 35922 42418 35934
rect 42366 35858 42418 35870
rect 43262 35922 43314 35934
rect 43262 35858 43314 35870
rect 54574 35922 54626 35934
rect 54574 35858 54626 35870
rect 57598 35922 57650 35934
rect 57598 35858 57650 35870
rect 58942 35922 58994 35934
rect 64542 35922 64594 35934
rect 61282 35870 61294 35922
rect 61346 35870 61358 35922
rect 58942 35858 58994 35870
rect 64542 35858 64594 35870
rect 70814 35922 70866 35934
rect 70814 35858 70866 35870
rect 73950 35922 74002 35934
rect 73950 35858 74002 35870
rect 80334 35922 80386 35934
rect 80334 35858 80386 35870
rect 92990 35922 93042 35934
rect 92990 35858 93042 35870
rect 97246 35922 97298 35934
rect 97246 35858 97298 35870
rect 99822 35922 99874 35934
rect 99822 35858 99874 35870
rect 100606 35922 100658 35934
rect 100606 35858 100658 35870
rect 101166 35922 101218 35934
rect 101166 35858 101218 35870
rect 104190 35922 104242 35934
rect 104190 35858 104242 35870
rect 111358 35922 111410 35934
rect 111358 35858 111410 35870
rect 113150 35922 113202 35934
rect 113150 35858 113202 35870
rect 116846 35922 116898 35934
rect 116846 35858 116898 35870
rect 119870 35922 119922 35934
rect 119870 35858 119922 35870
rect 121102 35922 121154 35934
rect 121102 35858 121154 35870
rect 122334 35922 122386 35934
rect 122334 35858 122386 35870
rect 132974 35922 133026 35934
rect 132974 35858 133026 35870
rect 137902 35922 137954 35934
rect 137902 35858 137954 35870
rect 142158 35922 142210 35934
rect 142158 35858 142210 35870
rect 144958 35922 145010 35934
rect 144958 35858 145010 35870
rect 145854 35922 145906 35934
rect 145854 35858 145906 35870
rect 146638 35922 146690 35934
rect 146638 35858 146690 35870
rect 10558 35810 10610 35822
rect 7522 35758 7534 35810
rect 7586 35758 7598 35810
rect 10558 35746 10610 35758
rect 13246 35810 13298 35822
rect 20414 35810 20466 35822
rect 39902 35810 39954 35822
rect 17826 35758 17838 35810
rect 17890 35758 17902 35810
rect 30146 35758 30158 35810
rect 30210 35758 30222 35810
rect 34514 35758 34526 35810
rect 34578 35758 34590 35810
rect 36530 35758 36542 35810
rect 36594 35758 36606 35810
rect 13246 35746 13298 35758
rect 20414 35746 20466 35758
rect 39902 35746 39954 35758
rect 40798 35810 40850 35822
rect 46398 35810 46450 35822
rect 53678 35810 53730 35822
rect 43922 35758 43934 35810
rect 43986 35758 43998 35810
rect 44370 35758 44382 35810
rect 44434 35758 44446 35810
rect 50306 35758 50318 35810
rect 50370 35758 50382 35810
rect 51874 35758 51886 35810
rect 51938 35758 51950 35810
rect 52434 35758 52446 35810
rect 52498 35758 52510 35810
rect 40798 35746 40850 35758
rect 46398 35746 46450 35758
rect 53678 35746 53730 35758
rect 54014 35810 54066 35822
rect 58606 35810 58658 35822
rect 64206 35810 64258 35822
rect 69918 35810 69970 35822
rect 55794 35758 55806 35810
rect 55858 35758 55870 35810
rect 62402 35758 62414 35810
rect 62466 35758 62478 35810
rect 65762 35758 65774 35810
rect 65826 35758 65838 35810
rect 67890 35758 67902 35810
rect 67954 35758 67966 35810
rect 54014 35746 54066 35758
rect 58606 35746 58658 35758
rect 64206 35746 64258 35758
rect 69918 35746 69970 35758
rect 70478 35810 70530 35822
rect 83470 35810 83522 35822
rect 74722 35758 74734 35810
rect 74786 35758 74798 35810
rect 76850 35758 76862 35810
rect 76914 35758 76926 35810
rect 70478 35746 70530 35758
rect 83470 35746 83522 35758
rect 86382 35810 86434 35822
rect 95342 35810 95394 35822
rect 89394 35758 89406 35810
rect 89458 35758 89470 35810
rect 89954 35758 89966 35810
rect 90018 35758 90030 35810
rect 93650 35758 93662 35810
rect 93714 35758 93726 35810
rect 86382 35746 86434 35758
rect 95342 35746 95394 35758
rect 101614 35810 101666 35822
rect 105534 35810 105586 35822
rect 108334 35810 108386 35822
rect 112254 35810 112306 35822
rect 102834 35758 102846 35810
rect 102898 35758 102910 35810
rect 106306 35758 106318 35810
rect 106370 35758 106382 35810
rect 109330 35758 109342 35810
rect 109394 35758 109406 35810
rect 101614 35746 101666 35758
rect 105534 35746 105586 35758
rect 108334 35746 108386 35758
rect 112254 35746 112306 35758
rect 116286 35810 116338 35822
rect 129614 35810 129666 35822
rect 135662 35810 135714 35822
rect 146190 35810 146242 35822
rect 124450 35758 124462 35810
rect 124514 35758 124526 35810
rect 126242 35758 126254 35810
rect 126306 35758 126318 35810
rect 130834 35758 130846 35810
rect 130898 35758 130910 35810
rect 131394 35758 131406 35810
rect 131458 35758 131470 35810
rect 134754 35758 134766 35810
rect 134818 35758 134830 35810
rect 138674 35758 138686 35810
rect 138738 35758 138750 35810
rect 140578 35758 140590 35810
rect 140642 35758 140654 35810
rect 143714 35758 143726 35810
rect 143778 35758 143790 35810
rect 116286 35746 116338 35758
rect 129614 35746 129666 35758
rect 135662 35746 135714 35758
rect 146190 35746 146242 35758
rect 20078 35698 20130 35710
rect 26238 35698 26290 35710
rect 29374 35698 29426 35710
rect 38670 35698 38722 35710
rect 6626 35646 6638 35698
rect 6690 35646 6702 35698
rect 8754 35646 8766 35698
rect 8818 35646 8830 35698
rect 10322 35646 10334 35698
rect 10386 35646 10398 35698
rect 11106 35646 11118 35698
rect 11170 35646 11182 35698
rect 13010 35646 13022 35698
rect 13074 35646 13086 35698
rect 13794 35646 13806 35698
rect 13858 35646 13870 35698
rect 15922 35646 15934 35698
rect 15986 35646 15998 35698
rect 18162 35646 18174 35698
rect 18226 35646 18238 35698
rect 20962 35646 20974 35698
rect 21026 35646 21038 35698
rect 22866 35646 22878 35698
rect 22930 35646 22942 35698
rect 23650 35646 23662 35698
rect 23714 35646 23726 35698
rect 28130 35646 28142 35698
rect 28194 35646 28206 35698
rect 29810 35646 29822 35698
rect 29874 35646 29886 35698
rect 30818 35646 30830 35698
rect 30882 35646 30894 35698
rect 33618 35646 33630 35698
rect 33682 35646 33694 35698
rect 37426 35646 37438 35698
rect 37490 35646 37502 35698
rect 20078 35634 20130 35646
rect 26238 35634 26290 35646
rect 29374 35634 29426 35646
rect 38670 35634 38722 35646
rect 39566 35698 39618 35710
rect 42702 35698 42754 35710
rect 52670 35698 52722 35710
rect 40562 35646 40574 35698
rect 40626 35646 40638 35698
rect 46162 35646 46174 35698
rect 46226 35646 46238 35698
rect 46946 35646 46958 35698
rect 47010 35646 47022 35698
rect 51202 35646 51214 35698
rect 51266 35646 51278 35698
rect 39566 35634 39618 35646
rect 42702 35634 42754 35646
rect 52670 35634 52722 35646
rect 54910 35698 54962 35710
rect 69582 35698 69634 35710
rect 77534 35698 77586 35710
rect 90190 35698 90242 35710
rect 94334 35698 94386 35710
rect 105198 35698 105250 35710
rect 107998 35698 108050 35710
rect 111022 35698 111074 35710
rect 113486 35698 113538 35710
rect 121998 35698 122050 35710
rect 127934 35698 127986 35710
rect 56690 35646 56702 35698
rect 56754 35646 56766 35698
rect 57810 35646 57822 35698
rect 57874 35646 57886 35698
rect 60722 35646 60734 35698
rect 60786 35646 60798 35698
rect 61506 35646 61518 35698
rect 61570 35646 61582 35698
rect 62738 35646 62750 35698
rect 62802 35646 62814 35698
rect 66098 35646 66110 35698
rect 66162 35646 66174 35698
rect 68786 35646 68798 35698
rect 68850 35646 68862 35698
rect 72594 35646 72606 35698
rect 72658 35646 72670 35698
rect 73714 35646 73726 35698
rect 73778 35646 73790 35698
rect 74610 35646 74622 35698
rect 74674 35646 74686 35698
rect 76738 35646 76750 35698
rect 76802 35646 76814 35698
rect 78530 35646 78542 35698
rect 78594 35646 78606 35698
rect 81330 35646 81342 35698
rect 81394 35646 81406 35698
rect 83234 35646 83246 35698
rect 83298 35646 83310 35698
rect 84578 35646 84590 35698
rect 84642 35646 84654 35698
rect 86594 35646 86606 35698
rect 86658 35646 86670 35698
rect 87378 35646 87390 35698
rect 87442 35646 87454 35698
rect 91186 35646 91198 35698
rect 91250 35646 91262 35698
rect 93538 35646 93550 35698
rect 93602 35646 93614 35698
rect 95554 35646 95566 35698
rect 95618 35646 95630 35698
rect 98018 35646 98030 35698
rect 98082 35646 98094 35698
rect 100034 35646 100046 35698
rect 100098 35646 100110 35698
rect 101826 35646 101838 35698
rect 101890 35646 101902 35698
rect 103506 35646 103518 35698
rect 103570 35646 103582 35698
rect 106194 35646 106206 35698
rect 106258 35646 106270 35698
rect 109218 35646 109230 35698
rect 109282 35646 109294 35698
rect 112018 35646 112030 35698
rect 112082 35646 112094 35698
rect 114258 35646 114270 35698
rect 114322 35646 114334 35698
rect 116050 35646 116062 35698
rect 116114 35646 116126 35698
rect 117058 35646 117070 35698
rect 117122 35646 117134 35698
rect 117730 35646 117742 35698
rect 117794 35646 117806 35698
rect 119634 35646 119646 35698
rect 119698 35646 119710 35698
rect 121314 35646 121326 35698
rect 121378 35646 121390 35698
rect 124562 35646 124574 35698
rect 124626 35646 124638 35698
rect 125346 35646 125358 35698
rect 125410 35646 125422 35698
rect 54910 35634 54962 35646
rect 69582 35634 69634 35646
rect 77534 35634 77586 35646
rect 90190 35634 90242 35646
rect 94334 35634 94386 35646
rect 105198 35634 105250 35646
rect 107998 35634 108050 35646
rect 111022 35634 111074 35646
rect 113486 35634 113538 35646
rect 121998 35634 122050 35646
rect 127934 35634 127986 35646
rect 129054 35698 129106 35710
rect 129054 35634 129106 35646
rect 130062 35698 130114 35710
rect 130062 35634 130114 35646
rect 132638 35698 132690 35710
rect 136894 35698 136946 35710
rect 133858 35646 133870 35698
rect 133922 35646 133934 35698
rect 135874 35646 135886 35698
rect 135938 35646 135950 35698
rect 137666 35646 137678 35698
rect 137730 35646 137742 35698
rect 138562 35646 138574 35698
rect 138626 35646 138638 35698
rect 140466 35646 140478 35698
rect 140530 35646 140542 35698
rect 142818 35646 142830 35698
rect 142882 35646 142894 35698
rect 145170 35646 145182 35698
rect 145234 35646 145246 35698
rect 132638 35634 132690 35646
rect 136894 35634 136946 35646
rect 9662 35586 9714 35598
rect 25678 35586 25730 35598
rect 32622 35586 32674 35598
rect 11778 35534 11790 35586
rect 11842 35534 11854 35586
rect 14466 35534 14478 35586
rect 14530 35534 14542 35586
rect 16370 35534 16382 35586
rect 16434 35534 16446 35586
rect 21634 35534 21646 35586
rect 21698 35534 21710 35586
rect 24322 35534 24334 35586
rect 24386 35534 24398 35586
rect 27346 35534 27358 35586
rect 27410 35534 27422 35586
rect 31490 35534 31502 35586
rect 31554 35534 31566 35586
rect 9662 35522 9714 35534
rect 25678 35522 25730 35534
rect 32622 35522 32674 35534
rect 38110 35586 38162 35598
rect 38110 35522 38162 35534
rect 45614 35586 45666 35598
rect 48750 35586 48802 35598
rect 47618 35534 47630 35586
rect 47682 35534 47694 35586
rect 45614 35522 45666 35534
rect 48750 35522 48802 35534
rect 49422 35586 49474 35598
rect 83918 35586 83970 35598
rect 96126 35586 96178 35598
rect 107326 35586 107378 35598
rect 120318 35586 120370 35598
rect 59714 35534 59726 35586
rect 59778 35534 59790 35586
rect 71810 35534 71822 35586
rect 71874 35534 71886 35586
rect 79202 35534 79214 35586
rect 79266 35534 79278 35586
rect 82002 35534 82014 35586
rect 82066 35534 82078 35586
rect 85250 35534 85262 35586
rect 85314 35534 85326 35586
rect 87938 35534 87950 35586
rect 88002 35534 88014 35586
rect 91858 35534 91870 35586
rect 91922 35534 91934 35586
rect 98690 35534 98702 35586
rect 98754 35534 98766 35586
rect 114818 35534 114830 35586
rect 114882 35534 114894 35586
rect 118402 35534 118414 35586
rect 118466 35534 118478 35586
rect 49422 35522 49474 35534
rect 83918 35522 83970 35534
rect 96126 35522 96178 35534
rect 107326 35522 107378 35534
rect 120318 35522 120370 35534
rect 122782 35586 122834 35598
rect 122782 35522 122834 35534
rect 127374 35586 127426 35598
rect 127374 35522 127426 35534
rect 131630 35586 131682 35598
rect 131630 35522 131682 35534
rect 141262 35586 141314 35598
rect 141262 35522 141314 35534
rect 18622 35474 18674 35486
rect 18622 35410 18674 35422
rect 18958 35474 19010 35486
rect 18958 35410 19010 35422
rect 29038 35474 29090 35486
rect 29038 35410 29090 35422
rect 44606 35474 44658 35486
rect 44606 35410 44658 35422
rect 44942 35474 44994 35486
rect 44942 35410 44994 35422
rect 53006 35474 53058 35486
rect 53006 35410 53058 35422
rect 63198 35474 63250 35486
rect 63198 35410 63250 35422
rect 63534 35474 63586 35486
rect 63534 35410 63586 35422
rect 66558 35474 66610 35486
rect 66558 35410 66610 35422
rect 66894 35474 66946 35486
rect 66894 35410 66946 35422
rect 75406 35474 75458 35486
rect 75406 35410 75458 35422
rect 75742 35474 75794 35486
rect 75742 35410 75794 35422
rect 77870 35474 77922 35486
rect 77870 35410 77922 35422
rect 90526 35474 90578 35486
rect 90526 35410 90578 35422
rect 94670 35474 94722 35486
rect 94670 35410 94722 35422
rect 106990 35474 107042 35486
rect 106990 35410 107042 35422
rect 110014 35474 110066 35486
rect 110014 35410 110066 35422
rect 110350 35474 110402 35486
rect 110350 35410 110402 35422
rect 123566 35474 123618 35486
rect 123566 35410 123618 35422
rect 123902 35474 123954 35486
rect 123902 35410 123954 35422
rect 131966 35474 132018 35486
rect 131966 35410 132018 35422
rect 139358 35474 139410 35486
rect 139358 35410 139410 35422
rect 139694 35474 139746 35486
rect 139694 35410 139746 35422
rect 141598 35474 141650 35486
rect 141598 35410 141650 35422
rect 1344 35306 148624 35340
rect 1344 35254 19624 35306
rect 19676 35254 19728 35306
rect 19780 35254 19832 35306
rect 19884 35254 56444 35306
rect 56496 35254 56548 35306
rect 56600 35254 56652 35306
rect 56704 35254 93264 35306
rect 93316 35254 93368 35306
rect 93420 35254 93472 35306
rect 93524 35254 130084 35306
rect 130136 35254 130188 35306
rect 130240 35254 130292 35306
rect 130344 35254 148624 35306
rect 1344 35220 148624 35254
rect 53790 35138 53842 35150
rect 53790 35074 53842 35086
rect 11006 35026 11058 35038
rect 31390 35026 31442 35038
rect 10098 34974 10110 35026
rect 10162 34974 10174 35026
rect 18498 34974 18510 35026
rect 18562 34974 18574 35026
rect 20290 34974 20302 35026
rect 20354 34974 20366 35026
rect 11006 34962 11058 34974
rect 31390 34962 31442 34974
rect 42030 35026 42082 35038
rect 42030 34962 42082 34974
rect 43374 35026 43426 35038
rect 43374 34962 43426 34974
rect 43822 35026 43874 35038
rect 53454 35026 53506 35038
rect 45714 34974 45726 35026
rect 45778 34974 45790 35026
rect 43822 34962 43874 34974
rect 53454 34962 53506 34974
rect 56030 35026 56082 35038
rect 56030 34962 56082 34974
rect 59614 35026 59666 35038
rect 66670 35026 66722 35038
rect 63410 34974 63422 35026
rect 63474 34974 63486 35026
rect 65090 34974 65102 35026
rect 65154 34974 65166 35026
rect 59614 34962 59666 34974
rect 66670 34962 66722 34974
rect 68686 35026 68738 35038
rect 68686 34962 68738 34974
rect 70142 35026 70194 35038
rect 70142 34962 70194 34974
rect 71038 35026 71090 35038
rect 71038 34962 71090 34974
rect 71598 35026 71650 35038
rect 71598 34962 71650 34974
rect 72046 35026 72098 35038
rect 72046 34962 72098 34974
rect 72494 35026 72546 35038
rect 99598 35026 99650 35038
rect 77970 34974 77982 35026
rect 78034 34974 78046 35026
rect 82562 34974 82574 35026
rect 82626 34974 82638 35026
rect 88834 34974 88846 35026
rect 88898 34974 88910 35026
rect 90178 34974 90190 35026
rect 90242 34974 90254 35026
rect 93986 34974 93998 35026
rect 94050 34974 94062 35026
rect 96002 34974 96014 35026
rect 96066 34974 96078 35026
rect 72494 34962 72546 34974
rect 99598 34962 99650 34974
rect 103854 35026 103906 35038
rect 117070 35026 117122 35038
rect 105858 34974 105870 35026
rect 105922 34974 105934 35026
rect 107650 34974 107662 35026
rect 107714 34974 107726 35026
rect 109778 34974 109790 35026
rect 109842 34974 109854 35026
rect 103854 34962 103906 34974
rect 117070 34962 117122 34974
rect 120430 35026 120482 35038
rect 120430 34962 120482 34974
rect 120990 35026 121042 35038
rect 139134 35026 139186 35038
rect 131058 34974 131070 35026
rect 131122 34974 131134 35026
rect 136322 34974 136334 35026
rect 136386 34974 136398 35026
rect 138114 34974 138126 35026
rect 138178 34974 138190 35026
rect 120990 34962 121042 34974
rect 139134 34962 139186 34974
rect 145518 35026 145570 35038
rect 145518 34962 145570 34974
rect 6190 34914 6242 34926
rect 6190 34850 6242 34862
rect 6974 34914 7026 34926
rect 6974 34850 7026 34862
rect 7870 34914 7922 34926
rect 12910 34914 12962 34926
rect 8530 34862 8542 34914
rect 8594 34862 8606 34914
rect 9314 34862 9326 34914
rect 9378 34862 9390 34914
rect 11778 34862 11790 34914
rect 11842 34862 11854 34914
rect 7870 34850 7922 34862
rect 12910 34850 12962 34862
rect 13582 34914 13634 34926
rect 13582 34850 13634 34862
rect 14590 34914 14642 34926
rect 22766 34914 22818 34926
rect 15250 34862 15262 34914
rect 15314 34862 15326 34914
rect 17154 34862 17166 34914
rect 17218 34862 17230 34914
rect 18050 34862 18062 34914
rect 18114 34862 18126 34914
rect 19618 34862 19630 34914
rect 19682 34862 19694 34914
rect 14590 34850 14642 34862
rect 22766 34850 22818 34862
rect 23998 34914 24050 34926
rect 23998 34850 24050 34862
rect 25454 34914 25506 34926
rect 25454 34850 25506 34862
rect 29934 34914 29986 34926
rect 37774 34914 37826 34926
rect 42478 34914 42530 34926
rect 30594 34862 30606 34914
rect 30658 34862 30670 34914
rect 32834 34862 32846 34914
rect 32898 34862 32910 34914
rect 36530 34862 36542 34914
rect 36594 34862 36606 34914
rect 38322 34862 38334 34914
rect 38386 34862 38398 34914
rect 40114 34862 40126 34914
rect 40178 34862 40190 34914
rect 29934 34850 29986 34862
rect 37774 34850 37826 34862
rect 42478 34850 42530 34862
rect 44270 34914 44322 34926
rect 49534 34914 49586 34926
rect 54574 34914 54626 34926
rect 46610 34862 46622 34914
rect 46674 34862 46686 34914
rect 50642 34862 50654 34914
rect 50706 34862 50718 34914
rect 44270 34850 44322 34862
rect 49534 34850 49586 34862
rect 54574 34850 54626 34862
rect 55022 34914 55074 34926
rect 55022 34850 55074 34862
rect 57374 34914 57426 34926
rect 57374 34850 57426 34862
rect 58606 34914 58658 34926
rect 58606 34850 58658 34862
rect 62190 34914 62242 34926
rect 67118 34914 67170 34926
rect 64306 34862 64318 34914
rect 64370 34862 64382 34914
rect 66098 34862 66110 34914
rect 66162 34862 66174 34914
rect 62190 34850 62242 34862
rect 67118 34850 67170 34862
rect 67566 34914 67618 34926
rect 67566 34850 67618 34862
rect 69358 34914 69410 34926
rect 69358 34850 69410 34862
rect 72942 34914 72994 34926
rect 72942 34850 72994 34862
rect 73838 34914 73890 34926
rect 73838 34850 73890 34862
rect 74734 34914 74786 34926
rect 74734 34850 74786 34862
rect 75854 34914 75906 34926
rect 75854 34850 75906 34862
rect 76190 34914 76242 34926
rect 117854 34914 117906 34926
rect 129390 34914 129442 34926
rect 131966 34914 132018 34926
rect 140926 34914 140978 34926
rect 77298 34862 77310 34914
rect 77362 34862 77374 34914
rect 79538 34862 79550 34914
rect 79602 34862 79614 34914
rect 81890 34862 81902 34914
rect 81954 34862 81966 34914
rect 88162 34862 88174 34914
rect 88226 34862 88238 34914
rect 90962 34862 90974 34914
rect 91026 34862 91038 34914
rect 93426 34862 93438 34914
rect 93490 34862 93502 34914
rect 95330 34862 95342 34914
rect 95394 34862 95406 34914
rect 97346 34862 97358 34914
rect 97410 34862 97422 34914
rect 104514 34862 104526 34914
rect 104578 34862 104590 34914
rect 105186 34862 105198 34914
rect 105250 34862 105262 34914
rect 106978 34862 106990 34914
rect 107042 34862 107054 34914
rect 109218 34862 109230 34914
rect 109282 34862 109294 34914
rect 111682 34862 111694 34914
rect 111746 34862 111758 34914
rect 115266 34862 115278 34914
rect 115330 34862 115342 34914
rect 119858 34862 119870 34914
rect 119922 34862 119934 34914
rect 122658 34862 122670 34914
rect 122722 34862 122734 34914
rect 125234 34862 125246 34914
rect 125298 34862 125310 34914
rect 127026 34862 127038 34914
rect 127090 34862 127102 34914
rect 128818 34862 128830 34914
rect 128882 34862 128894 34914
rect 130498 34862 130510 34914
rect 130562 34862 130574 34914
rect 133186 34862 133198 34914
rect 133250 34862 133262 34914
rect 135762 34862 135774 34914
rect 135826 34862 135838 34914
rect 137442 34862 137454 34914
rect 137506 34862 137518 34914
rect 140018 34862 140030 34914
rect 140082 34862 140094 34914
rect 143938 34862 143950 34914
rect 144002 34862 144014 34914
rect 76190 34850 76242 34862
rect 117854 34850 117906 34862
rect 129390 34850 129442 34862
rect 131966 34850 132018 34862
rect 140926 34850 140978 34862
rect 6638 34802 6690 34814
rect 6638 34738 6690 34750
rect 7534 34802 7586 34814
rect 7534 34738 7586 34750
rect 8766 34802 8818 34814
rect 8766 34738 8818 34750
rect 12014 34802 12066 34814
rect 12014 34738 12066 34750
rect 12574 34802 12626 34814
rect 12574 34738 12626 34750
rect 14254 34802 14306 34814
rect 14254 34738 14306 34750
rect 16046 34802 16098 34814
rect 16046 34738 16098 34750
rect 16382 34802 16434 34814
rect 16382 34738 16434 34750
rect 16942 34802 16994 34814
rect 16942 34738 16994 34750
rect 21870 34802 21922 34814
rect 21870 34738 21922 34750
rect 22206 34802 22258 34814
rect 22206 34738 22258 34750
rect 23102 34802 23154 34814
rect 23102 34738 23154 34750
rect 23662 34802 23714 34814
rect 23662 34738 23714 34750
rect 24558 34802 24610 34814
rect 24558 34738 24610 34750
rect 24894 34802 24946 34814
rect 24894 34738 24946 34750
rect 25790 34802 25842 34814
rect 25790 34738 25842 34750
rect 26574 34802 26626 34814
rect 26574 34738 26626 34750
rect 26910 34802 26962 34814
rect 26910 34738 26962 34750
rect 27806 34802 27858 34814
rect 27806 34738 27858 34750
rect 28142 34802 28194 34814
rect 28142 34738 28194 34750
rect 29598 34802 29650 34814
rect 29598 34738 29650 34750
rect 30830 34802 30882 34814
rect 30830 34738 30882 34750
rect 31838 34802 31890 34814
rect 31838 34738 31890 34750
rect 32174 34802 32226 34814
rect 32174 34738 32226 34750
rect 33630 34802 33682 34814
rect 33630 34738 33682 34750
rect 33966 34802 34018 34814
rect 33966 34738 34018 34750
rect 34526 34802 34578 34814
rect 34526 34738 34578 34750
rect 35534 34802 35586 34814
rect 35534 34738 35586 34750
rect 35870 34802 35922 34814
rect 35870 34738 35922 34750
rect 39118 34802 39170 34814
rect 39118 34738 39170 34750
rect 39454 34802 39506 34814
rect 39454 34738 39506 34750
rect 40910 34802 40962 34814
rect 40910 34738 40962 34750
rect 41246 34802 41298 34814
rect 41246 34738 41298 34750
rect 47742 34802 47794 34814
rect 47742 34738 47794 34750
rect 48638 34802 48690 34814
rect 48638 34738 48690 34750
rect 48974 34802 49026 34814
rect 48974 34738 49026 34750
rect 51438 34802 51490 34814
rect 51438 34738 51490 34750
rect 51774 34802 51826 34814
rect 51774 34738 51826 34750
rect 52334 34802 52386 34814
rect 52334 34738 52386 34750
rect 54014 34802 54066 34814
rect 54014 34738 54066 34750
rect 56478 34802 56530 34814
rect 56478 34738 56530 34750
rect 60062 34802 60114 34814
rect 60062 34738 60114 34750
rect 73278 34802 73330 34814
rect 73278 34738 73330 34750
rect 84030 34802 84082 34814
rect 84030 34738 84082 34750
rect 85262 34802 85314 34814
rect 85262 34738 85314 34750
rect 85598 34802 85650 34814
rect 85598 34738 85650 34750
rect 86942 34802 86994 34814
rect 86942 34738 86994 34750
rect 87278 34802 87330 34814
rect 87278 34738 87330 34750
rect 92430 34802 92482 34814
rect 92430 34738 92482 34750
rect 102398 34802 102450 34814
rect 102398 34738 102450 34750
rect 102958 34802 103010 34814
rect 102958 34738 103010 34750
rect 103294 34802 103346 34814
rect 103294 34738 103346 34750
rect 111470 34802 111522 34814
rect 111470 34738 111522 34750
rect 113150 34802 113202 34814
rect 113150 34738 113202 34750
rect 114382 34802 114434 34814
rect 114382 34738 114434 34750
rect 115838 34802 115890 34814
rect 115838 34738 115890 34750
rect 118750 34802 118802 34814
rect 118750 34738 118802 34750
rect 119086 34802 119138 34814
rect 119086 34738 119138 34750
rect 121550 34802 121602 34814
rect 121550 34738 121602 34750
rect 121886 34802 121938 34814
rect 121886 34738 121938 34750
rect 122446 34802 122498 34814
rect 122446 34738 122498 34750
rect 123342 34802 123394 34814
rect 123342 34738 123394 34750
rect 123678 34802 123730 34814
rect 123678 34738 123730 34750
rect 126254 34802 126306 34814
rect 126254 34738 126306 34750
rect 127710 34802 127762 34814
rect 127710 34738 127762 34750
rect 128046 34802 128098 34814
rect 128046 34738 128098 34750
rect 132974 34802 133026 34814
rect 132974 34738 133026 34750
rect 134430 34802 134482 34814
rect 134430 34738 134482 34750
rect 139806 34802 139858 34814
rect 139806 34738 139858 34750
rect 141262 34802 141314 34814
rect 141262 34738 141314 34750
rect 142158 34802 142210 34814
rect 142158 34738 142210 34750
rect 142494 34802 142546 34814
rect 142494 34738 142546 34750
rect 142942 34802 142994 34814
rect 142942 34738 142994 34750
rect 15486 34690 15538 34702
rect 15486 34626 15538 34638
rect 28702 34690 28754 34702
rect 28702 34626 28754 34638
rect 33070 34690 33122 34702
rect 33070 34626 33122 34638
rect 34862 34690 34914 34702
rect 34862 34626 34914 34638
rect 36766 34690 36818 34702
rect 36766 34626 36818 34638
rect 38558 34690 38610 34702
rect 38558 34626 38610 34638
rect 40350 34690 40402 34702
rect 40350 34626 40402 34638
rect 42814 34690 42866 34702
rect 42814 34626 42866 34638
rect 44606 34690 44658 34702
rect 44606 34626 44658 34638
rect 47294 34690 47346 34702
rect 47294 34626 47346 34638
rect 48078 34690 48130 34702
rect 48078 34626 48130 34638
rect 49870 34690 49922 34702
rect 49870 34626 49922 34638
rect 50878 34690 50930 34702
rect 50878 34626 50930 34638
rect 52670 34690 52722 34702
rect 52670 34626 52722 34638
rect 55358 34690 55410 34702
rect 55358 34626 55410 34638
rect 56814 34690 56866 34702
rect 56814 34626 56866 34638
rect 57710 34690 57762 34702
rect 57710 34626 57762 34638
rect 58942 34690 58994 34702
rect 58942 34626 58994 34638
rect 60622 34690 60674 34702
rect 60622 34626 60674 34638
rect 61630 34690 61682 34702
rect 61630 34626 61682 34638
rect 62526 34690 62578 34702
rect 62526 34626 62578 34638
rect 67902 34690 67954 34702
rect 67902 34626 67954 34638
rect 69694 34690 69746 34702
rect 69694 34626 69746 34638
rect 74174 34690 74226 34702
rect 74174 34626 74226 34638
rect 75294 34690 75346 34702
rect 75294 34626 75346 34638
rect 75966 34690 76018 34702
rect 75966 34626 76018 34638
rect 76638 34690 76690 34702
rect 76638 34626 76690 34638
rect 79774 34690 79826 34702
rect 79774 34626 79826 34638
rect 80222 34690 80274 34702
rect 80222 34626 80274 34638
rect 80670 34690 80722 34702
rect 80670 34626 80722 34638
rect 81342 34690 81394 34702
rect 81342 34626 81394 34638
rect 83694 34690 83746 34702
rect 83694 34626 83746 34638
rect 84590 34690 84642 34702
rect 84590 34626 84642 34638
rect 86158 34690 86210 34702
rect 86158 34626 86210 34638
rect 92094 34690 92146 34702
rect 92094 34626 92146 34638
rect 97134 34690 97186 34702
rect 97134 34626 97186 34638
rect 98030 34690 98082 34702
rect 98030 34626 98082 34638
rect 98366 34690 98418 34702
rect 98366 34626 98418 34638
rect 101166 34690 101218 34702
rect 101166 34626 101218 34638
rect 101614 34690 101666 34702
rect 101614 34626 101666 34638
rect 102062 34690 102114 34702
rect 102062 34626 102114 34638
rect 104302 34690 104354 34702
rect 104302 34626 104354 34638
rect 110798 34690 110850 34702
rect 110798 34626 110850 34638
rect 112254 34690 112306 34702
rect 112254 34626 112306 34638
rect 113486 34690 113538 34702
rect 113486 34626 113538 34638
rect 114046 34690 114098 34702
rect 114046 34626 114098 34638
rect 115054 34690 115106 34702
rect 115054 34626 115106 34638
rect 116286 34690 116338 34702
rect 116286 34626 116338 34638
rect 118190 34690 118242 34702
rect 118190 34626 118242 34638
rect 119646 34690 119698 34702
rect 119646 34626 119698 34638
rect 124238 34690 124290 34702
rect 124238 34626 124290 34638
rect 125022 34690 125074 34702
rect 125022 34626 125074 34638
rect 125918 34690 125970 34702
rect 125918 34626 125970 34638
rect 126814 34690 126866 34702
rect 126814 34626 126866 34638
rect 128606 34690 128658 34702
rect 128606 34626 128658 34638
rect 133758 34690 133810 34702
rect 133758 34626 133810 34638
rect 134766 34690 134818 34702
rect 134766 34626 134818 34638
rect 143726 34690 143778 34702
rect 143726 34626 143778 34638
rect 1344 34522 148784 34556
rect 1344 34470 38034 34522
rect 38086 34470 38138 34522
rect 38190 34470 38242 34522
rect 38294 34470 74854 34522
rect 74906 34470 74958 34522
rect 75010 34470 75062 34522
rect 75114 34470 111674 34522
rect 111726 34470 111778 34522
rect 111830 34470 111882 34522
rect 111934 34470 148494 34522
rect 148546 34470 148598 34522
rect 148650 34470 148702 34522
rect 148754 34470 148784 34522
rect 1344 34436 148784 34470
rect 7534 34354 7586 34366
rect 7534 34290 7586 34302
rect 7982 34354 8034 34366
rect 7982 34290 8034 34302
rect 9662 34354 9714 34366
rect 9662 34290 9714 34302
rect 12238 34354 12290 34366
rect 12238 34290 12290 34302
rect 14814 34354 14866 34366
rect 14814 34290 14866 34302
rect 15710 34354 15762 34366
rect 15710 34290 15762 34302
rect 18062 34354 18114 34366
rect 18062 34290 18114 34302
rect 19518 34354 19570 34366
rect 19518 34290 19570 34302
rect 20974 34354 21026 34366
rect 20974 34290 21026 34302
rect 22878 34354 22930 34366
rect 22878 34290 22930 34302
rect 23326 34354 23378 34366
rect 23326 34290 23378 34302
rect 24222 34354 24274 34366
rect 24222 34290 24274 34302
rect 26014 34354 26066 34366
rect 26014 34290 26066 34302
rect 27694 34354 27746 34366
rect 27694 34290 27746 34302
rect 28478 34354 28530 34366
rect 28478 34290 28530 34302
rect 29038 34354 29090 34366
rect 29038 34290 29090 34302
rect 29374 34354 29426 34366
rect 29374 34290 29426 34302
rect 29822 34354 29874 34366
rect 29822 34290 29874 34302
rect 30382 34354 30434 34366
rect 30382 34290 30434 34302
rect 31726 34354 31778 34366
rect 31726 34290 31778 34302
rect 33518 34354 33570 34366
rect 33518 34290 33570 34302
rect 36878 34354 36930 34366
rect 36878 34290 36930 34302
rect 37438 34354 37490 34366
rect 37438 34290 37490 34302
rect 40574 34354 40626 34366
rect 40574 34290 40626 34302
rect 46622 34354 46674 34366
rect 46622 34290 46674 34302
rect 48862 34354 48914 34366
rect 48862 34290 48914 34302
rect 49982 34354 50034 34366
rect 49982 34290 50034 34302
rect 50878 34354 50930 34366
rect 50878 34290 50930 34302
rect 51662 34354 51714 34366
rect 51662 34290 51714 34302
rect 52222 34354 52274 34366
rect 52222 34290 52274 34302
rect 54238 34354 54290 34366
rect 54238 34290 54290 34302
rect 54798 34354 54850 34366
rect 54798 34290 54850 34302
rect 56590 34354 56642 34366
rect 56590 34290 56642 34302
rect 57486 34354 57538 34366
rect 57486 34290 57538 34302
rect 58382 34354 58434 34366
rect 58382 34290 58434 34302
rect 59278 34354 59330 34366
rect 59278 34290 59330 34302
rect 62638 34354 62690 34366
rect 62638 34290 62690 34302
rect 63870 34354 63922 34366
rect 63870 34290 63922 34302
rect 64654 34354 64706 34366
rect 64654 34290 64706 34302
rect 65438 34354 65490 34366
rect 65438 34290 65490 34302
rect 67902 34354 67954 34366
rect 67902 34290 67954 34302
rect 73278 34354 73330 34366
rect 73278 34290 73330 34302
rect 73950 34354 74002 34366
rect 73950 34290 74002 34302
rect 74398 34354 74450 34366
rect 74398 34290 74450 34302
rect 75182 34354 75234 34366
rect 75182 34290 75234 34302
rect 75630 34354 75682 34366
rect 75630 34290 75682 34302
rect 76190 34354 76242 34366
rect 76190 34290 76242 34302
rect 76750 34354 76802 34366
rect 76750 34290 76802 34302
rect 78206 34354 78258 34366
rect 78206 34290 78258 34302
rect 78766 34354 78818 34366
rect 78766 34290 78818 34302
rect 81342 34354 81394 34366
rect 81342 34290 81394 34302
rect 81790 34354 81842 34366
rect 81790 34290 81842 34302
rect 82350 34354 82402 34366
rect 82350 34290 82402 34302
rect 83918 34354 83970 34366
rect 83918 34290 83970 34302
rect 84366 34354 84418 34366
rect 84366 34290 84418 34302
rect 86158 34354 86210 34366
rect 86158 34290 86210 34302
rect 87390 34354 87442 34366
rect 87390 34290 87442 34302
rect 87950 34354 88002 34366
rect 87950 34290 88002 34302
rect 89294 34354 89346 34366
rect 89294 34290 89346 34302
rect 90862 34354 90914 34366
rect 90862 34290 90914 34302
rect 93438 34354 93490 34366
rect 93438 34290 93490 34302
rect 95566 34354 95618 34366
rect 95566 34290 95618 34302
rect 96350 34354 96402 34366
rect 96350 34290 96402 34302
rect 97246 34354 97298 34366
rect 97246 34290 97298 34302
rect 103518 34354 103570 34366
rect 103518 34290 103570 34302
rect 105646 34354 105698 34366
rect 105646 34290 105698 34302
rect 107326 34354 107378 34366
rect 107326 34290 107378 34302
rect 108782 34354 108834 34366
rect 108782 34290 108834 34302
rect 109230 34354 109282 34366
rect 109230 34290 109282 34302
rect 111246 34354 111298 34366
rect 111246 34290 111298 34302
rect 114942 34354 114994 34366
rect 114942 34290 114994 34302
rect 117518 34354 117570 34366
rect 117518 34290 117570 34302
rect 122670 34354 122722 34366
rect 122670 34290 122722 34302
rect 123006 34354 123058 34366
rect 123006 34290 123058 34302
rect 124798 34354 124850 34366
rect 124798 34290 124850 34302
rect 125134 34354 125186 34366
rect 125134 34290 125186 34302
rect 127822 34354 127874 34366
rect 127822 34290 127874 34302
rect 129390 34354 129442 34366
rect 129390 34290 129442 34302
rect 130286 34354 130338 34366
rect 130286 34290 130338 34302
rect 131742 34354 131794 34366
rect 131742 34290 131794 34302
rect 132526 34354 132578 34366
rect 132526 34290 132578 34302
rect 132974 34354 133026 34366
rect 132974 34290 133026 34302
rect 135214 34354 135266 34366
rect 135214 34290 135266 34302
rect 135662 34354 135714 34366
rect 135662 34290 135714 34302
rect 137342 34354 137394 34366
rect 137342 34290 137394 34302
rect 138910 34354 138962 34366
rect 138910 34290 138962 34302
rect 139358 34354 139410 34366
rect 139358 34290 139410 34302
rect 140366 34354 140418 34366
rect 140366 34290 140418 34302
rect 140814 34354 140866 34366
rect 140814 34290 140866 34302
rect 141486 34354 141538 34366
rect 141486 34290 141538 34302
rect 141934 34354 141986 34366
rect 141934 34290 141986 34302
rect 143502 34354 143554 34366
rect 143502 34290 143554 34302
rect 8430 34242 8482 34254
rect 8430 34178 8482 34190
rect 8766 34242 8818 34254
rect 8766 34178 8818 34190
rect 19182 34242 19234 34254
rect 19182 34178 19234 34190
rect 20078 34242 20130 34254
rect 20078 34178 20130 34190
rect 20414 34242 20466 34254
rect 20414 34178 20466 34190
rect 28142 34242 28194 34254
rect 28142 34178 28194 34190
rect 30830 34242 30882 34254
rect 30830 34178 30882 34190
rect 31166 34242 31218 34254
rect 31166 34178 31218 34190
rect 39454 34242 39506 34254
rect 39454 34178 39506 34190
rect 46062 34242 46114 34254
rect 46062 34178 46114 34190
rect 49646 34242 49698 34254
rect 49646 34178 49698 34190
rect 52558 34242 52610 34254
rect 52558 34178 52610 34190
rect 53118 34242 53170 34254
rect 53118 34178 53170 34190
rect 53454 34242 53506 34254
rect 53454 34178 53506 34190
rect 73838 34242 73890 34254
rect 73838 34178 73890 34190
rect 79214 34242 79266 34254
rect 79214 34178 79266 34190
rect 82798 34242 82850 34254
rect 82798 34178 82850 34190
rect 83134 34242 83186 34254
rect 83134 34178 83186 34190
rect 89854 34242 89906 34254
rect 106094 34242 106146 34254
rect 92642 34190 92654 34242
rect 92706 34190 92718 34242
rect 89854 34178 89906 34190
rect 106094 34178 106146 34190
rect 106430 34242 106482 34254
rect 106430 34178 106482 34190
rect 107886 34242 107938 34254
rect 107886 34178 107938 34190
rect 109678 34242 109730 34254
rect 109678 34178 109730 34190
rect 113598 34242 113650 34254
rect 113598 34178 113650 34190
rect 126142 34242 126194 34254
rect 126142 34178 126194 34190
rect 130846 34242 130898 34254
rect 130846 34178 130898 34190
rect 131182 34242 131234 34254
rect 131182 34178 131234 34190
rect 132078 34242 132130 34254
rect 132078 34178 132130 34190
rect 138350 34242 138402 34254
rect 138350 34178 138402 34190
rect 142270 34242 142322 34254
rect 142270 34178 142322 34190
rect 18398 34130 18450 34142
rect 18398 34066 18450 34078
rect 21310 34130 21362 34142
rect 21310 34066 21362 34078
rect 25566 34130 25618 34142
rect 25566 34066 25618 34078
rect 37774 34130 37826 34142
rect 37774 34066 37826 34078
rect 39118 34130 39170 34142
rect 39118 34066 39170 34078
rect 44718 34130 44770 34142
rect 46958 34130 47010 34142
rect 45826 34078 45838 34130
rect 45890 34078 45902 34130
rect 44718 34066 44770 34078
rect 46958 34066 47010 34078
rect 48190 34130 48242 34142
rect 48190 34066 48242 34078
rect 61182 34130 61234 34142
rect 61182 34066 61234 34078
rect 62302 34130 62354 34142
rect 106990 34130 107042 34142
rect 113934 34130 113986 34142
rect 79426 34078 79438 34130
rect 79490 34078 79502 34130
rect 91746 34078 91758 34130
rect 91810 34078 91822 34130
rect 108098 34078 108110 34130
rect 108162 34078 108174 34130
rect 109890 34078 109902 34130
rect 109954 34078 109966 34130
rect 62302 34066 62354 34078
rect 106990 34066 107042 34078
rect 113934 34066 113986 34078
rect 125582 34130 125634 34142
rect 125582 34066 125634 34078
rect 126478 34130 126530 34142
rect 126478 34066 126530 34078
rect 129054 34130 129106 34142
rect 130050 34078 130062 34130
rect 130114 34078 130126 34130
rect 129054 34066 129106 34078
rect 13470 34018 13522 34030
rect 13470 33954 13522 33966
rect 16494 34018 16546 34030
rect 16494 33954 16546 33966
rect 17054 34018 17106 34030
rect 17054 33954 17106 33966
rect 21758 34018 21810 34030
rect 21758 33954 21810 33966
rect 22430 34018 22482 34030
rect 22430 33954 22482 33966
rect 27134 34018 27186 34030
rect 27134 33954 27186 33966
rect 32398 34018 32450 34030
rect 32398 33954 32450 33966
rect 34190 34018 34242 34030
rect 34190 33954 34242 33966
rect 35086 34018 35138 34030
rect 35086 33954 35138 33966
rect 36094 34018 36146 34030
rect 36094 33954 36146 33966
rect 38558 34018 38610 34030
rect 38558 33954 38610 33966
rect 39902 34018 39954 34030
rect 39902 33954 39954 33966
rect 41470 34018 41522 34030
rect 41470 33954 41522 33966
rect 41918 34018 41970 34030
rect 41918 33954 41970 33966
rect 42926 34018 42978 34030
rect 42926 33954 42978 33966
rect 45278 34018 45330 34030
rect 45278 33954 45330 33966
rect 47406 34018 47458 34030
rect 47406 33954 47458 33966
rect 51214 34018 51266 34030
rect 51214 33954 51266 33966
rect 55134 34018 55186 34030
rect 55134 33954 55186 33966
rect 55806 34018 55858 34030
rect 55806 33954 55858 33966
rect 56142 34018 56194 34030
rect 56142 33954 56194 33966
rect 57822 34018 57874 34030
rect 57822 33954 57874 33966
rect 58718 34018 58770 34030
rect 58718 33954 58770 33966
rect 59838 34018 59890 34030
rect 59838 33954 59890 33966
rect 60174 34018 60226 34030
rect 60174 33954 60226 33966
rect 60622 34018 60674 34030
rect 60622 33954 60674 33966
rect 61742 34018 61794 34030
rect 61742 33954 61794 33966
rect 63310 34018 63362 34030
rect 63310 33954 63362 33966
rect 65886 34018 65938 34030
rect 65886 33954 65938 33966
rect 66446 34018 66498 34030
rect 66446 33954 66498 33966
rect 67454 34018 67506 34030
rect 67454 33954 67506 33966
rect 69022 34018 69074 34030
rect 69022 33954 69074 33966
rect 72718 34018 72770 34030
rect 72718 33954 72770 33966
rect 77198 34018 77250 34030
rect 77198 33954 77250 33966
rect 86606 34018 86658 34030
rect 86606 33954 86658 33966
rect 88510 34018 88562 34030
rect 88510 33954 88562 33966
rect 90302 34018 90354 34030
rect 90302 33954 90354 33966
rect 91198 34018 91250 34030
rect 91198 33954 91250 33966
rect 93886 34018 93938 34030
rect 93886 33954 93938 33966
rect 95118 34018 95170 34030
rect 95118 33954 95170 33966
rect 96014 34018 96066 34030
rect 96014 33954 96066 33966
rect 102622 34018 102674 34030
rect 102622 33954 102674 33966
rect 104414 34018 104466 34030
rect 104414 33954 104466 33966
rect 105198 34018 105250 34030
rect 105198 33954 105250 33966
rect 110798 34018 110850 34030
rect 110798 33954 110850 33966
rect 111582 34018 111634 34030
rect 111582 33954 111634 33966
rect 113038 34018 113090 34030
rect 113038 33954 113090 33966
rect 114382 34018 114434 34030
rect 114382 33954 114434 33966
rect 119310 34018 119362 34030
rect 119310 33954 119362 33966
rect 122110 34018 122162 34030
rect 122110 33954 122162 33966
rect 123566 34018 123618 34030
rect 123566 33954 123618 33966
rect 126926 34018 126978 34030
rect 126926 33954 126978 33966
rect 127374 34018 127426 34030
rect 127374 33954 127426 33966
rect 128270 34018 128322 34030
rect 128270 33954 128322 33966
rect 134094 34018 134146 34030
rect 134094 33954 134146 33966
rect 138014 34018 138066 34030
rect 138014 33954 138066 33966
rect 139918 34018 139970 34030
rect 139918 33954 139970 33966
rect 138002 33854 138014 33906
rect 138066 33903 138078 33906
rect 138674 33903 138686 33906
rect 138066 33857 138686 33903
rect 138066 33854 138078 33857
rect 138674 33854 138686 33857
rect 138738 33854 138750 33906
rect 139906 33854 139918 33906
rect 139970 33903 139982 33906
rect 140578 33903 140590 33906
rect 139970 33857 140590 33903
rect 139970 33854 139982 33857
rect 140578 33854 140590 33857
rect 140642 33854 140654 33906
rect 1344 33738 148624 33772
rect 1344 33686 19624 33738
rect 19676 33686 19728 33738
rect 19780 33686 19832 33738
rect 19884 33686 56444 33738
rect 56496 33686 56548 33738
rect 56600 33686 56652 33738
rect 56704 33686 93264 33738
rect 93316 33686 93368 33738
rect 93420 33686 93472 33738
rect 93524 33686 130084 33738
rect 130136 33686 130188 33738
rect 130240 33686 130292 33738
rect 130344 33686 148624 33738
rect 1344 33652 148624 33686
rect 106642 33518 106654 33570
rect 106706 33567 106718 33570
rect 106978 33567 106990 33570
rect 106706 33521 106990 33567
rect 106706 33518 106718 33521
rect 106978 33518 106990 33521
rect 107042 33518 107054 33570
rect 17502 33458 17554 33470
rect 17502 33394 17554 33406
rect 18958 33458 19010 33470
rect 18958 33394 19010 33406
rect 19294 33458 19346 33470
rect 19294 33394 19346 33406
rect 19854 33458 19906 33470
rect 19854 33394 19906 33406
rect 20638 33458 20690 33470
rect 20638 33394 20690 33406
rect 30606 33458 30658 33470
rect 30606 33394 30658 33406
rect 31054 33458 31106 33470
rect 31054 33394 31106 33406
rect 46286 33458 46338 33470
rect 46286 33394 46338 33406
rect 46846 33458 46898 33470
rect 46846 33394 46898 33406
rect 49198 33458 49250 33470
rect 49198 33394 49250 33406
rect 51998 33458 52050 33470
rect 51998 33394 52050 33406
rect 53342 33458 53394 33470
rect 53342 33394 53394 33406
rect 53902 33458 53954 33470
rect 53902 33394 53954 33406
rect 59278 33458 59330 33470
rect 59278 33394 59330 33406
rect 60286 33458 60338 33470
rect 60286 33394 60338 33406
rect 61742 33458 61794 33470
rect 61742 33394 61794 33406
rect 63086 33458 63138 33470
rect 63086 33394 63138 33406
rect 64542 33458 64594 33470
rect 64542 33394 64594 33406
rect 65102 33458 65154 33470
rect 65102 33394 65154 33406
rect 65550 33458 65602 33470
rect 65550 33394 65602 33406
rect 73838 33458 73890 33470
rect 73838 33394 73890 33406
rect 74286 33458 74338 33470
rect 74286 33394 74338 33406
rect 74622 33458 74674 33470
rect 74622 33394 74674 33406
rect 87950 33458 88002 33470
rect 87950 33394 88002 33406
rect 89070 33458 89122 33470
rect 89070 33394 89122 33406
rect 91758 33458 91810 33470
rect 91758 33394 91810 33406
rect 93214 33458 93266 33470
rect 93214 33394 93266 33406
rect 105758 33458 105810 33470
rect 105758 33394 105810 33406
rect 106206 33458 106258 33470
rect 106206 33394 106258 33406
rect 107214 33458 107266 33470
rect 107214 33394 107266 33406
rect 107662 33458 107714 33470
rect 107662 33394 107714 33406
rect 109454 33458 109506 33470
rect 109454 33394 109506 33406
rect 110126 33458 110178 33470
rect 110126 33394 110178 33406
rect 126590 33458 126642 33470
rect 126590 33394 126642 33406
rect 127038 33458 127090 33470
rect 127038 33394 127090 33406
rect 128718 33458 128770 33470
rect 128718 33394 128770 33406
rect 131070 33458 131122 33470
rect 131070 33394 131122 33406
rect 131518 33458 131570 33470
rect 131518 33394 131570 33406
rect 51550 33346 51602 33358
rect 51550 33282 51602 33294
rect 52782 33346 52834 33358
rect 52782 33282 52834 33294
rect 54462 33346 54514 33358
rect 54462 33282 54514 33294
rect 62190 33346 62242 33358
rect 62190 33282 62242 33294
rect 63758 33346 63810 33358
rect 63758 33282 63810 33294
rect 129278 33346 129330 33358
rect 129278 33282 129330 33294
rect 18398 33234 18450 33246
rect 18398 33170 18450 33182
rect 89518 33234 89570 33246
rect 89518 33170 89570 33182
rect 110910 33234 110962 33246
rect 110910 33170 110962 33182
rect 129614 33234 129666 33246
rect 129614 33170 129666 33182
rect 20302 33122 20354 33134
rect 20302 33058 20354 33070
rect 37998 33122 38050 33134
rect 37998 33058 38050 33070
rect 38446 33122 38498 33134
rect 38446 33058 38498 33070
rect 60622 33122 60674 33134
rect 60622 33058 60674 33070
rect 62526 33122 62578 33134
rect 62526 33058 62578 33070
rect 64206 33122 64258 33134
rect 64206 33058 64258 33070
rect 76078 33122 76130 33134
rect 76078 33058 76130 33070
rect 105086 33122 105138 33134
rect 105086 33058 105138 33070
rect 106654 33122 106706 33134
rect 106654 33058 106706 33070
rect 107998 33122 108050 33134
rect 107998 33058 108050 33070
rect 109118 33122 109170 33134
rect 109118 33058 109170 33070
rect 130174 33122 130226 33134
rect 130174 33058 130226 33070
rect 130510 33122 130562 33134
rect 130510 33058 130562 33070
rect 1344 32954 148784 32988
rect 1344 32902 38034 32954
rect 38086 32902 38138 32954
rect 38190 32902 38242 32954
rect 38294 32902 74854 32954
rect 74906 32902 74958 32954
rect 75010 32902 75062 32954
rect 75114 32902 111674 32954
rect 111726 32902 111778 32954
rect 111830 32902 111882 32954
rect 111934 32902 148494 32954
rect 148546 32902 148598 32954
rect 148650 32902 148702 32954
rect 148754 32902 148784 32954
rect 1344 32868 148784 32902
rect 53454 32786 53506 32798
rect 53454 32722 53506 32734
rect 62078 32786 62130 32798
rect 62078 32722 62130 32734
rect 62526 32786 62578 32798
rect 62526 32722 62578 32734
rect 62974 32786 63026 32798
rect 62974 32722 63026 32734
rect 108222 32786 108274 32798
rect 108222 32722 108274 32734
rect 1344 32170 148624 32204
rect 1344 32118 19624 32170
rect 19676 32118 19728 32170
rect 19780 32118 19832 32170
rect 19884 32118 56444 32170
rect 56496 32118 56548 32170
rect 56600 32118 56652 32170
rect 56704 32118 93264 32170
rect 93316 32118 93368 32170
rect 93420 32118 93472 32170
rect 93524 32118 130084 32170
rect 130136 32118 130188 32170
rect 130240 32118 130292 32170
rect 130344 32118 148624 32170
rect 1344 32084 148624 32118
rect 1344 31386 148784 31420
rect 1344 31334 38034 31386
rect 38086 31334 38138 31386
rect 38190 31334 38242 31386
rect 38294 31334 74854 31386
rect 74906 31334 74958 31386
rect 75010 31334 75062 31386
rect 75114 31334 111674 31386
rect 111726 31334 111778 31386
rect 111830 31334 111882 31386
rect 111934 31334 148494 31386
rect 148546 31334 148598 31386
rect 148650 31334 148702 31386
rect 148754 31334 148784 31386
rect 1344 31300 148784 31334
rect 1344 30602 148624 30636
rect 1344 30550 19624 30602
rect 19676 30550 19728 30602
rect 19780 30550 19832 30602
rect 19884 30550 56444 30602
rect 56496 30550 56548 30602
rect 56600 30550 56652 30602
rect 56704 30550 93264 30602
rect 93316 30550 93368 30602
rect 93420 30550 93472 30602
rect 93524 30550 130084 30602
rect 130136 30550 130188 30602
rect 130240 30550 130292 30602
rect 130344 30550 148624 30602
rect 1344 30516 148624 30550
rect 1344 29818 148784 29852
rect 1344 29766 38034 29818
rect 38086 29766 38138 29818
rect 38190 29766 38242 29818
rect 38294 29766 74854 29818
rect 74906 29766 74958 29818
rect 75010 29766 75062 29818
rect 75114 29766 111674 29818
rect 111726 29766 111778 29818
rect 111830 29766 111882 29818
rect 111934 29766 148494 29818
rect 148546 29766 148598 29818
rect 148650 29766 148702 29818
rect 148754 29766 148784 29818
rect 1344 29732 148784 29766
rect 1344 29034 148624 29068
rect 1344 28982 19624 29034
rect 19676 28982 19728 29034
rect 19780 28982 19832 29034
rect 19884 28982 56444 29034
rect 56496 28982 56548 29034
rect 56600 28982 56652 29034
rect 56704 28982 93264 29034
rect 93316 28982 93368 29034
rect 93420 28982 93472 29034
rect 93524 28982 130084 29034
rect 130136 28982 130188 29034
rect 130240 28982 130292 29034
rect 130344 28982 148624 29034
rect 1344 28948 148624 28982
rect 1344 28250 148784 28284
rect 1344 28198 38034 28250
rect 38086 28198 38138 28250
rect 38190 28198 38242 28250
rect 38294 28198 74854 28250
rect 74906 28198 74958 28250
rect 75010 28198 75062 28250
rect 75114 28198 111674 28250
rect 111726 28198 111778 28250
rect 111830 28198 111882 28250
rect 111934 28198 148494 28250
rect 148546 28198 148598 28250
rect 148650 28198 148702 28250
rect 148754 28198 148784 28250
rect 1344 28164 148784 28198
rect 1344 27466 148624 27500
rect 1344 27414 19624 27466
rect 19676 27414 19728 27466
rect 19780 27414 19832 27466
rect 19884 27414 56444 27466
rect 56496 27414 56548 27466
rect 56600 27414 56652 27466
rect 56704 27414 93264 27466
rect 93316 27414 93368 27466
rect 93420 27414 93472 27466
rect 93524 27414 130084 27466
rect 130136 27414 130188 27466
rect 130240 27414 130292 27466
rect 130344 27414 148624 27466
rect 1344 27380 148624 27414
rect 1344 26682 148784 26716
rect 1344 26630 38034 26682
rect 38086 26630 38138 26682
rect 38190 26630 38242 26682
rect 38294 26630 74854 26682
rect 74906 26630 74958 26682
rect 75010 26630 75062 26682
rect 75114 26630 111674 26682
rect 111726 26630 111778 26682
rect 111830 26630 111882 26682
rect 111934 26630 148494 26682
rect 148546 26630 148598 26682
rect 148650 26630 148702 26682
rect 148754 26630 148784 26682
rect 1344 26596 148784 26630
rect 1344 25898 148624 25932
rect 1344 25846 19624 25898
rect 19676 25846 19728 25898
rect 19780 25846 19832 25898
rect 19884 25846 56444 25898
rect 56496 25846 56548 25898
rect 56600 25846 56652 25898
rect 56704 25846 93264 25898
rect 93316 25846 93368 25898
rect 93420 25846 93472 25898
rect 93524 25846 130084 25898
rect 130136 25846 130188 25898
rect 130240 25846 130292 25898
rect 130344 25846 148624 25898
rect 1344 25812 148624 25846
rect 1344 25114 148784 25148
rect 1344 25062 38034 25114
rect 38086 25062 38138 25114
rect 38190 25062 38242 25114
rect 38294 25062 74854 25114
rect 74906 25062 74958 25114
rect 75010 25062 75062 25114
rect 75114 25062 111674 25114
rect 111726 25062 111778 25114
rect 111830 25062 111882 25114
rect 111934 25062 148494 25114
rect 148546 25062 148598 25114
rect 148650 25062 148702 25114
rect 148754 25062 148784 25114
rect 1344 25028 148784 25062
rect 1344 24330 148624 24364
rect 1344 24278 19624 24330
rect 19676 24278 19728 24330
rect 19780 24278 19832 24330
rect 19884 24278 56444 24330
rect 56496 24278 56548 24330
rect 56600 24278 56652 24330
rect 56704 24278 93264 24330
rect 93316 24278 93368 24330
rect 93420 24278 93472 24330
rect 93524 24278 130084 24330
rect 130136 24278 130188 24330
rect 130240 24278 130292 24330
rect 130344 24278 148624 24330
rect 1344 24244 148624 24278
rect 1344 23546 148784 23580
rect 1344 23494 38034 23546
rect 38086 23494 38138 23546
rect 38190 23494 38242 23546
rect 38294 23494 74854 23546
rect 74906 23494 74958 23546
rect 75010 23494 75062 23546
rect 75114 23494 111674 23546
rect 111726 23494 111778 23546
rect 111830 23494 111882 23546
rect 111934 23494 148494 23546
rect 148546 23494 148598 23546
rect 148650 23494 148702 23546
rect 148754 23494 148784 23546
rect 1344 23460 148784 23494
rect 1344 22762 148624 22796
rect 1344 22710 19624 22762
rect 19676 22710 19728 22762
rect 19780 22710 19832 22762
rect 19884 22710 56444 22762
rect 56496 22710 56548 22762
rect 56600 22710 56652 22762
rect 56704 22710 93264 22762
rect 93316 22710 93368 22762
rect 93420 22710 93472 22762
rect 93524 22710 130084 22762
rect 130136 22710 130188 22762
rect 130240 22710 130292 22762
rect 130344 22710 148624 22762
rect 1344 22676 148624 22710
rect 1344 21978 148784 22012
rect 1344 21926 38034 21978
rect 38086 21926 38138 21978
rect 38190 21926 38242 21978
rect 38294 21926 74854 21978
rect 74906 21926 74958 21978
rect 75010 21926 75062 21978
rect 75114 21926 111674 21978
rect 111726 21926 111778 21978
rect 111830 21926 111882 21978
rect 111934 21926 148494 21978
rect 148546 21926 148598 21978
rect 148650 21926 148702 21978
rect 148754 21926 148784 21978
rect 1344 21892 148784 21926
rect 1344 21194 148624 21228
rect 1344 21142 19624 21194
rect 19676 21142 19728 21194
rect 19780 21142 19832 21194
rect 19884 21142 56444 21194
rect 56496 21142 56548 21194
rect 56600 21142 56652 21194
rect 56704 21142 93264 21194
rect 93316 21142 93368 21194
rect 93420 21142 93472 21194
rect 93524 21142 130084 21194
rect 130136 21142 130188 21194
rect 130240 21142 130292 21194
rect 130344 21142 148624 21194
rect 1344 21108 148624 21142
rect 1344 20410 148784 20444
rect 1344 20358 38034 20410
rect 38086 20358 38138 20410
rect 38190 20358 38242 20410
rect 38294 20358 74854 20410
rect 74906 20358 74958 20410
rect 75010 20358 75062 20410
rect 75114 20358 111674 20410
rect 111726 20358 111778 20410
rect 111830 20358 111882 20410
rect 111934 20358 148494 20410
rect 148546 20358 148598 20410
rect 148650 20358 148702 20410
rect 148754 20358 148784 20410
rect 1344 20324 148784 20358
rect 1344 19626 148624 19660
rect 1344 19574 19624 19626
rect 19676 19574 19728 19626
rect 19780 19574 19832 19626
rect 19884 19574 56444 19626
rect 56496 19574 56548 19626
rect 56600 19574 56652 19626
rect 56704 19574 93264 19626
rect 93316 19574 93368 19626
rect 93420 19574 93472 19626
rect 93524 19574 130084 19626
rect 130136 19574 130188 19626
rect 130240 19574 130292 19626
rect 130344 19574 148624 19626
rect 1344 19540 148624 19574
rect 1344 18842 148784 18876
rect 1344 18790 38034 18842
rect 38086 18790 38138 18842
rect 38190 18790 38242 18842
rect 38294 18790 74854 18842
rect 74906 18790 74958 18842
rect 75010 18790 75062 18842
rect 75114 18790 111674 18842
rect 111726 18790 111778 18842
rect 111830 18790 111882 18842
rect 111934 18790 148494 18842
rect 148546 18790 148598 18842
rect 148650 18790 148702 18842
rect 148754 18790 148784 18842
rect 1344 18756 148784 18790
rect 1344 18058 148624 18092
rect 1344 18006 19624 18058
rect 19676 18006 19728 18058
rect 19780 18006 19832 18058
rect 19884 18006 56444 18058
rect 56496 18006 56548 18058
rect 56600 18006 56652 18058
rect 56704 18006 93264 18058
rect 93316 18006 93368 18058
rect 93420 18006 93472 18058
rect 93524 18006 130084 18058
rect 130136 18006 130188 18058
rect 130240 18006 130292 18058
rect 130344 18006 148624 18058
rect 1344 17972 148624 18006
rect 1344 17274 148784 17308
rect 1344 17222 38034 17274
rect 38086 17222 38138 17274
rect 38190 17222 38242 17274
rect 38294 17222 74854 17274
rect 74906 17222 74958 17274
rect 75010 17222 75062 17274
rect 75114 17222 111674 17274
rect 111726 17222 111778 17274
rect 111830 17222 111882 17274
rect 111934 17222 148494 17274
rect 148546 17222 148598 17274
rect 148650 17222 148702 17274
rect 148754 17222 148784 17274
rect 1344 17188 148784 17222
rect 1344 16490 148624 16524
rect 1344 16438 19624 16490
rect 19676 16438 19728 16490
rect 19780 16438 19832 16490
rect 19884 16438 56444 16490
rect 56496 16438 56548 16490
rect 56600 16438 56652 16490
rect 56704 16438 93264 16490
rect 93316 16438 93368 16490
rect 93420 16438 93472 16490
rect 93524 16438 130084 16490
rect 130136 16438 130188 16490
rect 130240 16438 130292 16490
rect 130344 16438 148624 16490
rect 1344 16404 148624 16438
rect 1344 15706 148784 15740
rect 1344 15654 38034 15706
rect 38086 15654 38138 15706
rect 38190 15654 38242 15706
rect 38294 15654 74854 15706
rect 74906 15654 74958 15706
rect 75010 15654 75062 15706
rect 75114 15654 111674 15706
rect 111726 15654 111778 15706
rect 111830 15654 111882 15706
rect 111934 15654 148494 15706
rect 148546 15654 148598 15706
rect 148650 15654 148702 15706
rect 148754 15654 148784 15706
rect 1344 15620 148784 15654
rect 1344 14922 148624 14956
rect 1344 14870 19624 14922
rect 19676 14870 19728 14922
rect 19780 14870 19832 14922
rect 19884 14870 56444 14922
rect 56496 14870 56548 14922
rect 56600 14870 56652 14922
rect 56704 14870 93264 14922
rect 93316 14870 93368 14922
rect 93420 14870 93472 14922
rect 93524 14870 130084 14922
rect 130136 14870 130188 14922
rect 130240 14870 130292 14922
rect 130344 14870 148624 14922
rect 1344 14836 148624 14870
rect 1344 14138 148784 14172
rect 1344 14086 38034 14138
rect 38086 14086 38138 14138
rect 38190 14086 38242 14138
rect 38294 14086 74854 14138
rect 74906 14086 74958 14138
rect 75010 14086 75062 14138
rect 75114 14086 111674 14138
rect 111726 14086 111778 14138
rect 111830 14086 111882 14138
rect 111934 14086 148494 14138
rect 148546 14086 148598 14138
rect 148650 14086 148702 14138
rect 148754 14086 148784 14138
rect 1344 14052 148784 14086
rect 1344 13354 148624 13388
rect 1344 13302 19624 13354
rect 19676 13302 19728 13354
rect 19780 13302 19832 13354
rect 19884 13302 56444 13354
rect 56496 13302 56548 13354
rect 56600 13302 56652 13354
rect 56704 13302 93264 13354
rect 93316 13302 93368 13354
rect 93420 13302 93472 13354
rect 93524 13302 130084 13354
rect 130136 13302 130188 13354
rect 130240 13302 130292 13354
rect 130344 13302 148624 13354
rect 1344 13268 148624 13302
rect 1344 12570 148784 12604
rect 1344 12518 38034 12570
rect 38086 12518 38138 12570
rect 38190 12518 38242 12570
rect 38294 12518 74854 12570
rect 74906 12518 74958 12570
rect 75010 12518 75062 12570
rect 75114 12518 111674 12570
rect 111726 12518 111778 12570
rect 111830 12518 111882 12570
rect 111934 12518 148494 12570
rect 148546 12518 148598 12570
rect 148650 12518 148702 12570
rect 148754 12518 148784 12570
rect 1344 12484 148784 12518
rect 1344 11786 148624 11820
rect 1344 11734 19624 11786
rect 19676 11734 19728 11786
rect 19780 11734 19832 11786
rect 19884 11734 56444 11786
rect 56496 11734 56548 11786
rect 56600 11734 56652 11786
rect 56704 11734 93264 11786
rect 93316 11734 93368 11786
rect 93420 11734 93472 11786
rect 93524 11734 130084 11786
rect 130136 11734 130188 11786
rect 130240 11734 130292 11786
rect 130344 11734 148624 11786
rect 1344 11700 148624 11734
rect 1344 11002 148784 11036
rect 1344 10950 38034 11002
rect 38086 10950 38138 11002
rect 38190 10950 38242 11002
rect 38294 10950 74854 11002
rect 74906 10950 74958 11002
rect 75010 10950 75062 11002
rect 75114 10950 111674 11002
rect 111726 10950 111778 11002
rect 111830 10950 111882 11002
rect 111934 10950 148494 11002
rect 148546 10950 148598 11002
rect 148650 10950 148702 11002
rect 148754 10950 148784 11002
rect 1344 10916 148784 10950
rect 1344 10218 148624 10252
rect 1344 10166 19624 10218
rect 19676 10166 19728 10218
rect 19780 10166 19832 10218
rect 19884 10166 56444 10218
rect 56496 10166 56548 10218
rect 56600 10166 56652 10218
rect 56704 10166 93264 10218
rect 93316 10166 93368 10218
rect 93420 10166 93472 10218
rect 93524 10166 130084 10218
rect 130136 10166 130188 10218
rect 130240 10166 130292 10218
rect 130344 10166 148624 10218
rect 1344 10132 148624 10166
rect 64990 9602 65042 9614
rect 64990 9538 65042 9550
rect 1344 9434 148784 9468
rect 1344 9382 38034 9434
rect 38086 9382 38138 9434
rect 38190 9382 38242 9434
rect 38294 9382 74854 9434
rect 74906 9382 74958 9434
rect 75010 9382 75062 9434
rect 75114 9382 111674 9434
rect 111726 9382 111778 9434
rect 111830 9382 111882 9434
rect 111934 9382 148494 9434
rect 148546 9382 148598 9434
rect 148650 9382 148702 9434
rect 148754 9382 148784 9434
rect 1344 9348 148784 9382
rect 64542 9154 64594 9166
rect 64542 9090 64594 9102
rect 65774 9154 65826 9166
rect 124674 9102 124686 9154
rect 124738 9102 124750 9154
rect 65774 9090 65826 9102
rect 65438 9042 65490 9054
rect 124898 8990 124910 9042
rect 124962 8990 124974 9042
rect 65438 8978 65490 8990
rect 62190 8930 62242 8942
rect 62190 8866 62242 8878
rect 63086 8930 63138 8942
rect 63086 8866 63138 8878
rect 63534 8930 63586 8942
rect 63534 8866 63586 8878
rect 66334 8930 66386 8942
rect 66334 8866 66386 8878
rect 105198 8930 105250 8942
rect 105198 8866 105250 8878
rect 123118 8930 123170 8942
rect 123118 8866 123170 8878
rect 124126 8930 124178 8942
rect 124126 8866 124178 8878
rect 125470 8930 125522 8942
rect 125470 8866 125522 8878
rect 125918 8930 125970 8942
rect 125918 8866 125970 8878
rect 64654 8818 64706 8830
rect 64654 8754 64706 8766
rect 123790 8818 123842 8830
rect 123790 8754 123842 8766
rect 1344 8650 148624 8684
rect 1344 8598 19624 8650
rect 19676 8598 19728 8650
rect 19780 8598 19832 8650
rect 19884 8598 56444 8650
rect 56496 8598 56548 8650
rect 56600 8598 56652 8650
rect 56704 8598 93264 8650
rect 93316 8598 93368 8650
rect 93420 8598 93472 8650
rect 93524 8598 130084 8650
rect 130136 8598 130188 8650
rect 130240 8598 130292 8650
rect 130344 8598 148624 8650
rect 1344 8564 148624 8598
rect 64878 8482 64930 8494
rect 64878 8418 64930 8430
rect 62638 8370 62690 8382
rect 62638 8306 62690 8318
rect 121886 8370 121938 8382
rect 121886 8306 121938 8318
rect 122782 8370 122834 8382
rect 122782 8306 122834 8318
rect 124126 8370 124178 8382
rect 124126 8306 124178 8318
rect 64542 8258 64594 8270
rect 67006 8258 67058 8270
rect 63858 8206 63870 8258
rect 63922 8206 63934 8258
rect 65986 8206 65998 8258
rect 66050 8206 66062 8258
rect 64542 8194 64594 8206
rect 67006 8194 67058 8206
rect 87950 8258 88002 8270
rect 87950 8194 88002 8206
rect 89406 8258 89458 8270
rect 89406 8194 89458 8206
rect 94782 8258 94834 8270
rect 96126 8258 96178 8270
rect 105758 8258 105810 8270
rect 95554 8206 95566 8258
rect 95618 8206 95630 8258
rect 104514 8206 104526 8258
rect 104578 8206 104590 8258
rect 94782 8194 94834 8206
rect 96126 8194 96178 8206
rect 105758 8194 105810 8206
rect 107102 8258 107154 8270
rect 123554 8206 123566 8258
rect 123618 8206 123630 8258
rect 125234 8206 125246 8258
rect 125298 8206 125310 8258
rect 107102 8194 107154 8206
rect 65550 8146 65602 8158
rect 63970 8094 63982 8146
rect 64034 8094 64046 8146
rect 65550 8082 65602 8094
rect 66558 8146 66610 8158
rect 89854 8146 89906 8158
rect 88274 8094 88286 8146
rect 88338 8094 88350 8146
rect 88498 8094 88510 8146
rect 88562 8094 88574 8146
rect 66558 8082 66610 8094
rect 89854 8082 89906 8094
rect 93774 8146 93826 8158
rect 95330 8094 95342 8146
rect 95394 8094 95406 8146
rect 105970 8094 105982 8146
rect 106034 8094 106046 8146
rect 106306 8094 106318 8146
rect 106370 8094 106382 8146
rect 123442 8094 123454 8146
rect 123506 8094 123518 8146
rect 93774 8082 93826 8094
rect 28030 8034 28082 8046
rect 28030 7970 28082 7982
rect 28590 8034 28642 8046
rect 28590 7970 28642 7982
rect 60734 8034 60786 8046
rect 60734 7970 60786 7982
rect 61630 8034 61682 8046
rect 61630 7970 61682 7982
rect 62078 8034 62130 8046
rect 62078 7970 62130 7982
rect 62750 8034 62802 8046
rect 62750 7970 62802 7982
rect 86606 8034 86658 8046
rect 86606 7970 86658 7982
rect 87054 8034 87106 8046
rect 87054 7970 87106 7982
rect 87614 8034 87666 8046
rect 87614 7970 87666 7982
rect 94446 8034 94498 8046
rect 94446 7970 94498 7982
rect 96686 8034 96738 8046
rect 96686 7970 96738 7982
rect 103966 8034 104018 8046
rect 103966 7970 104018 7982
rect 104750 8034 104802 8046
rect 104750 7970 104802 7982
rect 105422 8034 105474 8046
rect 105422 7970 105474 7982
rect 122446 8034 122498 8046
rect 122446 7970 122498 7982
rect 125022 8034 125074 8046
rect 125022 7970 125074 7982
rect 125918 8034 125970 8046
rect 125918 7970 125970 7982
rect 126254 8034 126306 8046
rect 126254 7970 126306 7982
rect 126814 8034 126866 8046
rect 126814 7970 126866 7982
rect 127262 8034 127314 8046
rect 127262 7970 127314 7982
rect 1344 7866 148784 7900
rect 1344 7814 38034 7866
rect 38086 7814 38138 7866
rect 38190 7814 38242 7866
rect 38294 7814 74854 7866
rect 74906 7814 74958 7866
rect 75010 7814 75062 7866
rect 75114 7814 111674 7866
rect 111726 7814 111778 7866
rect 111830 7814 111882 7866
rect 111934 7814 148494 7866
rect 148546 7814 148598 7866
rect 148650 7814 148702 7866
rect 148754 7814 148784 7866
rect 1344 7780 148784 7814
rect 67230 7698 67282 7710
rect 67230 7634 67282 7646
rect 78430 7698 78482 7710
rect 78430 7634 78482 7646
rect 85486 7698 85538 7710
rect 85486 7634 85538 7646
rect 86046 7698 86098 7710
rect 86046 7634 86098 7646
rect 89182 7698 89234 7710
rect 89182 7634 89234 7646
rect 92542 7698 92594 7710
rect 92542 7634 92594 7646
rect 93102 7698 93154 7710
rect 93102 7634 93154 7646
rect 96014 7698 96066 7710
rect 96014 7634 96066 7646
rect 107102 7698 107154 7710
rect 126814 7698 126866 7710
rect 125794 7646 125806 7698
rect 125858 7646 125870 7698
rect 107102 7634 107154 7646
rect 126814 7634 126866 7646
rect 137118 7698 137170 7710
rect 137118 7634 137170 7646
rect 139134 7698 139186 7710
rect 139134 7634 139186 7646
rect 44270 7586 44322 7598
rect 26898 7534 26910 7586
rect 26962 7534 26974 7586
rect 27234 7534 27246 7586
rect 27298 7534 27310 7586
rect 28802 7534 28814 7586
rect 28866 7534 28878 7586
rect 29362 7534 29374 7586
rect 29426 7534 29438 7586
rect 44270 7522 44322 7534
rect 59166 7586 59218 7598
rect 62862 7586 62914 7598
rect 93662 7586 93714 7598
rect 104078 7586 104130 7598
rect 61842 7534 61854 7586
rect 61906 7534 61918 7586
rect 63522 7534 63534 7586
rect 63586 7534 63598 7586
rect 65650 7534 65662 7586
rect 65714 7534 65726 7586
rect 76290 7534 76302 7586
rect 76354 7534 76366 7586
rect 76850 7534 76862 7586
rect 76914 7534 76926 7586
rect 87826 7534 87838 7586
rect 87890 7534 87902 7586
rect 88386 7534 88398 7586
rect 88450 7534 88462 7586
rect 94434 7534 94446 7586
rect 94498 7534 94510 7586
rect 94882 7534 94894 7586
rect 94946 7534 94958 7586
rect 59166 7522 59218 7534
rect 62862 7522 62914 7534
rect 93662 7522 93714 7534
rect 104078 7522 104130 7534
rect 104414 7586 104466 7598
rect 121774 7586 121826 7598
rect 105970 7534 105982 7586
rect 106034 7534 106046 7586
rect 106306 7534 106318 7586
rect 106370 7534 106382 7586
rect 116610 7534 116622 7586
rect 116674 7534 116686 7586
rect 116946 7534 116958 7586
rect 117010 7534 117022 7586
rect 104414 7522 104466 7534
rect 121774 7522 121826 7534
rect 122110 7586 122162 7598
rect 122110 7522 122162 7534
rect 26686 7474 26738 7486
rect 26686 7410 26738 7422
rect 28590 7474 28642 7486
rect 28590 7410 28642 7422
rect 30382 7474 30434 7486
rect 30382 7410 30434 7422
rect 44606 7474 44658 7486
rect 44606 7410 44658 7422
rect 59502 7474 59554 7486
rect 59502 7410 59554 7422
rect 60958 7474 61010 7486
rect 60958 7410 61010 7422
rect 61294 7474 61346 7486
rect 64206 7474 64258 7486
rect 66334 7474 66386 7486
rect 62066 7422 62078 7474
rect 62130 7422 62142 7474
rect 63410 7422 63422 7474
rect 63474 7422 63486 7474
rect 65538 7422 65550 7474
rect 65602 7422 65614 7474
rect 61294 7410 61346 7422
rect 64206 7410 64258 7422
rect 66334 7410 66386 7422
rect 77086 7474 77138 7486
rect 77086 7410 77138 7422
rect 87614 7474 87666 7486
rect 87614 7410 87666 7422
rect 95118 7474 95170 7486
rect 95118 7410 95170 7422
rect 96462 7474 96514 7486
rect 96462 7410 96514 7422
rect 105758 7474 105810 7486
rect 105758 7410 105810 7422
rect 107550 7474 107602 7486
rect 107550 7410 107602 7422
rect 116398 7474 116450 7486
rect 116398 7410 116450 7422
rect 117742 7474 117794 7486
rect 117742 7410 117794 7422
rect 122670 7474 122722 7486
rect 123330 7422 123342 7474
rect 123394 7422 123406 7474
rect 137330 7422 137342 7474
rect 137394 7422 137406 7474
rect 122670 7410 122722 7422
rect 18398 7362 18450 7374
rect 18398 7298 18450 7310
rect 19294 7362 19346 7374
rect 19294 7298 19346 7310
rect 20302 7362 20354 7374
rect 20302 7298 20354 7310
rect 29934 7362 29986 7374
rect 29934 7298 29986 7310
rect 45166 7362 45218 7374
rect 45166 7298 45218 7310
rect 47182 7362 47234 7374
rect 47182 7298 47234 7310
rect 58158 7362 58210 7374
rect 58158 7298 58210 7310
rect 58718 7362 58770 7374
rect 58718 7298 58770 7310
rect 60286 7362 60338 7374
rect 60286 7298 60338 7310
rect 75630 7362 75682 7374
rect 75630 7298 75682 7310
rect 77982 7362 78034 7374
rect 89630 7362 89682 7374
rect 86482 7310 86494 7362
rect 86546 7310 86558 7362
rect 77982 7298 78034 7310
rect 89630 7298 89682 7310
rect 103518 7362 103570 7374
rect 103518 7298 103570 7310
rect 105422 7362 105474 7374
rect 105422 7298 105474 7310
rect 115390 7362 115442 7374
rect 115390 7298 115442 7310
rect 118190 7362 118242 7374
rect 118190 7298 118242 7310
rect 121214 7362 121266 7374
rect 121214 7298 121266 7310
rect 126926 7362 126978 7374
rect 126926 7298 126978 7310
rect 127486 7362 127538 7374
rect 127486 7298 127538 7310
rect 138126 7362 138178 7374
rect 138126 7298 138178 7310
rect 138686 7362 138738 7374
rect 138686 7298 138738 7310
rect 26350 7250 26402 7262
rect 26350 7186 26402 7198
rect 28254 7250 28306 7262
rect 28254 7186 28306 7198
rect 64542 7250 64594 7262
rect 64542 7186 64594 7198
rect 66670 7250 66722 7262
rect 66670 7186 66722 7198
rect 77422 7250 77474 7262
rect 77422 7186 77474 7198
rect 87278 7250 87330 7262
rect 87278 7186 87330 7198
rect 95454 7250 95506 7262
rect 95454 7186 95506 7198
rect 116062 7250 116114 7262
rect 116062 7186 116114 7198
rect 126366 7250 126418 7262
rect 126366 7186 126418 7198
rect 127598 7250 127650 7262
rect 127598 7186 127650 7198
rect 1344 7082 148624 7116
rect 1344 7030 19624 7082
rect 19676 7030 19728 7082
rect 19780 7030 19832 7082
rect 19884 7030 56444 7082
rect 56496 7030 56548 7082
rect 56600 7030 56652 7082
rect 56704 7030 93264 7082
rect 93316 7030 93368 7082
rect 93420 7030 93472 7082
rect 93524 7030 130084 7082
rect 130136 7030 130188 7082
rect 130240 7030 130292 7082
rect 130344 7030 148624 7082
rect 1344 6996 148624 7030
rect 19630 6914 19682 6926
rect 19630 6850 19682 6862
rect 43374 6914 43426 6926
rect 43374 6850 43426 6862
rect 45950 6914 46002 6926
rect 45950 6850 46002 6862
rect 124350 6914 124402 6926
rect 124350 6850 124402 6862
rect 137454 6914 137506 6926
rect 137454 6850 137506 6862
rect 75630 6802 75682 6814
rect 28354 6750 28366 6802
rect 28418 6750 28430 6802
rect 75630 6738 75682 6750
rect 78094 6802 78146 6814
rect 78094 6738 78146 6750
rect 93998 6802 94050 6814
rect 93998 6738 94050 6750
rect 139358 6802 139410 6814
rect 139358 6738 139410 6750
rect 18286 6690 18338 6702
rect 17602 6638 17614 6690
rect 17666 6638 17678 6690
rect 18286 6626 18338 6638
rect 20526 6690 20578 6702
rect 44830 6690 44882 6702
rect 26338 6638 26350 6690
rect 26402 6638 26414 6690
rect 27122 6638 27134 6690
rect 27186 6638 27198 6690
rect 44146 6638 44158 6690
rect 44210 6638 44222 6690
rect 20526 6626 20578 6638
rect 44830 6626 44882 6638
rect 45614 6690 45666 6702
rect 45614 6626 45666 6638
rect 47966 6690 48018 6702
rect 47966 6626 48018 6638
rect 53454 6690 53506 6702
rect 61966 6690 62018 6702
rect 57138 6638 57150 6690
rect 57202 6638 57214 6690
rect 57698 6638 57710 6690
rect 57762 6638 57774 6690
rect 53454 6626 53506 6638
rect 61966 6626 62018 6638
rect 62414 6690 62466 6702
rect 66110 6690 66162 6702
rect 67678 6690 67730 6702
rect 63074 6638 63086 6690
rect 63138 6638 63150 6690
rect 66658 6638 66670 6690
rect 66722 6638 66734 6690
rect 62414 6626 62466 6638
rect 66110 6626 66162 6638
rect 67678 6626 67730 6638
rect 68126 6690 68178 6702
rect 78542 6690 78594 6702
rect 87054 6690 87106 6702
rect 90750 6690 90802 6702
rect 95454 6690 95506 6702
rect 98926 6690 98978 6702
rect 106654 6690 106706 6702
rect 69346 6638 69358 6690
rect 69410 6638 69422 6690
rect 76402 6638 76414 6690
rect 76466 6638 76478 6690
rect 77410 6638 77422 6690
rect 77474 6638 77486 6690
rect 86370 6638 86382 6690
rect 86434 6638 86446 6690
rect 87714 6638 87726 6690
rect 87778 6638 87790 6690
rect 94546 6638 94558 6690
rect 94610 6638 94622 6690
rect 95778 6638 95790 6690
rect 95842 6638 95854 6690
rect 105970 6638 105982 6690
rect 106034 6638 106046 6690
rect 68126 6626 68178 6638
rect 78542 6626 78594 6638
rect 87054 6626 87106 6638
rect 90750 6626 90802 6638
rect 95454 6626 95506 6638
rect 98926 6626 98978 6638
rect 106654 6626 106706 6638
rect 115054 6690 115106 6702
rect 115054 6626 115106 6638
rect 120654 6690 120706 6702
rect 124910 6690 124962 6702
rect 140814 6690 140866 6702
rect 121314 6638 121326 6690
rect 121378 6638 121390 6690
rect 125458 6638 125470 6690
rect 125522 6638 125534 6690
rect 136770 6638 136782 6690
rect 136834 6638 136846 6690
rect 120654 6626 120706 6638
rect 124910 6626 124962 6638
rect 140814 6626 140866 6638
rect 29598 6578 29650 6590
rect 19058 6526 19070 6578
rect 19122 6526 19134 6578
rect 19282 6526 19294 6578
rect 19346 6526 19358 6578
rect 29598 6514 29650 6526
rect 42254 6578 42306 6590
rect 42254 6514 42306 6526
rect 43038 6578 43090 6590
rect 59950 6578 60002 6590
rect 44034 6526 44046 6578
rect 44098 6526 44110 6578
rect 46162 6526 46174 6578
rect 46226 6526 46238 6578
rect 46498 6526 46510 6578
rect 46562 6526 46574 6578
rect 43038 6514 43090 6526
rect 59950 6514 60002 6526
rect 61854 6578 61906 6590
rect 61854 6514 61906 6526
rect 65326 6578 65378 6590
rect 107438 6578 107490 6590
rect 72594 6526 72606 6578
rect 72658 6526 72670 6578
rect 76290 6526 76302 6578
rect 76354 6526 76366 6578
rect 65326 6514 65378 6526
rect 107438 6514 107490 6526
rect 135662 6578 135714 6590
rect 135662 6514 135714 6526
rect 135998 6578 136050 6590
rect 137790 6578 137842 6590
rect 136658 6526 136670 6578
rect 136722 6526 136734 6578
rect 138674 6526 138686 6578
rect 138738 6526 138750 6578
rect 139122 6526 139134 6578
rect 139186 6526 139198 6578
rect 135998 6514 136050 6526
rect 137790 6514 137842 6526
rect 14590 6466 14642 6478
rect 19966 6466 20018 6478
rect 15362 6414 15374 6466
rect 15426 6414 15438 6466
rect 14590 6402 14642 6414
rect 19966 6402 20018 6414
rect 26126 6466 26178 6478
rect 26126 6402 26178 6414
rect 27358 6466 27410 6478
rect 27358 6402 27410 6414
rect 27918 6466 27970 6478
rect 27918 6402 27970 6414
rect 41918 6466 41970 6478
rect 41918 6402 41970 6414
rect 47518 6466 47570 6478
rect 47518 6402 47570 6414
rect 50542 6466 50594 6478
rect 50542 6402 50594 6414
rect 50990 6466 51042 6478
rect 52670 6466 52722 6478
rect 51314 6414 51326 6466
rect 51378 6414 51390 6466
rect 50990 6402 51042 6414
rect 52670 6402 52722 6414
rect 54014 6466 54066 6478
rect 54014 6402 54066 6414
rect 60734 6466 60786 6478
rect 60734 6402 60786 6414
rect 61294 6466 61346 6478
rect 61294 6402 61346 6414
rect 66894 6466 66946 6478
rect 66894 6402 66946 6414
rect 67566 6466 67618 6478
rect 67566 6402 67618 6414
rect 68574 6466 68626 6478
rect 68574 6402 68626 6414
rect 75294 6466 75346 6478
rect 75294 6402 75346 6414
rect 77646 6466 77698 6478
rect 77646 6402 77698 6414
rect 79102 6466 79154 6478
rect 79102 6402 79154 6414
rect 86606 6466 86658 6478
rect 94782 6466 94834 6478
rect 102510 6466 102562 6478
rect 90178 6414 90190 6466
rect 90242 6414 90254 6466
rect 98242 6414 98254 6466
rect 98306 6414 98318 6466
rect 86606 6402 86658 6414
rect 94782 6402 94834 6414
rect 102510 6402 102562 6414
rect 102958 6466 103010 6478
rect 107102 6466 107154 6478
rect 103730 6414 103742 6466
rect 103794 6414 103806 6466
rect 102958 6402 103010 6414
rect 107102 6402 107154 6414
rect 109118 6466 109170 6478
rect 109118 6402 109170 6414
rect 110798 6466 110850 6478
rect 110798 6402 110850 6414
rect 114718 6466 114770 6478
rect 114718 6402 114770 6414
rect 117294 6466 117346 6478
rect 117294 6402 117346 6414
rect 120206 6466 120258 6478
rect 128606 6466 128658 6478
rect 123778 6414 123790 6466
rect 123842 6414 123854 6466
rect 128034 6414 128046 6466
rect 128098 6414 128110 6466
rect 120206 6402 120258 6414
rect 128606 6402 128658 6414
rect 129054 6466 129106 6478
rect 129054 6402 129106 6414
rect 129390 6466 129442 6478
rect 129390 6402 129442 6414
rect 139694 6466 139746 6478
rect 139694 6402 139746 6414
rect 141262 6466 141314 6478
rect 141262 6402 141314 6414
rect 1344 6298 148784 6332
rect 1344 6246 38034 6298
rect 38086 6246 38138 6298
rect 38190 6246 38242 6298
rect 38294 6246 74854 6298
rect 74906 6246 74958 6298
rect 75010 6246 75062 6298
rect 75114 6246 111674 6298
rect 111726 6246 111778 6298
rect 111830 6246 111882 6298
rect 111934 6246 148494 6298
rect 148546 6246 148598 6298
rect 148650 6246 148702 6298
rect 148754 6246 148784 6298
rect 1344 6212 148784 6246
rect 16158 6130 16210 6142
rect 16158 6066 16210 6078
rect 31390 6130 31442 6142
rect 31390 6066 31442 6078
rect 38894 6130 38946 6142
rect 38894 6066 38946 6078
rect 39454 6130 39506 6142
rect 53566 6130 53618 6142
rect 39778 6078 39790 6130
rect 39842 6078 39854 6130
rect 46722 6078 46734 6130
rect 46786 6078 46798 6130
rect 39454 6066 39506 6078
rect 53566 6066 53618 6078
rect 55134 6130 55186 6142
rect 63982 6130 64034 6142
rect 62738 6078 62750 6130
rect 62802 6078 62814 6130
rect 55134 6066 55186 6078
rect 63982 6066 64034 6078
rect 65326 6130 65378 6142
rect 87838 6130 87890 6142
rect 66098 6078 66110 6130
rect 66162 6078 66174 6130
rect 65326 6066 65378 6078
rect 87838 6066 87890 6078
rect 95342 6130 95394 6142
rect 95342 6066 95394 6078
rect 95790 6130 95842 6142
rect 95790 6066 95842 6078
rect 98254 6130 98306 6142
rect 98254 6066 98306 6078
rect 104414 6130 104466 6142
rect 109230 6130 109282 6142
rect 108210 6078 108222 6130
rect 108274 6078 108286 6130
rect 104414 6066 104466 6078
rect 109230 6066 109282 6078
rect 117854 6130 117906 6142
rect 117854 6066 117906 6078
rect 118302 6130 118354 6142
rect 126142 6130 126194 6142
rect 125570 6078 125582 6130
rect 125634 6078 125646 6130
rect 118302 6066 118354 6078
rect 126142 6066 126194 6078
rect 126590 6130 126642 6142
rect 126590 6066 126642 6078
rect 127262 6130 127314 6142
rect 127262 6066 127314 6078
rect 129390 6130 129442 6142
rect 129390 6066 129442 6078
rect 134206 6130 134258 6142
rect 134206 6066 134258 6078
rect 135774 6130 135826 6142
rect 135774 6066 135826 6078
rect 138574 6130 138626 6142
rect 138574 6066 138626 6078
rect 19630 6018 19682 6030
rect 18722 5966 18734 6018
rect 18786 5966 18798 6018
rect 19630 5954 19682 5966
rect 19966 6018 20018 6030
rect 19966 5954 20018 5966
rect 30606 6018 30658 6030
rect 30606 5954 30658 5966
rect 31726 6018 31778 6030
rect 31726 5954 31778 5966
rect 53118 6018 53170 6030
rect 53118 5954 53170 5966
rect 64318 6018 64370 6030
rect 64318 5954 64370 5966
rect 75294 6018 75346 6030
rect 75294 5954 75346 5966
rect 76526 6018 76578 6030
rect 76526 5954 76578 5966
rect 79886 6018 79938 6030
rect 79886 5954 79938 5966
rect 87502 6018 87554 6030
rect 87502 5954 87554 5966
rect 109342 6018 109394 6030
rect 109342 5954 109394 5966
rect 110238 6018 110290 6030
rect 110238 5954 110290 5966
rect 115950 6018 116002 6030
rect 140142 6018 140194 6030
rect 132962 5966 132974 6018
rect 133026 5966 133038 6018
rect 137442 5966 137454 6018
rect 137506 5966 137518 6018
rect 138002 5966 138014 6018
rect 138066 5966 138078 6018
rect 115950 5954 116002 5966
rect 140142 5954 140194 5966
rect 140702 6018 140754 6030
rect 140702 5954 140754 5966
rect 141262 6018 141314 6030
rect 141262 5954 141314 5966
rect 17838 5906 17890 5918
rect 15922 5854 15934 5906
rect 15986 5854 15998 5906
rect 17838 5842 17890 5854
rect 18174 5906 18226 5918
rect 21534 5906 21586 5918
rect 18946 5854 18958 5906
rect 19010 5854 19022 5906
rect 18174 5842 18226 5854
rect 21534 5842 21586 5854
rect 27694 5906 27746 5918
rect 43822 5906 43874 5918
rect 47630 5906 47682 5918
rect 28242 5854 28254 5906
rect 28306 5854 28318 5906
rect 44258 5854 44270 5906
rect 44322 5854 44334 5906
rect 27694 5842 27746 5854
rect 43822 5842 43874 5854
rect 47630 5842 47682 5854
rect 57822 5906 57874 5918
rect 57822 5842 57874 5854
rect 59838 5906 59890 5918
rect 69022 5906 69074 5918
rect 79438 5906 79490 5918
rect 105310 5906 105362 5918
rect 111022 5906 111074 5918
rect 60498 5854 60510 5906
rect 60562 5854 60574 5906
rect 68338 5854 68350 5906
rect 68402 5854 68414 5906
rect 75058 5854 75070 5906
rect 75122 5854 75134 5906
rect 78754 5854 78766 5906
rect 78818 5854 78830 5906
rect 95106 5854 95118 5906
rect 95170 5854 95182 5906
rect 105746 5854 105758 5906
rect 105810 5854 105822 5906
rect 59838 5842 59890 5854
rect 69022 5842 69074 5854
rect 79438 5842 79490 5854
rect 105310 5842 105362 5854
rect 111022 5842 111074 5854
rect 112366 5906 112418 5918
rect 112366 5842 112418 5854
rect 113262 5906 113314 5918
rect 117518 5906 117570 5918
rect 113698 5854 113710 5906
rect 113762 5854 113774 5906
rect 113262 5842 113314 5854
rect 117518 5842 117570 5854
rect 121998 5906 122050 5918
rect 121998 5842 122050 5854
rect 122446 5906 122498 5918
rect 132414 5906 132466 5918
rect 139582 5906 139634 5918
rect 123106 5854 123118 5906
rect 123170 5854 123182 5906
rect 129154 5854 129166 5906
rect 129218 5854 129230 5906
rect 133186 5854 133198 5906
rect 133250 5854 133262 5906
rect 122446 5842 122498 5854
rect 132414 5842 132466 5854
rect 139582 5842 139634 5854
rect 9774 5794 9826 5806
rect 9774 5730 9826 5742
rect 10110 5794 10162 5806
rect 10110 5730 10162 5742
rect 11678 5794 11730 5806
rect 11678 5730 11730 5742
rect 16942 5794 16994 5806
rect 16942 5730 16994 5742
rect 20638 5794 20690 5806
rect 20638 5730 20690 5742
rect 21198 5794 21250 5806
rect 21198 5730 21250 5742
rect 55694 5794 55746 5806
rect 55694 5730 55746 5742
rect 56366 5794 56418 5806
rect 56366 5730 56418 5742
rect 56814 5794 56866 5806
rect 56814 5730 56866 5742
rect 57486 5794 57538 5806
rect 57486 5730 57538 5742
rect 58270 5794 58322 5806
rect 58270 5730 58322 5742
rect 58830 5794 58882 5806
rect 58830 5730 58882 5742
rect 59390 5794 59442 5806
rect 59390 5730 59442 5742
rect 69358 5794 69410 5806
rect 69358 5730 69410 5742
rect 79998 5794 80050 5806
rect 79998 5730 80050 5742
rect 80446 5794 80498 5806
rect 80446 5730 80498 5742
rect 81342 5794 81394 5806
rect 81342 5730 81394 5742
rect 86830 5794 86882 5806
rect 86830 5730 86882 5742
rect 89406 5794 89458 5806
rect 89406 5730 89458 5742
rect 89966 5794 90018 5806
rect 89966 5730 90018 5742
rect 96574 5794 96626 5806
rect 96574 5730 96626 5742
rect 97246 5794 97298 5806
rect 97246 5730 97298 5742
rect 98366 5794 98418 5806
rect 98366 5730 98418 5742
rect 98926 5794 98978 5806
rect 98926 5730 98978 5742
rect 102734 5794 102786 5806
rect 102734 5730 102786 5742
rect 103182 5794 103234 5806
rect 103182 5730 103234 5742
rect 103630 5794 103682 5806
rect 103630 5730 103682 5742
rect 104302 5794 104354 5806
rect 104302 5730 104354 5742
rect 109902 5794 109954 5806
rect 109902 5730 109954 5742
rect 111582 5794 111634 5806
rect 111582 5730 111634 5742
rect 121550 5794 121602 5806
rect 121550 5730 121602 5742
rect 126702 5794 126754 5806
rect 126702 5730 126754 5742
rect 127374 5794 127426 5806
rect 127374 5730 127426 5742
rect 128046 5794 128098 5806
rect 128046 5730 128098 5742
rect 129838 5794 129890 5806
rect 129838 5730 129890 5742
rect 130286 5794 130338 5806
rect 130286 5730 130338 5742
rect 133758 5794 133810 5806
rect 133758 5730 133810 5742
rect 134654 5794 134706 5806
rect 134654 5730 134706 5742
rect 136222 5794 136274 5806
rect 136222 5730 136274 5742
rect 20526 5682 20578 5694
rect 20526 5618 20578 5630
rect 47294 5682 47346 5694
rect 59278 5682 59330 5694
rect 56354 5630 56366 5682
rect 56418 5679 56430 5682
rect 56914 5679 56926 5682
rect 56418 5633 56926 5679
rect 56418 5630 56430 5633
rect 56914 5630 56926 5633
rect 56978 5630 56990 5682
rect 47294 5618 47346 5630
rect 59278 5618 59330 5630
rect 63534 5682 63586 5694
rect 63534 5618 63586 5630
rect 75742 5682 75794 5694
rect 75742 5618 75794 5630
rect 89294 5682 89346 5694
rect 89294 5618 89346 5630
rect 97358 5682 97410 5694
rect 97358 5618 97410 5630
rect 103742 5682 103794 5694
rect 103742 5618 103794 5630
rect 108782 5682 108834 5694
rect 108782 5618 108834 5630
rect 116734 5682 116786 5694
rect 116734 5618 116786 5630
rect 127934 5682 127986 5694
rect 127934 5618 127986 5630
rect 132078 5682 132130 5694
rect 132078 5618 132130 5630
rect 138238 5682 138290 5694
rect 138238 5618 138290 5630
rect 1344 5514 148624 5548
rect 1344 5462 19624 5514
rect 19676 5462 19728 5514
rect 19780 5462 19832 5514
rect 19884 5462 56444 5514
rect 56496 5462 56548 5514
rect 56600 5462 56652 5514
rect 56704 5462 93264 5514
rect 93316 5462 93368 5514
rect 93420 5462 93472 5514
rect 93524 5462 130084 5514
rect 130136 5462 130188 5514
rect 130240 5462 130292 5514
rect 130344 5462 148624 5514
rect 1344 5428 148624 5462
rect 20750 5346 20802 5358
rect 20750 5282 20802 5294
rect 29710 5346 29762 5358
rect 29710 5282 29762 5294
rect 47070 5346 47122 5358
rect 47070 5282 47122 5294
rect 58830 5346 58882 5358
rect 58830 5282 58882 5294
rect 67678 5346 67730 5358
rect 67678 5282 67730 5294
rect 80894 5346 80946 5358
rect 80894 5282 80946 5294
rect 90302 5346 90354 5358
rect 90302 5282 90354 5294
rect 98030 5346 98082 5358
rect 98030 5282 98082 5294
rect 103070 5346 103122 5358
rect 103070 5282 103122 5294
rect 109566 5346 109618 5358
rect 109566 5282 109618 5294
rect 115614 5346 115666 5358
rect 115614 5282 115666 5294
rect 118526 5346 118578 5358
rect 118526 5282 118578 5294
rect 130846 5346 130898 5358
rect 130846 5282 130898 5294
rect 133422 5346 133474 5358
rect 133422 5282 133474 5294
rect 137118 5346 137170 5358
rect 137118 5282 137170 5294
rect 16718 5234 16770 5246
rect 16718 5170 16770 5182
rect 28590 5234 28642 5246
rect 28590 5170 28642 5182
rect 46398 5234 46450 5246
rect 46398 5170 46450 5182
rect 47182 5234 47234 5246
rect 47182 5170 47234 5182
rect 47630 5234 47682 5246
rect 47630 5170 47682 5182
rect 52670 5234 52722 5246
rect 52670 5170 52722 5182
rect 53678 5234 53730 5246
rect 67790 5234 67842 5246
rect 63970 5182 63982 5234
rect 64034 5182 64046 5234
rect 53678 5170 53730 5182
rect 67790 5170 67842 5182
rect 68238 5234 68290 5246
rect 68238 5170 68290 5182
rect 69694 5234 69746 5246
rect 108222 5234 108274 5246
rect 75506 5182 75518 5234
rect 75570 5182 75582 5234
rect 69694 5170 69746 5182
rect 108222 5170 108274 5182
rect 109230 5234 109282 5246
rect 109230 5170 109282 5182
rect 110910 5234 110962 5246
rect 110910 5170 110962 5182
rect 111358 5234 111410 5246
rect 111358 5170 111410 5182
rect 114942 5234 114994 5246
rect 114942 5170 114994 5182
rect 115502 5234 115554 5246
rect 115502 5170 115554 5182
rect 116286 5234 116338 5246
rect 116286 5170 116338 5182
rect 116958 5234 117010 5246
rect 116958 5170 117010 5182
rect 119534 5234 119586 5246
rect 119534 5170 119586 5182
rect 124350 5234 124402 5246
rect 124350 5170 124402 5182
rect 131854 5234 131906 5246
rect 131854 5170 131906 5182
rect 132190 5234 132242 5246
rect 132190 5170 132242 5182
rect 134766 5234 134818 5246
rect 134766 5170 134818 5182
rect 135214 5234 135266 5246
rect 135214 5170 135266 5182
rect 138462 5234 138514 5246
rect 138462 5170 138514 5182
rect 139022 5234 139074 5246
rect 139022 5170 139074 5182
rect 139470 5234 139522 5246
rect 139470 5170 139522 5182
rect 139806 5234 139858 5246
rect 139806 5170 139858 5182
rect 140814 5234 140866 5246
rect 140814 5170 140866 5182
rect 16158 5122 16210 5134
rect 7746 5070 7758 5122
rect 7810 5070 7822 5122
rect 8194 5070 8206 5122
rect 8258 5070 8270 5122
rect 10434 5070 10446 5122
rect 10498 5070 10510 5122
rect 16158 5058 16210 5070
rect 17278 5122 17330 5134
rect 21534 5122 21586 5134
rect 17714 5070 17726 5122
rect 17778 5070 17790 5122
rect 17278 5058 17330 5070
rect 21534 5058 21586 5070
rect 25118 5122 25170 5134
rect 41022 5122 41074 5134
rect 44718 5122 44770 5134
rect 25554 5070 25566 5122
rect 25618 5070 25630 5122
rect 41682 5070 41694 5122
rect 41746 5070 41758 5122
rect 25118 5058 25170 5070
rect 41022 5058 41074 5070
rect 44718 5058 44770 5070
rect 45390 5122 45442 5134
rect 45390 5058 45442 5070
rect 46510 5122 46562 5134
rect 46510 5058 46562 5070
rect 52334 5122 52386 5134
rect 52334 5058 52386 5070
rect 55358 5122 55410 5134
rect 67118 5122 67170 5134
rect 77422 5122 77474 5134
rect 86382 5122 86434 5134
rect 89854 5122 89906 5134
rect 55682 5070 55694 5122
rect 55746 5070 55758 5122
rect 62850 5070 62862 5122
rect 62914 5070 62926 5122
rect 72594 5070 72606 5122
rect 72658 5070 72670 5122
rect 77746 5070 77758 5122
rect 77810 5070 77822 5122
rect 86706 5070 86718 5122
rect 86770 5070 86782 5122
rect 55358 5058 55410 5070
rect 67118 5058 67170 5070
rect 77422 5058 77474 5070
rect 86382 5058 86434 5070
rect 89854 5058 89906 5070
rect 90414 5122 90466 5134
rect 90414 5058 90466 5070
rect 93886 5122 93938 5134
rect 93886 5058 93938 5070
rect 94558 5122 94610 5134
rect 102622 5122 102674 5134
rect 106766 5122 106818 5134
rect 116174 5122 116226 5134
rect 94882 5070 94894 5122
rect 94946 5070 94958 5122
rect 106082 5070 106094 5122
rect 106146 5070 106158 5122
rect 110226 5070 110238 5122
rect 110290 5070 110302 5122
rect 94558 5058 94610 5070
rect 102622 5058 102674 5070
rect 106766 5058 106818 5070
rect 116174 5058 116226 5070
rect 120206 5122 120258 5134
rect 120206 5058 120258 5070
rect 120878 5122 120930 5134
rect 124910 5122 124962 5134
rect 128382 5122 128434 5134
rect 130958 5122 131010 5134
rect 121202 5070 121214 5122
rect 121266 5070 121278 5122
rect 128034 5070 128046 5122
rect 128098 5070 128110 5122
rect 129266 5070 129278 5122
rect 129330 5070 129342 5122
rect 120878 5058 120930 5070
rect 124910 5058 124962 5070
rect 128382 5058 128434 5070
rect 130958 5058 131010 5070
rect 133086 5122 133138 5134
rect 134194 5070 134206 5122
rect 134258 5070 134270 5122
rect 137778 5070 137790 5122
rect 137842 5070 137854 5122
rect 133086 5058 133138 5070
rect 12126 5010 12178 5022
rect 12126 4946 12178 4958
rect 29598 5010 29650 5022
rect 29598 4946 29650 4958
rect 54350 5010 54402 5022
rect 54350 4946 54402 4958
rect 54686 5010 54738 5022
rect 54686 4946 54738 4958
rect 59278 5010 59330 5022
rect 59278 4946 59330 4958
rect 60286 5010 60338 5022
rect 60286 4946 60338 4958
rect 60622 5010 60674 5022
rect 60622 4946 60674 4958
rect 85262 5010 85314 5022
rect 85262 4946 85314 4958
rect 85598 5010 85650 5022
rect 85598 4946 85650 4958
rect 107550 5010 107602 5022
rect 129054 5010 129106 5022
rect 110114 4958 110126 5010
rect 110178 4958 110190 5010
rect 117730 4958 117742 5010
rect 117794 4958 117806 5010
rect 118290 4958 118302 5010
rect 118354 4958 118366 5010
rect 107550 4946 107602 4958
rect 129054 4946 129106 4958
rect 130286 5010 130338 5022
rect 135774 5010 135826 5022
rect 133970 4958 133982 5010
rect 134034 4958 134046 5010
rect 130286 4946 130338 4958
rect 135774 4946 135826 4958
rect 136110 5010 136162 5022
rect 136110 4946 136162 4958
rect 136782 5010 136834 5022
rect 137890 4958 137902 5010
rect 137954 4958 137966 5010
rect 136782 4946 136834 4958
rect 6190 4898 6242 4910
rect 6190 4834 6242 4846
rect 11342 4898 11394 4910
rect 11342 4834 11394 4846
rect 12238 4898 12290 4910
rect 12238 4834 12290 4846
rect 12686 4898 12738 4910
rect 22094 4898 22146 4910
rect 30158 4898 30210 4910
rect 59614 4898 59666 4910
rect 20066 4846 20078 4898
rect 20130 4846 20142 4898
rect 28018 4846 28030 4898
rect 28082 4846 28094 4898
rect 44146 4846 44158 4898
rect 44210 4846 44222 4898
rect 58258 4846 58270 4898
rect 58322 4846 58334 4898
rect 12686 4834 12738 4846
rect 22094 4834 22146 4846
rect 30158 4834 30210 4846
rect 59614 4834 59666 4846
rect 69358 4898 69410 4910
rect 84478 4898 84530 4910
rect 90862 4898 90914 4910
rect 107214 4898 107266 4910
rect 80098 4846 80110 4898
rect 80162 4846 80174 4898
rect 89282 4846 89294 4898
rect 89346 4846 89358 4898
rect 97346 4846 97358 4898
rect 97410 4846 97422 4898
rect 103730 4846 103742 4898
rect 103794 4846 103806 4898
rect 69358 4834 69410 4846
rect 84478 4834 84530 4846
rect 90862 4834 90914 4846
rect 107214 4834 107266 4846
rect 108110 4898 108162 4910
rect 108110 4834 108162 4846
rect 118862 4898 118914 4910
rect 129950 4898 130002 4910
rect 123778 4846 123790 4898
rect 123842 4846 123854 4898
rect 125682 4846 125694 4898
rect 125746 4846 125758 4898
rect 118862 4834 118914 4846
rect 129950 4834 130002 4846
rect 1344 4730 148784 4764
rect 1344 4678 38034 4730
rect 38086 4678 38138 4730
rect 38190 4678 38242 4730
rect 38294 4678 74854 4730
rect 74906 4678 74958 4730
rect 75010 4678 75062 4730
rect 75114 4678 111674 4730
rect 111726 4678 111778 4730
rect 111830 4678 111882 4730
rect 111934 4678 148494 4730
rect 148546 4678 148598 4730
rect 148650 4678 148702 4730
rect 148754 4678 148784 4730
rect 1344 4644 148784 4678
rect 8206 4562 8258 4574
rect 13358 4562 13410 4574
rect 12562 4510 12574 4562
rect 12626 4510 12638 4562
rect 8206 4498 8258 4510
rect 13358 4498 13410 4510
rect 13694 4562 13746 4574
rect 13694 4498 13746 4510
rect 15710 4562 15762 4574
rect 15710 4498 15762 4510
rect 16270 4562 16322 4574
rect 21758 4562 21810 4574
rect 18162 4510 18174 4562
rect 18226 4510 18238 4562
rect 16270 4498 16322 4510
rect 21758 4498 21810 4510
rect 26462 4562 26514 4574
rect 26462 4498 26514 4510
rect 28030 4562 28082 4574
rect 28030 4498 28082 4510
rect 28702 4562 28754 4574
rect 28702 4498 28754 4510
rect 29150 4562 29202 4574
rect 29150 4498 29202 4510
rect 46734 4562 46786 4574
rect 46734 4498 46786 4510
rect 48190 4562 48242 4574
rect 48190 4498 48242 4510
rect 54126 4562 54178 4574
rect 54126 4498 54178 4510
rect 57934 4562 57986 4574
rect 57934 4498 57986 4510
rect 58830 4562 58882 4574
rect 58830 4498 58882 4510
rect 65326 4562 65378 4574
rect 69806 4562 69858 4574
rect 66098 4510 66110 4562
rect 66162 4510 66174 4562
rect 65326 4498 65378 4510
rect 69806 4498 69858 4510
rect 70254 4562 70306 4574
rect 70254 4498 70306 4510
rect 79998 4562 80050 4574
rect 79998 4498 80050 4510
rect 85934 4562 85986 4574
rect 85934 4498 85986 4510
rect 86382 4562 86434 4574
rect 86382 4498 86434 4510
rect 88510 4562 88562 4574
rect 88510 4498 88562 4510
rect 89630 4562 89682 4574
rect 89630 4498 89682 4510
rect 90078 4562 90130 4574
rect 90078 4498 90130 4510
rect 103966 4562 104018 4574
rect 103966 4498 104018 4510
rect 104414 4562 104466 4574
rect 110910 4562 110962 4574
rect 108098 4510 108110 4562
rect 108162 4510 108174 4562
rect 104414 4498 104466 4510
rect 110910 4498 110962 4510
rect 114830 4562 114882 4574
rect 118974 4562 119026 4574
rect 115602 4510 115614 4562
rect 115666 4510 115678 4562
rect 114830 4498 114882 4510
rect 118974 4498 119026 4510
rect 121326 4562 121378 4574
rect 128046 4562 128098 4574
rect 133646 4562 133698 4574
rect 125794 4510 125806 4562
rect 125858 4510 125870 4562
rect 131954 4510 131966 4562
rect 132018 4510 132030 4562
rect 121326 4498 121378 4510
rect 128046 4498 128098 4510
rect 133646 4498 133698 4510
rect 137118 4562 137170 4574
rect 137118 4498 137170 4510
rect 138350 4562 138402 4574
rect 138350 4498 138402 4510
rect 138798 4562 138850 4574
rect 138798 4498 138850 4510
rect 142046 4562 142098 4574
rect 142046 4498 142098 4510
rect 145742 4562 145794 4574
rect 145742 4498 145794 4510
rect 7758 4450 7810 4462
rect 7758 4386 7810 4398
rect 16830 4450 16882 4462
rect 16830 4386 16882 4398
rect 27134 4450 27186 4462
rect 27134 4386 27186 4398
rect 27470 4450 27522 4462
rect 27470 4386 27522 4398
rect 28142 4450 28194 4462
rect 28142 4386 28194 4398
rect 29598 4450 29650 4462
rect 56366 4450 56418 4462
rect 54674 4398 54686 4450
rect 54738 4398 54750 4450
rect 55234 4398 55246 4450
rect 55298 4398 55310 4450
rect 29598 4386 29650 4398
rect 56366 4386 56418 4398
rect 58494 4450 58546 4462
rect 79886 4450 79938 4462
rect 61282 4398 61294 4450
rect 61346 4398 61358 4450
rect 78418 4398 78430 4450
rect 78482 4398 78494 4450
rect 58494 4386 58546 4398
rect 79886 4386 79938 4398
rect 80446 4450 80498 4462
rect 80446 4386 80498 4398
rect 89294 4450 89346 4462
rect 89294 4386 89346 4398
rect 111358 4450 111410 4462
rect 111358 4386 111410 4398
rect 119310 4450 119362 4462
rect 119310 4386 119362 4398
rect 127486 4450 127538 4462
rect 127486 4386 127538 4398
rect 128158 4450 128210 4462
rect 128158 4386 128210 4398
rect 137454 4450 137506 4462
rect 137454 4386 137506 4398
rect 6974 4338 7026 4350
rect 8318 4338 8370 4350
rect 5842 4286 5854 4338
rect 5906 4286 5918 4338
rect 7522 4286 7534 4338
rect 7586 4286 7598 4338
rect 6974 4274 7026 4286
rect 8318 4274 8370 4286
rect 8542 4338 8594 4350
rect 8542 4274 8594 4286
rect 8766 4338 8818 4350
rect 8766 4274 8818 4286
rect 8990 4338 9042 4350
rect 8990 4274 9042 4286
rect 9886 4338 9938 4350
rect 15374 4338 15426 4350
rect 10210 4286 10222 4338
rect 10274 4286 10286 4338
rect 9886 4274 9938 4286
rect 15374 4274 15426 4286
rect 17614 4338 17666 4350
rect 21310 4338 21362 4350
rect 20626 4286 20638 4338
rect 20690 4286 20702 4338
rect 17614 4274 17666 4286
rect 21310 4274 21362 4286
rect 22094 4338 22146 4350
rect 22094 4274 22146 4286
rect 22542 4338 22594 4350
rect 22542 4274 22594 4286
rect 26126 4338 26178 4350
rect 53454 4338 53506 4350
rect 52882 4286 52894 4338
rect 52946 4286 52958 4338
rect 26126 4274 26178 4286
rect 53454 4274 53506 4286
rect 54462 4338 54514 4350
rect 54462 4274 54514 4286
rect 56702 4338 56754 4350
rect 56702 4274 56754 4286
rect 57598 4338 57650 4350
rect 69470 4338 69522 4350
rect 63858 4286 63870 4338
rect 63922 4286 63934 4338
rect 68338 4286 68350 4338
rect 68402 4286 68414 4338
rect 68898 4286 68910 4338
rect 68962 4286 68974 4338
rect 57598 4274 57650 4286
rect 69470 4274 69522 4286
rect 70702 4338 70754 4350
rect 70702 4274 70754 4286
rect 72606 4338 72658 4350
rect 79102 4338 79154 4350
rect 74834 4286 74846 4338
rect 74898 4286 74910 4338
rect 72606 4274 72658 4286
rect 79102 4274 79154 4286
rect 105310 4338 105362 4350
rect 114382 4338 114434 4350
rect 118526 4338 118578 4350
rect 105746 4286 105758 4338
rect 105810 4286 105822 4338
rect 110450 4286 110462 4338
rect 110514 4286 110526 4338
rect 117954 4286 117966 4338
rect 118018 4286 118030 4338
rect 105310 4274 105362 4286
rect 114382 4274 114434 4286
rect 118526 4274 118578 4286
rect 122222 4338 122274 4350
rect 122222 4274 122274 4286
rect 122894 4338 122946 4350
rect 128942 4338 128994 4350
rect 138014 4338 138066 4350
rect 123330 4286 123342 4338
rect 123394 4286 123406 4338
rect 127250 4286 127262 4338
rect 127314 4286 127326 4338
rect 129490 4286 129502 4338
rect 129554 4286 129566 4338
rect 133858 4286 133870 4338
rect 133922 4286 133934 4338
rect 122894 4274 122946 4286
rect 128942 4274 128994 4286
rect 138014 4274 138066 4286
rect 141710 4338 141762 4350
rect 145954 4286 145966 4338
rect 146018 4286 146030 4338
rect 141710 4274 141762 4286
rect 6526 4226 6578 4238
rect 4834 4174 4846 4226
rect 4898 4174 4910 4226
rect 6526 4162 6578 4174
rect 14478 4226 14530 4238
rect 14478 4162 14530 4174
rect 14926 4226 14978 4238
rect 14926 4162 14978 4174
rect 16942 4226 16994 4238
rect 16942 4162 16994 4174
rect 25006 4226 25058 4238
rect 25006 4162 25058 4174
rect 25678 4226 25730 4238
rect 25678 4162 25730 4174
rect 31726 4226 31778 4238
rect 31726 4162 31778 4174
rect 32958 4226 33010 4238
rect 32958 4162 33010 4174
rect 33966 4226 34018 4238
rect 33966 4162 34018 4174
rect 36878 4226 36930 4238
rect 36878 4162 36930 4174
rect 37214 4226 37266 4238
rect 37214 4162 37266 4174
rect 38670 4226 38722 4238
rect 38670 4162 38722 4174
rect 40798 4226 40850 4238
rect 40798 4162 40850 4174
rect 42590 4226 42642 4238
rect 42590 4162 42642 4174
rect 44718 4226 44770 4238
rect 44718 4162 44770 4174
rect 45054 4226 45106 4238
rect 45054 4162 45106 4174
rect 47182 4226 47234 4238
rect 47182 4162 47234 4174
rect 48750 4226 48802 4238
rect 55918 4226 55970 4238
rect 51874 4174 51886 4226
rect 51938 4174 51950 4226
rect 48750 4162 48802 4174
rect 55918 4162 55970 4174
rect 81790 4226 81842 4238
rect 81790 4162 81842 4174
rect 93550 4226 93602 4238
rect 93550 4162 93602 4174
rect 97582 4226 97634 4238
rect 97582 4162 97634 4174
rect 101614 4226 101666 4238
rect 113710 4226 113762 4238
rect 109442 4174 109454 4226
rect 109506 4174 109518 4226
rect 101614 4162 101666 4174
rect 113710 4162 113762 4174
rect 121774 4226 121826 4238
rect 121774 4162 121826 4174
rect 126366 4226 126418 4238
rect 126366 4162 126418 4174
rect 132974 4226 133026 4238
rect 132974 4162 133026 4174
rect 134430 4226 134482 4238
rect 134430 4162 134482 4174
rect 141262 4226 141314 4238
rect 141262 4162 141314 4174
rect 145294 4226 145346 4238
rect 145294 4162 145346 4174
rect 108782 4114 108834 4126
rect 108782 4050 108834 4062
rect 132638 4114 132690 4126
rect 132638 4050 132690 4062
rect 1344 3946 148624 3980
rect 1344 3894 19624 3946
rect 19676 3894 19728 3946
rect 19780 3894 19832 3946
rect 19884 3894 56444 3946
rect 56496 3894 56548 3946
rect 56600 3894 56652 3946
rect 56704 3894 93264 3946
rect 93316 3894 93368 3946
rect 93420 3894 93472 3946
rect 93524 3894 130084 3946
rect 130136 3894 130188 3946
rect 130240 3894 130292 3946
rect 130344 3894 148624 3946
rect 1344 3860 148624 3894
rect 12238 3778 12290 3790
rect 8082 3726 8094 3778
rect 8146 3726 8158 3778
rect 12238 3714 12290 3726
rect 17614 3778 17666 3790
rect 17614 3714 17666 3726
rect 17950 3778 18002 3790
rect 17950 3714 18002 3726
rect 18734 3778 18786 3790
rect 18734 3714 18786 3726
rect 54798 3778 54850 3790
rect 54798 3714 54850 3726
rect 55134 3778 55186 3790
rect 55134 3714 55186 3726
rect 108110 3778 108162 3790
rect 108110 3714 108162 3726
rect 108446 3778 108498 3790
rect 108446 3714 108498 3726
rect 127262 3778 127314 3790
rect 127262 3714 127314 3726
rect 12350 3666 12402 3678
rect 12350 3602 12402 3614
rect 12910 3666 12962 3678
rect 21534 3666 21586 3678
rect 75630 3666 75682 3678
rect 19618 3614 19630 3666
rect 19682 3614 19694 3666
rect 35298 3614 35310 3666
rect 35362 3614 35374 3666
rect 43362 3614 43374 3666
rect 43426 3614 43438 3666
rect 47394 3614 47406 3666
rect 47458 3614 47470 3666
rect 12910 3602 12962 3614
rect 21534 3602 21586 3614
rect 75630 3602 75682 3614
rect 78990 3666 79042 3678
rect 78990 3602 79042 3614
rect 94670 3666 94722 3678
rect 94670 3602 94722 3614
rect 102734 3666 102786 3678
rect 102734 3602 102786 3614
rect 110686 3666 110738 3678
rect 115726 3666 115778 3678
rect 112354 3614 112366 3666
rect 112418 3614 112430 3666
rect 110686 3602 110738 3614
rect 115726 3602 115778 3614
rect 119310 3666 119362 3678
rect 119310 3602 119362 3614
rect 123342 3666 123394 3678
rect 123342 3602 123394 3614
rect 123790 3666 123842 3678
rect 123790 3602 123842 3614
rect 127374 3666 127426 3678
rect 127374 3602 127426 3614
rect 131630 3666 131682 3678
rect 131630 3602 131682 3614
rect 135886 3666 135938 3678
rect 135886 3602 135938 3614
rect 138014 3666 138066 3678
rect 138014 3602 138066 3614
rect 139918 3666 139970 3678
rect 139918 3602 139970 3614
rect 143950 3666 144002 3678
rect 143950 3602 144002 3614
rect 5854 3554 5906 3566
rect 8542 3554 8594 3566
rect 7298 3502 7310 3554
rect 7362 3502 7374 3554
rect 5854 3490 5906 3502
rect 8542 3490 8594 3502
rect 8654 3554 8706 3566
rect 8654 3490 8706 3502
rect 8766 3554 8818 3566
rect 51998 3554 52050 3566
rect 15250 3502 15262 3554
rect 15314 3502 15326 3554
rect 16482 3502 16494 3554
rect 16546 3502 16558 3554
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 20626 3502 20638 3554
rect 20690 3502 20702 3554
rect 22306 3502 22318 3554
rect 22370 3502 22382 3554
rect 26562 3502 26574 3554
rect 26626 3502 26638 3554
rect 31378 3502 31390 3554
rect 31442 3502 31454 3554
rect 36306 3502 36318 3554
rect 36370 3502 36382 3554
rect 40226 3502 40238 3554
rect 40290 3502 40302 3554
rect 41234 3502 41246 3554
rect 41298 3502 41310 3554
rect 42242 3502 42254 3554
rect 42306 3502 42318 3554
rect 44146 3502 44158 3554
rect 44210 3502 44222 3554
rect 46162 3502 46174 3554
rect 46226 3502 46238 3554
rect 48066 3502 48078 3554
rect 48130 3502 48142 3554
rect 8766 3490 8818 3502
rect 51998 3490 52050 3502
rect 55918 3554 55970 3566
rect 58942 3554 58994 3566
rect 57922 3502 57934 3554
rect 57986 3502 57998 3554
rect 55918 3490 55970 3502
rect 58942 3490 58994 3502
rect 59838 3554 59890 3566
rect 62414 3554 62466 3566
rect 61618 3502 61630 3554
rect 61682 3502 61694 3554
rect 59838 3490 59890 3502
rect 62414 3490 62466 3502
rect 63646 3554 63698 3566
rect 67566 3554 67618 3566
rect 70254 3554 70306 3566
rect 65538 3502 65550 3554
rect 65602 3502 65614 3554
rect 66546 3502 66558 3554
rect 66610 3502 66622 3554
rect 69682 3502 69694 3554
rect 69746 3502 69758 3554
rect 63646 3490 63698 3502
rect 67566 3490 67618 3502
rect 70254 3490 70306 3502
rect 70590 3554 70642 3566
rect 70590 3490 70642 3502
rect 71710 3554 71762 3566
rect 82910 3554 82962 3566
rect 98702 3554 98754 3566
rect 118302 3554 118354 3566
rect 131070 3554 131122 3566
rect 73602 3502 73614 3554
rect 73666 3502 73678 3554
rect 77522 3502 77534 3554
rect 77586 3502 77598 3554
rect 81442 3502 81454 3554
rect 81506 3502 81518 3554
rect 85362 3502 85374 3554
rect 85426 3502 85438 3554
rect 89282 3502 89294 3554
rect 89346 3502 89358 3554
rect 93202 3502 93214 3554
rect 93266 3502 93278 3554
rect 97234 3502 97246 3554
rect 97298 3502 97310 3554
rect 101266 3502 101278 3554
rect 101330 3502 101342 3554
rect 105298 3502 105310 3554
rect 105362 3502 105374 3554
rect 109218 3502 109230 3554
rect 109282 3502 109294 3554
rect 113362 3502 113374 3554
rect 113426 3502 113438 3554
rect 117170 3502 117182 3554
rect 117234 3502 117246 3554
rect 121426 3502 121438 3554
rect 121490 3502 121502 3554
rect 125234 3502 125246 3554
rect 125298 3502 125310 3554
rect 126130 3502 126142 3554
rect 126194 3502 126206 3554
rect 129490 3502 129502 3554
rect 129554 3502 129566 3554
rect 133298 3502 133310 3554
rect 133362 3502 133374 3554
rect 137554 3502 137566 3554
rect 137618 3502 137630 3554
rect 140354 3502 140366 3554
rect 140418 3502 140430 3554
rect 144386 3502 144398 3554
rect 144450 3502 144462 3554
rect 71710 3490 71762 3502
rect 82910 3490 82962 3502
rect 98702 3490 98754 3502
rect 118302 3490 118354 3502
rect 131070 3490 131122 3502
rect 6302 3442 6354 3454
rect 6302 3378 6354 3390
rect 9998 3442 10050 3454
rect 9998 3378 10050 3390
rect 10334 3442 10386 3454
rect 10334 3378 10386 3390
rect 10894 3442 10946 3454
rect 10894 3378 10946 3390
rect 11678 3442 11730 3454
rect 15934 3442 15986 3454
rect 14354 3390 14366 3442
rect 14418 3390 14430 3442
rect 11678 3378 11730 3390
rect 15934 3378 15986 3390
rect 18846 3442 18898 3454
rect 18846 3378 18898 3390
rect 22990 3442 23042 3454
rect 22990 3378 23042 3390
rect 23438 3442 23490 3454
rect 27470 3442 27522 3454
rect 25666 3390 25678 3442
rect 25730 3390 25742 3442
rect 23438 3378 23490 3390
rect 27470 3378 27522 3390
rect 28590 3442 28642 3454
rect 28590 3378 28642 3390
rect 29598 3442 29650 3454
rect 31950 3442 32002 3454
rect 30482 3390 30494 3442
rect 30546 3390 30558 3442
rect 29598 3378 29650 3390
rect 31950 3378 32002 3390
rect 33182 3442 33234 3454
rect 33182 3378 33234 3390
rect 34190 3442 34242 3454
rect 34190 3378 34242 3390
rect 37102 3442 37154 3454
rect 37102 3378 37154 3390
rect 38446 3442 38498 3454
rect 44942 3442 44994 3454
rect 39330 3390 39342 3442
rect 39394 3390 39406 3442
rect 38446 3378 38498 3390
rect 44942 3378 44994 3390
rect 48974 3442 49026 3454
rect 48974 3378 49026 3390
rect 49870 3442 49922 3454
rect 49870 3378 49922 3390
rect 50318 3442 50370 3454
rect 50318 3378 50370 3390
rect 51214 3442 51266 3454
rect 51214 3378 51266 3390
rect 53342 3442 53394 3454
rect 62750 3442 62802 3454
rect 54002 3390 54014 3442
rect 54066 3390 54078 3442
rect 54562 3390 54574 3442
rect 54626 3390 54638 3442
rect 57026 3390 57038 3442
rect 57090 3390 57102 3442
rect 60946 3390 60958 3442
rect 61010 3390 61022 3442
rect 53342 3378 53394 3390
rect 62750 3378 62802 3390
rect 63310 3442 63362 3454
rect 74510 3442 74562 3454
rect 64866 3390 64878 3442
rect 64930 3390 64942 3442
rect 68786 3390 68798 3442
rect 68850 3390 68862 3442
rect 72706 3390 72718 3442
rect 72770 3390 72782 3442
rect 63310 3378 63362 3390
rect 74510 3378 74562 3390
rect 74958 3442 75010 3454
rect 78430 3442 78482 3454
rect 76626 3390 76638 3442
rect 76690 3390 76702 3442
rect 74958 3378 75010 3390
rect 78430 3378 78482 3390
rect 79326 3442 79378 3454
rect 82014 3442 82066 3454
rect 80546 3390 80558 3442
rect 80610 3390 80622 3442
rect 79326 3378 79378 3390
rect 82014 3378 82066 3390
rect 82350 3442 82402 3454
rect 86270 3442 86322 3454
rect 84466 3390 84478 3442
rect 84530 3390 84542 3442
rect 82350 3378 82402 3390
rect 86270 3378 86322 3390
rect 86718 3442 86770 3454
rect 90190 3442 90242 3454
rect 88386 3390 88398 3442
rect 88450 3390 88462 3442
rect 86718 3378 86770 3390
rect 90190 3378 90242 3390
rect 90638 3442 90690 3454
rect 93774 3442 93826 3454
rect 97806 3442 97858 3454
rect 101838 3442 101890 3454
rect 106206 3442 106258 3454
rect 92306 3390 92318 3442
rect 92370 3390 92382 3442
rect 96338 3390 96350 3442
rect 96402 3390 96414 3442
rect 100370 3390 100382 3442
rect 100434 3390 100446 3442
rect 104402 3390 104414 3442
rect 104466 3390 104478 3442
rect 90638 3378 90690 3390
rect 93774 3378 93826 3390
rect 97806 3378 97858 3390
rect 101838 3378 101890 3390
rect 106206 3378 106258 3390
rect 106654 3442 106706 3454
rect 109902 3442 109954 3454
rect 108994 3390 109006 3442
rect 109058 3390 109070 3442
rect 106654 3378 106706 3390
rect 109902 3378 109954 3390
rect 111470 3442 111522 3454
rect 111470 3378 111522 3390
rect 113934 3442 113986 3454
rect 121998 3442 122050 3454
rect 130062 3442 130114 3454
rect 116498 3390 116510 3442
rect 116562 3390 116574 3442
rect 120530 3390 120542 3442
rect 120594 3390 120606 3442
rect 124562 3390 124574 3442
rect 124626 3390 124638 3442
rect 128594 3390 128606 3442
rect 128658 3390 128670 3442
rect 132626 3390 132638 3442
rect 132690 3390 132702 3442
rect 136658 3390 136670 3442
rect 136722 3390 136734 3442
rect 141250 3390 141262 3442
rect 141314 3390 141326 3442
rect 145282 3390 145294 3442
rect 145346 3390 145358 3442
rect 113934 3378 113986 3390
rect 121998 3378 122050 3390
rect 130062 3378 130114 3390
rect 6638 3330 6690 3342
rect 6638 3266 6690 3278
rect 7534 3330 7586 3342
rect 7534 3266 7586 3278
rect 11342 3330 11394 3342
rect 11342 3266 11394 3278
rect 16718 3330 16770 3342
rect 16718 3266 16770 3278
rect 22094 3330 22146 3342
rect 22094 3266 22146 3278
rect 23774 3330 23826 3342
rect 23774 3266 23826 3278
rect 27806 3330 27858 3342
rect 27806 3266 27858 3278
rect 29262 3330 29314 3342
rect 29262 3266 29314 3278
rect 32286 3330 32338 3342
rect 32286 3266 32338 3278
rect 33518 3330 33570 3342
rect 33518 3266 33570 3278
rect 34526 3330 34578 3342
rect 34526 3266 34578 3278
rect 37438 3330 37490 3342
rect 37438 3266 37490 3278
rect 38110 3330 38162 3342
rect 38110 3266 38162 3278
rect 41022 3330 41074 3342
rect 41022 3266 41074 3278
rect 42030 3330 42082 3342
rect 42030 3266 42082 3278
rect 45278 3330 45330 3342
rect 45278 3266 45330 3278
rect 45950 3330 46002 3342
rect 45950 3266 46002 3278
rect 49310 3330 49362 3342
rect 49310 3266 49362 3278
rect 50654 3330 50706 3342
rect 50654 3266 50706 3278
rect 51662 3330 51714 3342
rect 51662 3266 51714 3278
rect 53006 3330 53058 3342
rect 53006 3266 53058 3278
rect 58606 3330 58658 3342
rect 58606 3266 58658 3278
rect 59502 3330 59554 3342
rect 59502 3266 59554 3278
rect 66334 3330 66386 3342
rect 66334 3266 66386 3278
rect 67230 3330 67282 3342
rect 67230 3266 67282 3278
rect 74174 3330 74226 3342
rect 74174 3266 74226 3278
rect 78094 3330 78146 3342
rect 78094 3266 78146 3278
rect 85934 3330 85986 3342
rect 85934 3266 85986 3278
rect 89854 3330 89906 3342
rect 89854 3266 89906 3278
rect 94110 3330 94162 3342
rect 94110 3266 94162 3278
rect 98142 3330 98194 3342
rect 98142 3266 98194 3278
rect 102174 3330 102226 3342
rect 102174 3266 102226 3278
rect 105870 3330 105922 3342
rect 105870 3266 105922 3278
rect 110238 3330 110290 3342
rect 110238 3266 110290 3278
rect 114270 3330 114322 3342
rect 114270 3266 114322 3278
rect 117966 3330 118018 3342
rect 117966 3266 118018 3278
rect 122334 3330 122386 3342
rect 122334 3266 122386 3278
rect 126366 3330 126418 3342
rect 126366 3266 126418 3278
rect 130398 3330 130450 3342
rect 130398 3266 130450 3278
rect 1344 3162 148784 3196
rect 1344 3110 38034 3162
rect 38086 3110 38138 3162
rect 38190 3110 38242 3162
rect 38294 3110 74854 3162
rect 74906 3110 74958 3162
rect 75010 3110 75062 3162
rect 75114 3110 111674 3162
rect 111726 3110 111778 3162
rect 111830 3110 111882 3162
rect 111934 3110 148494 3162
rect 148546 3110 148598 3162
rect 148650 3110 148702 3162
rect 148754 3110 148784 3162
rect 1344 3076 148784 3110
rect 105858 2942 105870 2994
rect 105922 2991 105934 2994
rect 106866 2991 106878 2994
rect 105922 2945 106878 2991
rect 105922 2942 105934 2945
rect 106866 2942 106878 2945
rect 106930 2942 106942 2994
<< via1 >>
rect 19624 36822 19676 36874
rect 19728 36822 19780 36874
rect 19832 36822 19884 36874
rect 56444 36822 56496 36874
rect 56548 36822 56600 36874
rect 56652 36822 56704 36874
rect 93264 36822 93316 36874
rect 93368 36822 93420 36874
rect 93472 36822 93524 36874
rect 130084 36822 130136 36874
rect 130188 36822 130240 36874
rect 130292 36822 130344 36874
rect 30158 36654 30210 36706
rect 35982 36654 36034 36706
rect 36542 36654 36594 36706
rect 75070 36654 75122 36706
rect 132414 36654 132466 36706
rect 5966 36542 6018 36594
rect 8206 36542 8258 36594
rect 10446 36542 10498 36594
rect 12126 36542 12178 36594
rect 14478 36542 14530 36594
rect 16046 36542 16098 36594
rect 22206 36542 22258 36594
rect 23886 36542 23938 36594
rect 26014 36542 26066 36594
rect 27806 36542 27858 36594
rect 31502 36542 31554 36594
rect 34638 36542 34690 36594
rect 36094 36542 36146 36594
rect 37774 36542 37826 36594
rect 39566 36542 39618 36594
rect 41358 36542 41410 36594
rect 43150 36542 43202 36594
rect 49534 36542 49586 36594
rect 51326 36542 51378 36594
rect 54910 36542 54962 36594
rect 57934 36542 57986 36594
rect 61070 36542 61122 36594
rect 64542 36542 64594 36594
rect 68910 36542 68962 36594
rect 70590 36542 70642 36594
rect 73390 36542 73442 36594
rect 80894 36542 80946 36594
rect 82686 36542 82738 36594
rect 84814 36542 84866 36594
rect 86158 36542 86210 36594
rect 96574 36542 96626 36594
rect 98366 36542 98418 36594
rect 100046 36542 100098 36594
rect 102398 36542 102450 36594
rect 104414 36542 104466 36594
rect 112254 36542 112306 36594
rect 114046 36542 114098 36594
rect 116622 36542 116674 36594
rect 120206 36542 120258 36594
rect 121998 36542 122050 36594
rect 126030 36542 126082 36594
rect 127934 36542 127986 36594
rect 129726 36542 129778 36594
rect 133758 36542 133810 36594
rect 141598 36542 141650 36594
rect 143614 36542 143666 36594
rect 145406 36542 145458 36594
rect 6974 36430 7026 36482
rect 7646 36430 7698 36482
rect 9774 36430 9826 36482
rect 12574 36430 12626 36482
rect 13918 36430 13970 36482
rect 16718 36430 16770 36482
rect 18062 36430 18114 36482
rect 19742 36430 19794 36482
rect 21758 36430 21810 36482
rect 24446 36430 24498 36482
rect 26462 36430 26514 36482
rect 28478 36430 28530 36482
rect 32174 36430 32226 36482
rect 33518 36430 33570 36482
rect 35534 36430 35586 36482
rect 38446 36430 38498 36482
rect 40238 36430 40290 36482
rect 42366 36430 42418 36482
rect 44158 36430 44210 36482
rect 45726 36430 45778 36482
rect 47518 36430 47570 36482
rect 48974 36430 49026 36482
rect 51998 36430 52050 36482
rect 53006 36430 53058 36482
rect 53678 36430 53730 36482
rect 55918 36430 55970 36482
rect 58830 36430 58882 36482
rect 61742 36430 61794 36482
rect 62750 36430 62802 36482
rect 63310 36430 63362 36482
rect 64990 36430 65042 36482
rect 66110 36430 66162 36482
rect 66782 36430 66834 36482
rect 69694 36430 69746 36482
rect 71486 36430 71538 36482
rect 72382 36430 72434 36482
rect 74398 36430 74450 36482
rect 76750 36430 76802 36482
rect 77422 36430 77474 36482
rect 80446 36430 80498 36482
rect 82014 36430 82066 36482
rect 84142 36430 84194 36482
rect 86942 36430 86994 36482
rect 87950 36430 88002 36482
rect 88958 36430 89010 36482
rect 89742 36430 89794 36482
rect 92206 36430 92258 36482
rect 93662 36430 93714 36482
rect 94334 36430 94386 36482
rect 96126 36430 96178 36482
rect 97918 36430 97970 36482
rect 100830 36430 100882 36482
rect 101614 36430 101666 36482
rect 103742 36430 103794 36482
rect 106430 36430 106482 36482
rect 108670 36430 108722 36482
rect 109342 36430 109394 36482
rect 111582 36430 111634 36482
rect 113374 36430 113426 36482
rect 115950 36430 116002 36482
rect 117854 36430 117906 36482
rect 119534 36430 119586 36482
rect 121326 36430 121378 36482
rect 123790 36430 123842 36482
rect 124574 36430 124626 36482
rect 125246 36430 125298 36482
rect 127262 36430 127314 36482
rect 129278 36430 129330 36482
rect 131406 36430 131458 36482
rect 132078 36430 132130 36482
rect 133086 36430 133138 36482
rect 136558 36430 136610 36482
rect 137790 36430 137842 36482
rect 139246 36430 139298 36482
rect 139918 36430 139970 36482
rect 141038 36430 141090 36482
rect 142942 36430 142994 36482
rect 144958 36430 145010 36482
rect 4846 36318 4898 36370
rect 17502 36318 17554 36370
rect 18958 36318 19010 36370
rect 19518 36318 19570 36370
rect 29486 36318 29538 36370
rect 29822 36318 29874 36370
rect 33854 36318 33906 36370
rect 46846 36318 46898 36370
rect 47182 36318 47234 36370
rect 52894 36318 52946 36370
rect 56814 36318 56866 36370
rect 57150 36318 57202 36370
rect 59502 36318 59554 36370
rect 62526 36318 62578 36370
rect 65326 36318 65378 36370
rect 65998 36318 66050 36370
rect 67790 36318 67842 36370
rect 74286 36318 74338 36370
rect 76638 36318 76690 36370
rect 78766 36318 78818 36370
rect 89518 36318 89570 36370
rect 90750 36318 90802 36370
rect 91198 36318 91250 36370
rect 91982 36318 92034 36370
rect 93774 36318 93826 36370
rect 105646 36318 105698 36370
rect 106206 36318 106258 36370
rect 108558 36318 108610 36370
rect 110350 36318 110402 36370
rect 110686 36318 110738 36370
rect 118078 36318 118130 36370
rect 124350 36318 124402 36370
rect 131294 36318 131346 36370
rect 135774 36318 135826 36370
rect 136222 36318 136274 36370
rect 139134 36318 139186 36370
rect 18286 36206 18338 36258
rect 20078 36206 20130 36258
rect 20750 36206 20802 36258
rect 30494 36206 30546 36258
rect 45278 36206 45330 36258
rect 46062 36206 46114 36258
rect 47854 36206 47906 36258
rect 54014 36206 54066 36258
rect 59838 36206 59890 36258
rect 63646 36206 63698 36258
rect 67118 36206 67170 36258
rect 75406 36206 75458 36258
rect 77758 36206 77810 36258
rect 78430 36206 78482 36258
rect 79214 36206 79266 36258
rect 88622 36206 88674 36258
rect 90414 36206 90466 36258
rect 92766 36206 92818 36258
rect 94670 36206 94722 36258
rect 106766 36206 106818 36258
rect 107550 36206 107602 36258
rect 109678 36206 109730 36258
rect 115502 36206 115554 36258
rect 118526 36206 118578 36258
rect 123454 36206 123506 36258
rect 134990 36206 135042 36258
rect 136894 36206 136946 36258
rect 137566 36206 137618 36258
rect 140254 36206 140306 36258
rect 38034 36038 38086 36090
rect 38138 36038 38190 36090
rect 38242 36038 38294 36090
rect 74854 36038 74906 36090
rect 74958 36038 75010 36090
rect 75062 36038 75114 36090
rect 111674 36038 111726 36090
rect 111778 36038 111830 36090
rect 111882 36038 111934 36090
rect 148494 36038 148546 36090
rect 148598 36038 148650 36090
rect 148702 36038 148754 36090
rect 6078 35870 6130 35922
rect 8990 35870 9042 35922
rect 19518 35870 19570 35922
rect 23102 35870 23154 35922
rect 26574 35870 26626 35922
rect 39006 35870 39058 35922
rect 41806 35870 41858 35922
rect 42366 35870 42418 35922
rect 43262 35870 43314 35922
rect 54574 35870 54626 35922
rect 57598 35870 57650 35922
rect 58942 35870 58994 35922
rect 61294 35870 61346 35922
rect 64542 35870 64594 35922
rect 70814 35870 70866 35922
rect 73950 35870 74002 35922
rect 80334 35870 80386 35922
rect 92990 35870 93042 35922
rect 97246 35870 97298 35922
rect 99822 35870 99874 35922
rect 100606 35870 100658 35922
rect 101166 35870 101218 35922
rect 104190 35870 104242 35922
rect 111358 35870 111410 35922
rect 113150 35870 113202 35922
rect 116846 35870 116898 35922
rect 119870 35870 119922 35922
rect 121102 35870 121154 35922
rect 122334 35870 122386 35922
rect 132974 35870 133026 35922
rect 137902 35870 137954 35922
rect 142158 35870 142210 35922
rect 144958 35870 145010 35922
rect 145854 35870 145906 35922
rect 146638 35870 146690 35922
rect 7534 35758 7586 35810
rect 10558 35758 10610 35810
rect 13246 35758 13298 35810
rect 17838 35758 17890 35810
rect 20414 35758 20466 35810
rect 30158 35758 30210 35810
rect 34526 35758 34578 35810
rect 36542 35758 36594 35810
rect 39902 35758 39954 35810
rect 40798 35758 40850 35810
rect 43934 35758 43986 35810
rect 44382 35758 44434 35810
rect 46398 35758 46450 35810
rect 50318 35758 50370 35810
rect 51886 35758 51938 35810
rect 52446 35758 52498 35810
rect 53678 35758 53730 35810
rect 54014 35758 54066 35810
rect 55806 35758 55858 35810
rect 58606 35758 58658 35810
rect 62414 35758 62466 35810
rect 64206 35758 64258 35810
rect 65774 35758 65826 35810
rect 67902 35758 67954 35810
rect 69918 35758 69970 35810
rect 70478 35758 70530 35810
rect 74734 35758 74786 35810
rect 76862 35758 76914 35810
rect 83470 35758 83522 35810
rect 86382 35758 86434 35810
rect 89406 35758 89458 35810
rect 89966 35758 90018 35810
rect 93662 35758 93714 35810
rect 95342 35758 95394 35810
rect 101614 35758 101666 35810
rect 102846 35758 102898 35810
rect 105534 35758 105586 35810
rect 106318 35758 106370 35810
rect 108334 35758 108386 35810
rect 109342 35758 109394 35810
rect 112254 35758 112306 35810
rect 116286 35758 116338 35810
rect 124462 35758 124514 35810
rect 126254 35758 126306 35810
rect 129614 35758 129666 35810
rect 130846 35758 130898 35810
rect 131406 35758 131458 35810
rect 134766 35758 134818 35810
rect 135662 35758 135714 35810
rect 138686 35758 138738 35810
rect 140590 35758 140642 35810
rect 143726 35758 143778 35810
rect 146190 35758 146242 35810
rect 6638 35646 6690 35698
rect 8766 35646 8818 35698
rect 10334 35646 10386 35698
rect 11118 35646 11170 35698
rect 13022 35646 13074 35698
rect 13806 35646 13858 35698
rect 15934 35646 15986 35698
rect 18174 35646 18226 35698
rect 20078 35646 20130 35698
rect 20974 35646 21026 35698
rect 22878 35646 22930 35698
rect 23662 35646 23714 35698
rect 26238 35646 26290 35698
rect 28142 35646 28194 35698
rect 29374 35646 29426 35698
rect 29822 35646 29874 35698
rect 30830 35646 30882 35698
rect 33630 35646 33682 35698
rect 37438 35646 37490 35698
rect 38670 35646 38722 35698
rect 39566 35646 39618 35698
rect 40574 35646 40626 35698
rect 42702 35646 42754 35698
rect 46174 35646 46226 35698
rect 46958 35646 47010 35698
rect 51214 35646 51266 35698
rect 52670 35646 52722 35698
rect 54910 35646 54962 35698
rect 56702 35646 56754 35698
rect 57822 35646 57874 35698
rect 60734 35646 60786 35698
rect 61518 35646 61570 35698
rect 62750 35646 62802 35698
rect 66110 35646 66162 35698
rect 68798 35646 68850 35698
rect 69582 35646 69634 35698
rect 72606 35646 72658 35698
rect 73726 35646 73778 35698
rect 74622 35646 74674 35698
rect 76750 35646 76802 35698
rect 77534 35646 77586 35698
rect 78542 35646 78594 35698
rect 81342 35646 81394 35698
rect 83246 35646 83298 35698
rect 84590 35646 84642 35698
rect 86606 35646 86658 35698
rect 87390 35646 87442 35698
rect 90190 35646 90242 35698
rect 91198 35646 91250 35698
rect 93550 35646 93602 35698
rect 94334 35646 94386 35698
rect 95566 35646 95618 35698
rect 98030 35646 98082 35698
rect 100046 35646 100098 35698
rect 101838 35646 101890 35698
rect 103518 35646 103570 35698
rect 105198 35646 105250 35698
rect 106206 35646 106258 35698
rect 107998 35646 108050 35698
rect 109230 35646 109282 35698
rect 111022 35646 111074 35698
rect 112030 35646 112082 35698
rect 113486 35646 113538 35698
rect 114270 35646 114322 35698
rect 116062 35646 116114 35698
rect 117070 35646 117122 35698
rect 117742 35646 117794 35698
rect 119646 35646 119698 35698
rect 121326 35646 121378 35698
rect 121998 35646 122050 35698
rect 124574 35646 124626 35698
rect 125358 35646 125410 35698
rect 127934 35646 127986 35698
rect 129054 35646 129106 35698
rect 130062 35646 130114 35698
rect 132638 35646 132690 35698
rect 133870 35646 133922 35698
rect 135886 35646 135938 35698
rect 136894 35646 136946 35698
rect 137678 35646 137730 35698
rect 138574 35646 138626 35698
rect 140478 35646 140530 35698
rect 142830 35646 142882 35698
rect 145182 35646 145234 35698
rect 9662 35534 9714 35586
rect 11790 35534 11842 35586
rect 14478 35534 14530 35586
rect 16382 35534 16434 35586
rect 21646 35534 21698 35586
rect 24334 35534 24386 35586
rect 25678 35534 25730 35586
rect 27358 35534 27410 35586
rect 31502 35534 31554 35586
rect 32622 35534 32674 35586
rect 38110 35534 38162 35586
rect 45614 35534 45666 35586
rect 47630 35534 47682 35586
rect 48750 35534 48802 35586
rect 49422 35534 49474 35586
rect 59726 35534 59778 35586
rect 71822 35534 71874 35586
rect 79214 35534 79266 35586
rect 82014 35534 82066 35586
rect 83918 35534 83970 35586
rect 85262 35534 85314 35586
rect 87950 35534 88002 35586
rect 91870 35534 91922 35586
rect 96126 35534 96178 35586
rect 98702 35534 98754 35586
rect 107326 35534 107378 35586
rect 114830 35534 114882 35586
rect 118414 35534 118466 35586
rect 120318 35534 120370 35586
rect 122782 35534 122834 35586
rect 127374 35534 127426 35586
rect 131630 35534 131682 35586
rect 141262 35534 141314 35586
rect 18622 35422 18674 35474
rect 18958 35422 19010 35474
rect 29038 35422 29090 35474
rect 44606 35422 44658 35474
rect 44942 35422 44994 35474
rect 53006 35422 53058 35474
rect 63198 35422 63250 35474
rect 63534 35422 63586 35474
rect 66558 35422 66610 35474
rect 66894 35422 66946 35474
rect 75406 35422 75458 35474
rect 75742 35422 75794 35474
rect 77870 35422 77922 35474
rect 90526 35422 90578 35474
rect 94670 35422 94722 35474
rect 106990 35422 107042 35474
rect 110014 35422 110066 35474
rect 110350 35422 110402 35474
rect 123566 35422 123618 35474
rect 123902 35422 123954 35474
rect 131966 35422 132018 35474
rect 139358 35422 139410 35474
rect 139694 35422 139746 35474
rect 141598 35422 141650 35474
rect 19624 35254 19676 35306
rect 19728 35254 19780 35306
rect 19832 35254 19884 35306
rect 56444 35254 56496 35306
rect 56548 35254 56600 35306
rect 56652 35254 56704 35306
rect 93264 35254 93316 35306
rect 93368 35254 93420 35306
rect 93472 35254 93524 35306
rect 130084 35254 130136 35306
rect 130188 35254 130240 35306
rect 130292 35254 130344 35306
rect 53790 35086 53842 35138
rect 10110 34974 10162 35026
rect 11006 34974 11058 35026
rect 18510 34974 18562 35026
rect 20302 34974 20354 35026
rect 31390 34974 31442 35026
rect 42030 34974 42082 35026
rect 43374 34974 43426 35026
rect 43822 34974 43874 35026
rect 45726 34974 45778 35026
rect 53454 34974 53506 35026
rect 56030 34974 56082 35026
rect 59614 34974 59666 35026
rect 63422 34974 63474 35026
rect 65102 34974 65154 35026
rect 66670 34974 66722 35026
rect 68686 34974 68738 35026
rect 70142 34974 70194 35026
rect 71038 34974 71090 35026
rect 71598 34974 71650 35026
rect 72046 34974 72098 35026
rect 72494 34974 72546 35026
rect 77982 34974 78034 35026
rect 82574 34974 82626 35026
rect 88846 34974 88898 35026
rect 90190 34974 90242 35026
rect 93998 34974 94050 35026
rect 96014 34974 96066 35026
rect 99598 34974 99650 35026
rect 103854 34974 103906 35026
rect 105870 34974 105922 35026
rect 107662 34974 107714 35026
rect 109790 34974 109842 35026
rect 117070 34974 117122 35026
rect 120430 34974 120482 35026
rect 120990 34974 121042 35026
rect 131070 34974 131122 35026
rect 136334 34974 136386 35026
rect 138126 34974 138178 35026
rect 139134 34974 139186 35026
rect 145518 34974 145570 35026
rect 6190 34862 6242 34914
rect 6974 34862 7026 34914
rect 7870 34862 7922 34914
rect 8542 34862 8594 34914
rect 9326 34862 9378 34914
rect 11790 34862 11842 34914
rect 12910 34862 12962 34914
rect 13582 34862 13634 34914
rect 14590 34862 14642 34914
rect 15262 34862 15314 34914
rect 17166 34862 17218 34914
rect 18062 34862 18114 34914
rect 19630 34862 19682 34914
rect 22766 34862 22818 34914
rect 23998 34862 24050 34914
rect 25454 34862 25506 34914
rect 29934 34862 29986 34914
rect 30606 34862 30658 34914
rect 32846 34862 32898 34914
rect 36542 34862 36594 34914
rect 37774 34862 37826 34914
rect 38334 34862 38386 34914
rect 40126 34862 40178 34914
rect 42478 34862 42530 34914
rect 44270 34862 44322 34914
rect 46622 34862 46674 34914
rect 49534 34862 49586 34914
rect 50654 34862 50706 34914
rect 54574 34862 54626 34914
rect 55022 34862 55074 34914
rect 57374 34862 57426 34914
rect 58606 34862 58658 34914
rect 62190 34862 62242 34914
rect 64318 34862 64370 34914
rect 66110 34862 66162 34914
rect 67118 34862 67170 34914
rect 67566 34862 67618 34914
rect 69358 34862 69410 34914
rect 72942 34862 72994 34914
rect 73838 34862 73890 34914
rect 74734 34862 74786 34914
rect 75854 34862 75906 34914
rect 76190 34862 76242 34914
rect 77310 34862 77362 34914
rect 79550 34862 79602 34914
rect 81902 34862 81954 34914
rect 88174 34862 88226 34914
rect 90974 34862 91026 34914
rect 93438 34862 93490 34914
rect 95342 34862 95394 34914
rect 97358 34862 97410 34914
rect 104526 34862 104578 34914
rect 105198 34862 105250 34914
rect 106990 34862 107042 34914
rect 109230 34862 109282 34914
rect 111694 34862 111746 34914
rect 115278 34862 115330 34914
rect 117854 34862 117906 34914
rect 119870 34862 119922 34914
rect 122670 34862 122722 34914
rect 125246 34862 125298 34914
rect 127038 34862 127090 34914
rect 128830 34862 128882 34914
rect 129390 34862 129442 34914
rect 130510 34862 130562 34914
rect 131966 34862 132018 34914
rect 133198 34862 133250 34914
rect 135774 34862 135826 34914
rect 137454 34862 137506 34914
rect 140030 34862 140082 34914
rect 140926 34862 140978 34914
rect 143950 34862 144002 34914
rect 6638 34750 6690 34802
rect 7534 34750 7586 34802
rect 8766 34750 8818 34802
rect 12014 34750 12066 34802
rect 12574 34750 12626 34802
rect 14254 34750 14306 34802
rect 16046 34750 16098 34802
rect 16382 34750 16434 34802
rect 16942 34750 16994 34802
rect 21870 34750 21922 34802
rect 22206 34750 22258 34802
rect 23102 34750 23154 34802
rect 23662 34750 23714 34802
rect 24558 34750 24610 34802
rect 24894 34750 24946 34802
rect 25790 34750 25842 34802
rect 26574 34750 26626 34802
rect 26910 34750 26962 34802
rect 27806 34750 27858 34802
rect 28142 34750 28194 34802
rect 29598 34750 29650 34802
rect 30830 34750 30882 34802
rect 31838 34750 31890 34802
rect 32174 34750 32226 34802
rect 33630 34750 33682 34802
rect 33966 34750 34018 34802
rect 34526 34750 34578 34802
rect 35534 34750 35586 34802
rect 35870 34750 35922 34802
rect 39118 34750 39170 34802
rect 39454 34750 39506 34802
rect 40910 34750 40962 34802
rect 41246 34750 41298 34802
rect 47742 34750 47794 34802
rect 48638 34750 48690 34802
rect 48974 34750 49026 34802
rect 51438 34750 51490 34802
rect 51774 34750 51826 34802
rect 52334 34750 52386 34802
rect 54014 34750 54066 34802
rect 56478 34750 56530 34802
rect 60062 34750 60114 34802
rect 73278 34750 73330 34802
rect 84030 34750 84082 34802
rect 85262 34750 85314 34802
rect 85598 34750 85650 34802
rect 86942 34750 86994 34802
rect 87278 34750 87330 34802
rect 92430 34750 92482 34802
rect 102398 34750 102450 34802
rect 102958 34750 103010 34802
rect 103294 34750 103346 34802
rect 111470 34750 111522 34802
rect 113150 34750 113202 34802
rect 114382 34750 114434 34802
rect 115838 34750 115890 34802
rect 118750 34750 118802 34802
rect 119086 34750 119138 34802
rect 121550 34750 121602 34802
rect 121886 34750 121938 34802
rect 122446 34750 122498 34802
rect 123342 34750 123394 34802
rect 123678 34750 123730 34802
rect 126254 34750 126306 34802
rect 127710 34750 127762 34802
rect 128046 34750 128098 34802
rect 132974 34750 133026 34802
rect 134430 34750 134482 34802
rect 139806 34750 139858 34802
rect 141262 34750 141314 34802
rect 142158 34750 142210 34802
rect 142494 34750 142546 34802
rect 142942 34750 142994 34802
rect 15486 34638 15538 34690
rect 28702 34638 28754 34690
rect 33070 34638 33122 34690
rect 34862 34638 34914 34690
rect 36766 34638 36818 34690
rect 38558 34638 38610 34690
rect 40350 34638 40402 34690
rect 42814 34638 42866 34690
rect 44606 34638 44658 34690
rect 47294 34638 47346 34690
rect 48078 34638 48130 34690
rect 49870 34638 49922 34690
rect 50878 34638 50930 34690
rect 52670 34638 52722 34690
rect 55358 34638 55410 34690
rect 56814 34638 56866 34690
rect 57710 34638 57762 34690
rect 58942 34638 58994 34690
rect 60622 34638 60674 34690
rect 61630 34638 61682 34690
rect 62526 34638 62578 34690
rect 67902 34638 67954 34690
rect 69694 34638 69746 34690
rect 74174 34638 74226 34690
rect 75294 34638 75346 34690
rect 75966 34638 76018 34690
rect 76638 34638 76690 34690
rect 79774 34638 79826 34690
rect 80222 34638 80274 34690
rect 80670 34638 80722 34690
rect 81342 34638 81394 34690
rect 83694 34638 83746 34690
rect 84590 34638 84642 34690
rect 86158 34638 86210 34690
rect 92094 34638 92146 34690
rect 97134 34638 97186 34690
rect 98030 34638 98082 34690
rect 98366 34638 98418 34690
rect 101166 34638 101218 34690
rect 101614 34638 101666 34690
rect 102062 34638 102114 34690
rect 104302 34638 104354 34690
rect 110798 34638 110850 34690
rect 112254 34638 112306 34690
rect 113486 34638 113538 34690
rect 114046 34638 114098 34690
rect 115054 34638 115106 34690
rect 116286 34638 116338 34690
rect 118190 34638 118242 34690
rect 119646 34638 119698 34690
rect 124238 34638 124290 34690
rect 125022 34638 125074 34690
rect 125918 34638 125970 34690
rect 126814 34638 126866 34690
rect 128606 34638 128658 34690
rect 133758 34638 133810 34690
rect 134766 34638 134818 34690
rect 143726 34638 143778 34690
rect 38034 34470 38086 34522
rect 38138 34470 38190 34522
rect 38242 34470 38294 34522
rect 74854 34470 74906 34522
rect 74958 34470 75010 34522
rect 75062 34470 75114 34522
rect 111674 34470 111726 34522
rect 111778 34470 111830 34522
rect 111882 34470 111934 34522
rect 148494 34470 148546 34522
rect 148598 34470 148650 34522
rect 148702 34470 148754 34522
rect 7534 34302 7586 34354
rect 7982 34302 8034 34354
rect 9662 34302 9714 34354
rect 12238 34302 12290 34354
rect 14814 34302 14866 34354
rect 15710 34302 15762 34354
rect 18062 34302 18114 34354
rect 19518 34302 19570 34354
rect 20974 34302 21026 34354
rect 22878 34302 22930 34354
rect 23326 34302 23378 34354
rect 24222 34302 24274 34354
rect 26014 34302 26066 34354
rect 27694 34302 27746 34354
rect 28478 34302 28530 34354
rect 29038 34302 29090 34354
rect 29374 34302 29426 34354
rect 29822 34302 29874 34354
rect 30382 34302 30434 34354
rect 31726 34302 31778 34354
rect 33518 34302 33570 34354
rect 36878 34302 36930 34354
rect 37438 34302 37490 34354
rect 40574 34302 40626 34354
rect 46622 34302 46674 34354
rect 48862 34302 48914 34354
rect 49982 34302 50034 34354
rect 50878 34302 50930 34354
rect 51662 34302 51714 34354
rect 52222 34302 52274 34354
rect 54238 34302 54290 34354
rect 54798 34302 54850 34354
rect 56590 34302 56642 34354
rect 57486 34302 57538 34354
rect 58382 34302 58434 34354
rect 59278 34302 59330 34354
rect 62638 34302 62690 34354
rect 63870 34302 63922 34354
rect 64654 34302 64706 34354
rect 65438 34302 65490 34354
rect 67902 34302 67954 34354
rect 73278 34302 73330 34354
rect 73950 34302 74002 34354
rect 74398 34302 74450 34354
rect 75182 34302 75234 34354
rect 75630 34302 75682 34354
rect 76190 34302 76242 34354
rect 76750 34302 76802 34354
rect 78206 34302 78258 34354
rect 78766 34302 78818 34354
rect 81342 34302 81394 34354
rect 81790 34302 81842 34354
rect 82350 34302 82402 34354
rect 83918 34302 83970 34354
rect 84366 34302 84418 34354
rect 86158 34302 86210 34354
rect 87390 34302 87442 34354
rect 87950 34302 88002 34354
rect 89294 34302 89346 34354
rect 90862 34302 90914 34354
rect 93438 34302 93490 34354
rect 95566 34302 95618 34354
rect 96350 34302 96402 34354
rect 97246 34302 97298 34354
rect 103518 34302 103570 34354
rect 105646 34302 105698 34354
rect 107326 34302 107378 34354
rect 108782 34302 108834 34354
rect 109230 34302 109282 34354
rect 111246 34302 111298 34354
rect 114942 34302 114994 34354
rect 117518 34302 117570 34354
rect 122670 34302 122722 34354
rect 123006 34302 123058 34354
rect 124798 34302 124850 34354
rect 125134 34302 125186 34354
rect 127822 34302 127874 34354
rect 129390 34302 129442 34354
rect 130286 34302 130338 34354
rect 131742 34302 131794 34354
rect 132526 34302 132578 34354
rect 132974 34302 133026 34354
rect 135214 34302 135266 34354
rect 135662 34302 135714 34354
rect 137342 34302 137394 34354
rect 138910 34302 138962 34354
rect 139358 34302 139410 34354
rect 140366 34302 140418 34354
rect 140814 34302 140866 34354
rect 141486 34302 141538 34354
rect 141934 34302 141986 34354
rect 143502 34302 143554 34354
rect 8430 34190 8482 34242
rect 8766 34190 8818 34242
rect 19182 34190 19234 34242
rect 20078 34190 20130 34242
rect 20414 34190 20466 34242
rect 28142 34190 28194 34242
rect 30830 34190 30882 34242
rect 31166 34190 31218 34242
rect 39454 34190 39506 34242
rect 46062 34190 46114 34242
rect 49646 34190 49698 34242
rect 52558 34190 52610 34242
rect 53118 34190 53170 34242
rect 53454 34190 53506 34242
rect 73838 34190 73890 34242
rect 79214 34190 79266 34242
rect 82798 34190 82850 34242
rect 83134 34190 83186 34242
rect 89854 34190 89906 34242
rect 92654 34190 92706 34242
rect 106094 34190 106146 34242
rect 106430 34190 106482 34242
rect 107886 34190 107938 34242
rect 109678 34190 109730 34242
rect 113598 34190 113650 34242
rect 126142 34190 126194 34242
rect 130846 34190 130898 34242
rect 131182 34190 131234 34242
rect 132078 34190 132130 34242
rect 138350 34190 138402 34242
rect 142270 34190 142322 34242
rect 18398 34078 18450 34130
rect 21310 34078 21362 34130
rect 25566 34078 25618 34130
rect 37774 34078 37826 34130
rect 39118 34078 39170 34130
rect 44718 34078 44770 34130
rect 45838 34078 45890 34130
rect 46958 34078 47010 34130
rect 48190 34078 48242 34130
rect 61182 34078 61234 34130
rect 62302 34078 62354 34130
rect 79438 34078 79490 34130
rect 91758 34078 91810 34130
rect 106990 34078 107042 34130
rect 108110 34078 108162 34130
rect 109902 34078 109954 34130
rect 113934 34078 113986 34130
rect 125582 34078 125634 34130
rect 126478 34078 126530 34130
rect 129054 34078 129106 34130
rect 130062 34078 130114 34130
rect 13470 33966 13522 34018
rect 16494 33966 16546 34018
rect 17054 33966 17106 34018
rect 21758 33966 21810 34018
rect 22430 33966 22482 34018
rect 27134 33966 27186 34018
rect 32398 33966 32450 34018
rect 34190 33966 34242 34018
rect 35086 33966 35138 34018
rect 36094 33966 36146 34018
rect 38558 33966 38610 34018
rect 39902 33966 39954 34018
rect 41470 33966 41522 34018
rect 41918 33966 41970 34018
rect 42926 33966 42978 34018
rect 45278 33966 45330 34018
rect 47406 33966 47458 34018
rect 51214 33966 51266 34018
rect 55134 33966 55186 34018
rect 55806 33966 55858 34018
rect 56142 33966 56194 34018
rect 57822 33966 57874 34018
rect 58718 33966 58770 34018
rect 59838 33966 59890 34018
rect 60174 33966 60226 34018
rect 60622 33966 60674 34018
rect 61742 33966 61794 34018
rect 63310 33966 63362 34018
rect 65886 33966 65938 34018
rect 66446 33966 66498 34018
rect 67454 33966 67506 34018
rect 69022 33966 69074 34018
rect 72718 33966 72770 34018
rect 77198 33966 77250 34018
rect 86606 33966 86658 34018
rect 88510 33966 88562 34018
rect 90302 33966 90354 34018
rect 91198 33966 91250 34018
rect 93886 33966 93938 34018
rect 95118 33966 95170 34018
rect 96014 33966 96066 34018
rect 102622 33966 102674 34018
rect 104414 33966 104466 34018
rect 105198 33966 105250 34018
rect 110798 33966 110850 34018
rect 111582 33966 111634 34018
rect 113038 33966 113090 34018
rect 114382 33966 114434 34018
rect 119310 33966 119362 34018
rect 122110 33966 122162 34018
rect 123566 33966 123618 34018
rect 126926 33966 126978 34018
rect 127374 33966 127426 34018
rect 128270 33966 128322 34018
rect 134094 33966 134146 34018
rect 138014 33966 138066 34018
rect 139918 33966 139970 34018
rect 138014 33854 138066 33906
rect 138686 33854 138738 33906
rect 139918 33854 139970 33906
rect 140590 33854 140642 33906
rect 19624 33686 19676 33738
rect 19728 33686 19780 33738
rect 19832 33686 19884 33738
rect 56444 33686 56496 33738
rect 56548 33686 56600 33738
rect 56652 33686 56704 33738
rect 93264 33686 93316 33738
rect 93368 33686 93420 33738
rect 93472 33686 93524 33738
rect 130084 33686 130136 33738
rect 130188 33686 130240 33738
rect 130292 33686 130344 33738
rect 106654 33518 106706 33570
rect 106990 33518 107042 33570
rect 17502 33406 17554 33458
rect 18958 33406 19010 33458
rect 19294 33406 19346 33458
rect 19854 33406 19906 33458
rect 20638 33406 20690 33458
rect 30606 33406 30658 33458
rect 31054 33406 31106 33458
rect 46286 33406 46338 33458
rect 46846 33406 46898 33458
rect 49198 33406 49250 33458
rect 51998 33406 52050 33458
rect 53342 33406 53394 33458
rect 53902 33406 53954 33458
rect 59278 33406 59330 33458
rect 60286 33406 60338 33458
rect 61742 33406 61794 33458
rect 63086 33406 63138 33458
rect 64542 33406 64594 33458
rect 65102 33406 65154 33458
rect 65550 33406 65602 33458
rect 73838 33406 73890 33458
rect 74286 33406 74338 33458
rect 74622 33406 74674 33458
rect 87950 33406 88002 33458
rect 89070 33406 89122 33458
rect 91758 33406 91810 33458
rect 93214 33406 93266 33458
rect 105758 33406 105810 33458
rect 106206 33406 106258 33458
rect 107214 33406 107266 33458
rect 107662 33406 107714 33458
rect 109454 33406 109506 33458
rect 110126 33406 110178 33458
rect 126590 33406 126642 33458
rect 127038 33406 127090 33458
rect 128718 33406 128770 33458
rect 131070 33406 131122 33458
rect 131518 33406 131570 33458
rect 51550 33294 51602 33346
rect 52782 33294 52834 33346
rect 54462 33294 54514 33346
rect 62190 33294 62242 33346
rect 63758 33294 63810 33346
rect 129278 33294 129330 33346
rect 18398 33182 18450 33234
rect 89518 33182 89570 33234
rect 110910 33182 110962 33234
rect 129614 33182 129666 33234
rect 20302 33070 20354 33122
rect 37998 33070 38050 33122
rect 38446 33070 38498 33122
rect 60622 33070 60674 33122
rect 62526 33070 62578 33122
rect 64206 33070 64258 33122
rect 76078 33070 76130 33122
rect 105086 33070 105138 33122
rect 106654 33070 106706 33122
rect 107998 33070 108050 33122
rect 109118 33070 109170 33122
rect 130174 33070 130226 33122
rect 130510 33070 130562 33122
rect 38034 32902 38086 32954
rect 38138 32902 38190 32954
rect 38242 32902 38294 32954
rect 74854 32902 74906 32954
rect 74958 32902 75010 32954
rect 75062 32902 75114 32954
rect 111674 32902 111726 32954
rect 111778 32902 111830 32954
rect 111882 32902 111934 32954
rect 148494 32902 148546 32954
rect 148598 32902 148650 32954
rect 148702 32902 148754 32954
rect 53454 32734 53506 32786
rect 62078 32734 62130 32786
rect 62526 32734 62578 32786
rect 62974 32734 63026 32786
rect 108222 32734 108274 32786
rect 19624 32118 19676 32170
rect 19728 32118 19780 32170
rect 19832 32118 19884 32170
rect 56444 32118 56496 32170
rect 56548 32118 56600 32170
rect 56652 32118 56704 32170
rect 93264 32118 93316 32170
rect 93368 32118 93420 32170
rect 93472 32118 93524 32170
rect 130084 32118 130136 32170
rect 130188 32118 130240 32170
rect 130292 32118 130344 32170
rect 38034 31334 38086 31386
rect 38138 31334 38190 31386
rect 38242 31334 38294 31386
rect 74854 31334 74906 31386
rect 74958 31334 75010 31386
rect 75062 31334 75114 31386
rect 111674 31334 111726 31386
rect 111778 31334 111830 31386
rect 111882 31334 111934 31386
rect 148494 31334 148546 31386
rect 148598 31334 148650 31386
rect 148702 31334 148754 31386
rect 19624 30550 19676 30602
rect 19728 30550 19780 30602
rect 19832 30550 19884 30602
rect 56444 30550 56496 30602
rect 56548 30550 56600 30602
rect 56652 30550 56704 30602
rect 93264 30550 93316 30602
rect 93368 30550 93420 30602
rect 93472 30550 93524 30602
rect 130084 30550 130136 30602
rect 130188 30550 130240 30602
rect 130292 30550 130344 30602
rect 38034 29766 38086 29818
rect 38138 29766 38190 29818
rect 38242 29766 38294 29818
rect 74854 29766 74906 29818
rect 74958 29766 75010 29818
rect 75062 29766 75114 29818
rect 111674 29766 111726 29818
rect 111778 29766 111830 29818
rect 111882 29766 111934 29818
rect 148494 29766 148546 29818
rect 148598 29766 148650 29818
rect 148702 29766 148754 29818
rect 19624 28982 19676 29034
rect 19728 28982 19780 29034
rect 19832 28982 19884 29034
rect 56444 28982 56496 29034
rect 56548 28982 56600 29034
rect 56652 28982 56704 29034
rect 93264 28982 93316 29034
rect 93368 28982 93420 29034
rect 93472 28982 93524 29034
rect 130084 28982 130136 29034
rect 130188 28982 130240 29034
rect 130292 28982 130344 29034
rect 38034 28198 38086 28250
rect 38138 28198 38190 28250
rect 38242 28198 38294 28250
rect 74854 28198 74906 28250
rect 74958 28198 75010 28250
rect 75062 28198 75114 28250
rect 111674 28198 111726 28250
rect 111778 28198 111830 28250
rect 111882 28198 111934 28250
rect 148494 28198 148546 28250
rect 148598 28198 148650 28250
rect 148702 28198 148754 28250
rect 19624 27414 19676 27466
rect 19728 27414 19780 27466
rect 19832 27414 19884 27466
rect 56444 27414 56496 27466
rect 56548 27414 56600 27466
rect 56652 27414 56704 27466
rect 93264 27414 93316 27466
rect 93368 27414 93420 27466
rect 93472 27414 93524 27466
rect 130084 27414 130136 27466
rect 130188 27414 130240 27466
rect 130292 27414 130344 27466
rect 38034 26630 38086 26682
rect 38138 26630 38190 26682
rect 38242 26630 38294 26682
rect 74854 26630 74906 26682
rect 74958 26630 75010 26682
rect 75062 26630 75114 26682
rect 111674 26630 111726 26682
rect 111778 26630 111830 26682
rect 111882 26630 111934 26682
rect 148494 26630 148546 26682
rect 148598 26630 148650 26682
rect 148702 26630 148754 26682
rect 19624 25846 19676 25898
rect 19728 25846 19780 25898
rect 19832 25846 19884 25898
rect 56444 25846 56496 25898
rect 56548 25846 56600 25898
rect 56652 25846 56704 25898
rect 93264 25846 93316 25898
rect 93368 25846 93420 25898
rect 93472 25846 93524 25898
rect 130084 25846 130136 25898
rect 130188 25846 130240 25898
rect 130292 25846 130344 25898
rect 38034 25062 38086 25114
rect 38138 25062 38190 25114
rect 38242 25062 38294 25114
rect 74854 25062 74906 25114
rect 74958 25062 75010 25114
rect 75062 25062 75114 25114
rect 111674 25062 111726 25114
rect 111778 25062 111830 25114
rect 111882 25062 111934 25114
rect 148494 25062 148546 25114
rect 148598 25062 148650 25114
rect 148702 25062 148754 25114
rect 19624 24278 19676 24330
rect 19728 24278 19780 24330
rect 19832 24278 19884 24330
rect 56444 24278 56496 24330
rect 56548 24278 56600 24330
rect 56652 24278 56704 24330
rect 93264 24278 93316 24330
rect 93368 24278 93420 24330
rect 93472 24278 93524 24330
rect 130084 24278 130136 24330
rect 130188 24278 130240 24330
rect 130292 24278 130344 24330
rect 38034 23494 38086 23546
rect 38138 23494 38190 23546
rect 38242 23494 38294 23546
rect 74854 23494 74906 23546
rect 74958 23494 75010 23546
rect 75062 23494 75114 23546
rect 111674 23494 111726 23546
rect 111778 23494 111830 23546
rect 111882 23494 111934 23546
rect 148494 23494 148546 23546
rect 148598 23494 148650 23546
rect 148702 23494 148754 23546
rect 19624 22710 19676 22762
rect 19728 22710 19780 22762
rect 19832 22710 19884 22762
rect 56444 22710 56496 22762
rect 56548 22710 56600 22762
rect 56652 22710 56704 22762
rect 93264 22710 93316 22762
rect 93368 22710 93420 22762
rect 93472 22710 93524 22762
rect 130084 22710 130136 22762
rect 130188 22710 130240 22762
rect 130292 22710 130344 22762
rect 38034 21926 38086 21978
rect 38138 21926 38190 21978
rect 38242 21926 38294 21978
rect 74854 21926 74906 21978
rect 74958 21926 75010 21978
rect 75062 21926 75114 21978
rect 111674 21926 111726 21978
rect 111778 21926 111830 21978
rect 111882 21926 111934 21978
rect 148494 21926 148546 21978
rect 148598 21926 148650 21978
rect 148702 21926 148754 21978
rect 19624 21142 19676 21194
rect 19728 21142 19780 21194
rect 19832 21142 19884 21194
rect 56444 21142 56496 21194
rect 56548 21142 56600 21194
rect 56652 21142 56704 21194
rect 93264 21142 93316 21194
rect 93368 21142 93420 21194
rect 93472 21142 93524 21194
rect 130084 21142 130136 21194
rect 130188 21142 130240 21194
rect 130292 21142 130344 21194
rect 38034 20358 38086 20410
rect 38138 20358 38190 20410
rect 38242 20358 38294 20410
rect 74854 20358 74906 20410
rect 74958 20358 75010 20410
rect 75062 20358 75114 20410
rect 111674 20358 111726 20410
rect 111778 20358 111830 20410
rect 111882 20358 111934 20410
rect 148494 20358 148546 20410
rect 148598 20358 148650 20410
rect 148702 20358 148754 20410
rect 19624 19574 19676 19626
rect 19728 19574 19780 19626
rect 19832 19574 19884 19626
rect 56444 19574 56496 19626
rect 56548 19574 56600 19626
rect 56652 19574 56704 19626
rect 93264 19574 93316 19626
rect 93368 19574 93420 19626
rect 93472 19574 93524 19626
rect 130084 19574 130136 19626
rect 130188 19574 130240 19626
rect 130292 19574 130344 19626
rect 38034 18790 38086 18842
rect 38138 18790 38190 18842
rect 38242 18790 38294 18842
rect 74854 18790 74906 18842
rect 74958 18790 75010 18842
rect 75062 18790 75114 18842
rect 111674 18790 111726 18842
rect 111778 18790 111830 18842
rect 111882 18790 111934 18842
rect 148494 18790 148546 18842
rect 148598 18790 148650 18842
rect 148702 18790 148754 18842
rect 19624 18006 19676 18058
rect 19728 18006 19780 18058
rect 19832 18006 19884 18058
rect 56444 18006 56496 18058
rect 56548 18006 56600 18058
rect 56652 18006 56704 18058
rect 93264 18006 93316 18058
rect 93368 18006 93420 18058
rect 93472 18006 93524 18058
rect 130084 18006 130136 18058
rect 130188 18006 130240 18058
rect 130292 18006 130344 18058
rect 38034 17222 38086 17274
rect 38138 17222 38190 17274
rect 38242 17222 38294 17274
rect 74854 17222 74906 17274
rect 74958 17222 75010 17274
rect 75062 17222 75114 17274
rect 111674 17222 111726 17274
rect 111778 17222 111830 17274
rect 111882 17222 111934 17274
rect 148494 17222 148546 17274
rect 148598 17222 148650 17274
rect 148702 17222 148754 17274
rect 19624 16438 19676 16490
rect 19728 16438 19780 16490
rect 19832 16438 19884 16490
rect 56444 16438 56496 16490
rect 56548 16438 56600 16490
rect 56652 16438 56704 16490
rect 93264 16438 93316 16490
rect 93368 16438 93420 16490
rect 93472 16438 93524 16490
rect 130084 16438 130136 16490
rect 130188 16438 130240 16490
rect 130292 16438 130344 16490
rect 38034 15654 38086 15706
rect 38138 15654 38190 15706
rect 38242 15654 38294 15706
rect 74854 15654 74906 15706
rect 74958 15654 75010 15706
rect 75062 15654 75114 15706
rect 111674 15654 111726 15706
rect 111778 15654 111830 15706
rect 111882 15654 111934 15706
rect 148494 15654 148546 15706
rect 148598 15654 148650 15706
rect 148702 15654 148754 15706
rect 19624 14870 19676 14922
rect 19728 14870 19780 14922
rect 19832 14870 19884 14922
rect 56444 14870 56496 14922
rect 56548 14870 56600 14922
rect 56652 14870 56704 14922
rect 93264 14870 93316 14922
rect 93368 14870 93420 14922
rect 93472 14870 93524 14922
rect 130084 14870 130136 14922
rect 130188 14870 130240 14922
rect 130292 14870 130344 14922
rect 38034 14086 38086 14138
rect 38138 14086 38190 14138
rect 38242 14086 38294 14138
rect 74854 14086 74906 14138
rect 74958 14086 75010 14138
rect 75062 14086 75114 14138
rect 111674 14086 111726 14138
rect 111778 14086 111830 14138
rect 111882 14086 111934 14138
rect 148494 14086 148546 14138
rect 148598 14086 148650 14138
rect 148702 14086 148754 14138
rect 19624 13302 19676 13354
rect 19728 13302 19780 13354
rect 19832 13302 19884 13354
rect 56444 13302 56496 13354
rect 56548 13302 56600 13354
rect 56652 13302 56704 13354
rect 93264 13302 93316 13354
rect 93368 13302 93420 13354
rect 93472 13302 93524 13354
rect 130084 13302 130136 13354
rect 130188 13302 130240 13354
rect 130292 13302 130344 13354
rect 38034 12518 38086 12570
rect 38138 12518 38190 12570
rect 38242 12518 38294 12570
rect 74854 12518 74906 12570
rect 74958 12518 75010 12570
rect 75062 12518 75114 12570
rect 111674 12518 111726 12570
rect 111778 12518 111830 12570
rect 111882 12518 111934 12570
rect 148494 12518 148546 12570
rect 148598 12518 148650 12570
rect 148702 12518 148754 12570
rect 19624 11734 19676 11786
rect 19728 11734 19780 11786
rect 19832 11734 19884 11786
rect 56444 11734 56496 11786
rect 56548 11734 56600 11786
rect 56652 11734 56704 11786
rect 93264 11734 93316 11786
rect 93368 11734 93420 11786
rect 93472 11734 93524 11786
rect 130084 11734 130136 11786
rect 130188 11734 130240 11786
rect 130292 11734 130344 11786
rect 38034 10950 38086 11002
rect 38138 10950 38190 11002
rect 38242 10950 38294 11002
rect 74854 10950 74906 11002
rect 74958 10950 75010 11002
rect 75062 10950 75114 11002
rect 111674 10950 111726 11002
rect 111778 10950 111830 11002
rect 111882 10950 111934 11002
rect 148494 10950 148546 11002
rect 148598 10950 148650 11002
rect 148702 10950 148754 11002
rect 19624 10166 19676 10218
rect 19728 10166 19780 10218
rect 19832 10166 19884 10218
rect 56444 10166 56496 10218
rect 56548 10166 56600 10218
rect 56652 10166 56704 10218
rect 93264 10166 93316 10218
rect 93368 10166 93420 10218
rect 93472 10166 93524 10218
rect 130084 10166 130136 10218
rect 130188 10166 130240 10218
rect 130292 10166 130344 10218
rect 64990 9550 65042 9602
rect 38034 9382 38086 9434
rect 38138 9382 38190 9434
rect 38242 9382 38294 9434
rect 74854 9382 74906 9434
rect 74958 9382 75010 9434
rect 75062 9382 75114 9434
rect 111674 9382 111726 9434
rect 111778 9382 111830 9434
rect 111882 9382 111934 9434
rect 148494 9382 148546 9434
rect 148598 9382 148650 9434
rect 148702 9382 148754 9434
rect 64542 9102 64594 9154
rect 65774 9102 65826 9154
rect 124686 9102 124738 9154
rect 65438 8990 65490 9042
rect 124910 8990 124962 9042
rect 62190 8878 62242 8930
rect 63086 8878 63138 8930
rect 63534 8878 63586 8930
rect 66334 8878 66386 8930
rect 105198 8878 105250 8930
rect 123118 8878 123170 8930
rect 124126 8878 124178 8930
rect 125470 8878 125522 8930
rect 125918 8878 125970 8930
rect 64654 8766 64706 8818
rect 123790 8766 123842 8818
rect 19624 8598 19676 8650
rect 19728 8598 19780 8650
rect 19832 8598 19884 8650
rect 56444 8598 56496 8650
rect 56548 8598 56600 8650
rect 56652 8598 56704 8650
rect 93264 8598 93316 8650
rect 93368 8598 93420 8650
rect 93472 8598 93524 8650
rect 130084 8598 130136 8650
rect 130188 8598 130240 8650
rect 130292 8598 130344 8650
rect 64878 8430 64930 8482
rect 62638 8318 62690 8370
rect 121886 8318 121938 8370
rect 122782 8318 122834 8370
rect 124126 8318 124178 8370
rect 63870 8206 63922 8258
rect 64542 8206 64594 8258
rect 65998 8206 66050 8258
rect 67006 8206 67058 8258
rect 87950 8206 88002 8258
rect 89406 8206 89458 8258
rect 94782 8206 94834 8258
rect 95566 8206 95618 8258
rect 96126 8206 96178 8258
rect 104526 8206 104578 8258
rect 105758 8206 105810 8258
rect 107102 8206 107154 8258
rect 123566 8206 123618 8258
rect 125246 8206 125298 8258
rect 63982 8094 64034 8146
rect 65550 8094 65602 8146
rect 66558 8094 66610 8146
rect 88286 8094 88338 8146
rect 88510 8094 88562 8146
rect 89854 8094 89906 8146
rect 93774 8094 93826 8146
rect 95342 8094 95394 8146
rect 105982 8094 106034 8146
rect 106318 8094 106370 8146
rect 123454 8094 123506 8146
rect 28030 7982 28082 8034
rect 28590 7982 28642 8034
rect 60734 7982 60786 8034
rect 61630 7982 61682 8034
rect 62078 7982 62130 8034
rect 62750 7982 62802 8034
rect 86606 7982 86658 8034
rect 87054 7982 87106 8034
rect 87614 7982 87666 8034
rect 94446 7982 94498 8034
rect 96686 7982 96738 8034
rect 103966 7982 104018 8034
rect 104750 7982 104802 8034
rect 105422 7982 105474 8034
rect 122446 7982 122498 8034
rect 125022 7982 125074 8034
rect 125918 7982 125970 8034
rect 126254 7982 126306 8034
rect 126814 7982 126866 8034
rect 127262 7982 127314 8034
rect 38034 7814 38086 7866
rect 38138 7814 38190 7866
rect 38242 7814 38294 7866
rect 74854 7814 74906 7866
rect 74958 7814 75010 7866
rect 75062 7814 75114 7866
rect 111674 7814 111726 7866
rect 111778 7814 111830 7866
rect 111882 7814 111934 7866
rect 148494 7814 148546 7866
rect 148598 7814 148650 7866
rect 148702 7814 148754 7866
rect 67230 7646 67282 7698
rect 78430 7646 78482 7698
rect 85486 7646 85538 7698
rect 86046 7646 86098 7698
rect 89182 7646 89234 7698
rect 92542 7646 92594 7698
rect 93102 7646 93154 7698
rect 96014 7646 96066 7698
rect 107102 7646 107154 7698
rect 125806 7646 125858 7698
rect 126814 7646 126866 7698
rect 137118 7646 137170 7698
rect 139134 7646 139186 7698
rect 26910 7534 26962 7586
rect 27246 7534 27298 7586
rect 28814 7534 28866 7586
rect 29374 7534 29426 7586
rect 44270 7534 44322 7586
rect 59166 7534 59218 7586
rect 61854 7534 61906 7586
rect 62862 7534 62914 7586
rect 63534 7534 63586 7586
rect 65662 7534 65714 7586
rect 76302 7534 76354 7586
rect 76862 7534 76914 7586
rect 87838 7534 87890 7586
rect 88398 7534 88450 7586
rect 93662 7534 93714 7586
rect 94446 7534 94498 7586
rect 94894 7534 94946 7586
rect 104078 7534 104130 7586
rect 104414 7534 104466 7586
rect 105982 7534 106034 7586
rect 106318 7534 106370 7586
rect 116622 7534 116674 7586
rect 116958 7534 117010 7586
rect 121774 7534 121826 7586
rect 122110 7534 122162 7586
rect 26686 7422 26738 7474
rect 28590 7422 28642 7474
rect 30382 7422 30434 7474
rect 44606 7422 44658 7474
rect 59502 7422 59554 7474
rect 60958 7422 61010 7474
rect 61294 7422 61346 7474
rect 62078 7422 62130 7474
rect 63422 7422 63474 7474
rect 64206 7422 64258 7474
rect 65550 7422 65602 7474
rect 66334 7422 66386 7474
rect 77086 7422 77138 7474
rect 87614 7422 87666 7474
rect 95118 7422 95170 7474
rect 96462 7422 96514 7474
rect 105758 7422 105810 7474
rect 107550 7422 107602 7474
rect 116398 7422 116450 7474
rect 117742 7422 117794 7474
rect 122670 7422 122722 7474
rect 123342 7422 123394 7474
rect 137342 7422 137394 7474
rect 18398 7310 18450 7362
rect 19294 7310 19346 7362
rect 20302 7310 20354 7362
rect 29934 7310 29986 7362
rect 45166 7310 45218 7362
rect 47182 7310 47234 7362
rect 58158 7310 58210 7362
rect 58718 7310 58770 7362
rect 60286 7310 60338 7362
rect 75630 7310 75682 7362
rect 77982 7310 78034 7362
rect 86494 7310 86546 7362
rect 89630 7310 89682 7362
rect 103518 7310 103570 7362
rect 105422 7310 105474 7362
rect 115390 7310 115442 7362
rect 118190 7310 118242 7362
rect 121214 7310 121266 7362
rect 126926 7310 126978 7362
rect 127486 7310 127538 7362
rect 138126 7310 138178 7362
rect 138686 7310 138738 7362
rect 26350 7198 26402 7250
rect 28254 7198 28306 7250
rect 64542 7198 64594 7250
rect 66670 7198 66722 7250
rect 77422 7198 77474 7250
rect 87278 7198 87330 7250
rect 95454 7198 95506 7250
rect 116062 7198 116114 7250
rect 126366 7198 126418 7250
rect 127598 7198 127650 7250
rect 19624 7030 19676 7082
rect 19728 7030 19780 7082
rect 19832 7030 19884 7082
rect 56444 7030 56496 7082
rect 56548 7030 56600 7082
rect 56652 7030 56704 7082
rect 93264 7030 93316 7082
rect 93368 7030 93420 7082
rect 93472 7030 93524 7082
rect 130084 7030 130136 7082
rect 130188 7030 130240 7082
rect 130292 7030 130344 7082
rect 19630 6862 19682 6914
rect 43374 6862 43426 6914
rect 45950 6862 46002 6914
rect 124350 6862 124402 6914
rect 137454 6862 137506 6914
rect 28366 6750 28418 6802
rect 75630 6750 75682 6802
rect 78094 6750 78146 6802
rect 93998 6750 94050 6802
rect 139358 6750 139410 6802
rect 17614 6638 17666 6690
rect 18286 6638 18338 6690
rect 20526 6638 20578 6690
rect 26350 6638 26402 6690
rect 27134 6638 27186 6690
rect 44158 6638 44210 6690
rect 44830 6638 44882 6690
rect 45614 6638 45666 6690
rect 47966 6638 48018 6690
rect 53454 6638 53506 6690
rect 57150 6638 57202 6690
rect 57710 6638 57762 6690
rect 61966 6638 62018 6690
rect 62414 6638 62466 6690
rect 63086 6638 63138 6690
rect 66110 6638 66162 6690
rect 66670 6638 66722 6690
rect 67678 6638 67730 6690
rect 68126 6638 68178 6690
rect 69358 6638 69410 6690
rect 76414 6638 76466 6690
rect 77422 6638 77474 6690
rect 78542 6638 78594 6690
rect 86382 6638 86434 6690
rect 87054 6638 87106 6690
rect 87726 6638 87778 6690
rect 90750 6638 90802 6690
rect 94558 6638 94610 6690
rect 95454 6638 95506 6690
rect 95790 6638 95842 6690
rect 98926 6638 98978 6690
rect 105982 6638 106034 6690
rect 106654 6638 106706 6690
rect 115054 6638 115106 6690
rect 120654 6638 120706 6690
rect 121326 6638 121378 6690
rect 124910 6638 124962 6690
rect 125470 6638 125522 6690
rect 136782 6638 136834 6690
rect 140814 6638 140866 6690
rect 19070 6526 19122 6578
rect 19294 6526 19346 6578
rect 29598 6526 29650 6578
rect 42254 6526 42306 6578
rect 43038 6526 43090 6578
rect 44046 6526 44098 6578
rect 46174 6526 46226 6578
rect 46510 6526 46562 6578
rect 59950 6526 60002 6578
rect 61854 6526 61906 6578
rect 65326 6526 65378 6578
rect 72606 6526 72658 6578
rect 76302 6526 76354 6578
rect 107438 6526 107490 6578
rect 135662 6526 135714 6578
rect 135998 6526 136050 6578
rect 136670 6526 136722 6578
rect 137790 6526 137842 6578
rect 138686 6526 138738 6578
rect 139134 6526 139186 6578
rect 14590 6414 14642 6466
rect 15374 6414 15426 6466
rect 19966 6414 20018 6466
rect 26126 6414 26178 6466
rect 27358 6414 27410 6466
rect 27918 6414 27970 6466
rect 41918 6414 41970 6466
rect 47518 6414 47570 6466
rect 50542 6414 50594 6466
rect 50990 6414 51042 6466
rect 51326 6414 51378 6466
rect 52670 6414 52722 6466
rect 54014 6414 54066 6466
rect 60734 6414 60786 6466
rect 61294 6414 61346 6466
rect 66894 6414 66946 6466
rect 67566 6414 67618 6466
rect 68574 6414 68626 6466
rect 75294 6414 75346 6466
rect 77646 6414 77698 6466
rect 79102 6414 79154 6466
rect 86606 6414 86658 6466
rect 90190 6414 90242 6466
rect 94782 6414 94834 6466
rect 98254 6414 98306 6466
rect 102510 6414 102562 6466
rect 102958 6414 103010 6466
rect 103742 6414 103794 6466
rect 107102 6414 107154 6466
rect 109118 6414 109170 6466
rect 110798 6414 110850 6466
rect 114718 6414 114770 6466
rect 117294 6414 117346 6466
rect 120206 6414 120258 6466
rect 123790 6414 123842 6466
rect 128046 6414 128098 6466
rect 128606 6414 128658 6466
rect 129054 6414 129106 6466
rect 129390 6414 129442 6466
rect 139694 6414 139746 6466
rect 141262 6414 141314 6466
rect 38034 6246 38086 6298
rect 38138 6246 38190 6298
rect 38242 6246 38294 6298
rect 74854 6246 74906 6298
rect 74958 6246 75010 6298
rect 75062 6246 75114 6298
rect 111674 6246 111726 6298
rect 111778 6246 111830 6298
rect 111882 6246 111934 6298
rect 148494 6246 148546 6298
rect 148598 6246 148650 6298
rect 148702 6246 148754 6298
rect 16158 6078 16210 6130
rect 31390 6078 31442 6130
rect 38894 6078 38946 6130
rect 39454 6078 39506 6130
rect 39790 6078 39842 6130
rect 46734 6078 46786 6130
rect 53566 6078 53618 6130
rect 55134 6078 55186 6130
rect 62750 6078 62802 6130
rect 63982 6078 64034 6130
rect 65326 6078 65378 6130
rect 66110 6078 66162 6130
rect 87838 6078 87890 6130
rect 95342 6078 95394 6130
rect 95790 6078 95842 6130
rect 98254 6078 98306 6130
rect 104414 6078 104466 6130
rect 108222 6078 108274 6130
rect 109230 6078 109282 6130
rect 117854 6078 117906 6130
rect 118302 6078 118354 6130
rect 125582 6078 125634 6130
rect 126142 6078 126194 6130
rect 126590 6078 126642 6130
rect 127262 6078 127314 6130
rect 129390 6078 129442 6130
rect 134206 6078 134258 6130
rect 135774 6078 135826 6130
rect 138574 6078 138626 6130
rect 18734 5966 18786 6018
rect 19630 5966 19682 6018
rect 19966 5966 20018 6018
rect 30606 5966 30658 6018
rect 31726 5966 31778 6018
rect 53118 5966 53170 6018
rect 64318 5966 64370 6018
rect 75294 5966 75346 6018
rect 76526 5966 76578 6018
rect 79886 5966 79938 6018
rect 87502 5966 87554 6018
rect 109342 5966 109394 6018
rect 110238 5966 110290 6018
rect 115950 5966 116002 6018
rect 132974 5966 133026 6018
rect 137454 5966 137506 6018
rect 138014 5966 138066 6018
rect 140142 5966 140194 6018
rect 140702 5966 140754 6018
rect 141262 5966 141314 6018
rect 15934 5854 15986 5906
rect 17838 5854 17890 5906
rect 18174 5854 18226 5906
rect 18958 5854 19010 5906
rect 21534 5854 21586 5906
rect 27694 5854 27746 5906
rect 28254 5854 28306 5906
rect 43822 5854 43874 5906
rect 44270 5854 44322 5906
rect 47630 5854 47682 5906
rect 57822 5854 57874 5906
rect 59838 5854 59890 5906
rect 60510 5854 60562 5906
rect 68350 5854 68402 5906
rect 69022 5854 69074 5906
rect 75070 5854 75122 5906
rect 78766 5854 78818 5906
rect 79438 5854 79490 5906
rect 95118 5854 95170 5906
rect 105310 5854 105362 5906
rect 105758 5854 105810 5906
rect 111022 5854 111074 5906
rect 112366 5854 112418 5906
rect 113262 5854 113314 5906
rect 113710 5854 113762 5906
rect 117518 5854 117570 5906
rect 121998 5854 122050 5906
rect 122446 5854 122498 5906
rect 123118 5854 123170 5906
rect 129166 5854 129218 5906
rect 132414 5854 132466 5906
rect 133198 5854 133250 5906
rect 139582 5854 139634 5906
rect 9774 5742 9826 5794
rect 10110 5742 10162 5794
rect 11678 5742 11730 5794
rect 16942 5742 16994 5794
rect 20638 5742 20690 5794
rect 21198 5742 21250 5794
rect 55694 5742 55746 5794
rect 56366 5742 56418 5794
rect 56814 5742 56866 5794
rect 57486 5742 57538 5794
rect 58270 5742 58322 5794
rect 58830 5742 58882 5794
rect 59390 5742 59442 5794
rect 69358 5742 69410 5794
rect 79998 5742 80050 5794
rect 80446 5742 80498 5794
rect 81342 5742 81394 5794
rect 86830 5742 86882 5794
rect 89406 5742 89458 5794
rect 89966 5742 90018 5794
rect 96574 5742 96626 5794
rect 97246 5742 97298 5794
rect 98366 5742 98418 5794
rect 98926 5742 98978 5794
rect 102734 5742 102786 5794
rect 103182 5742 103234 5794
rect 103630 5742 103682 5794
rect 104302 5742 104354 5794
rect 109902 5742 109954 5794
rect 111582 5742 111634 5794
rect 121550 5742 121602 5794
rect 126702 5742 126754 5794
rect 127374 5742 127426 5794
rect 128046 5742 128098 5794
rect 129838 5742 129890 5794
rect 130286 5742 130338 5794
rect 133758 5742 133810 5794
rect 134654 5742 134706 5794
rect 136222 5742 136274 5794
rect 20526 5630 20578 5682
rect 47294 5630 47346 5682
rect 56366 5630 56418 5682
rect 56926 5630 56978 5682
rect 59278 5630 59330 5682
rect 63534 5630 63586 5682
rect 75742 5630 75794 5682
rect 89294 5630 89346 5682
rect 97358 5630 97410 5682
rect 103742 5630 103794 5682
rect 108782 5630 108834 5682
rect 116734 5630 116786 5682
rect 127934 5630 127986 5682
rect 132078 5630 132130 5682
rect 138238 5630 138290 5682
rect 19624 5462 19676 5514
rect 19728 5462 19780 5514
rect 19832 5462 19884 5514
rect 56444 5462 56496 5514
rect 56548 5462 56600 5514
rect 56652 5462 56704 5514
rect 93264 5462 93316 5514
rect 93368 5462 93420 5514
rect 93472 5462 93524 5514
rect 130084 5462 130136 5514
rect 130188 5462 130240 5514
rect 130292 5462 130344 5514
rect 20750 5294 20802 5346
rect 29710 5294 29762 5346
rect 47070 5294 47122 5346
rect 58830 5294 58882 5346
rect 67678 5294 67730 5346
rect 80894 5294 80946 5346
rect 90302 5294 90354 5346
rect 98030 5294 98082 5346
rect 103070 5294 103122 5346
rect 109566 5294 109618 5346
rect 115614 5294 115666 5346
rect 118526 5294 118578 5346
rect 130846 5294 130898 5346
rect 133422 5294 133474 5346
rect 137118 5294 137170 5346
rect 16718 5182 16770 5234
rect 28590 5182 28642 5234
rect 46398 5182 46450 5234
rect 47182 5182 47234 5234
rect 47630 5182 47682 5234
rect 52670 5182 52722 5234
rect 53678 5182 53730 5234
rect 63982 5182 64034 5234
rect 67790 5182 67842 5234
rect 68238 5182 68290 5234
rect 69694 5182 69746 5234
rect 75518 5182 75570 5234
rect 108222 5182 108274 5234
rect 109230 5182 109282 5234
rect 110910 5182 110962 5234
rect 111358 5182 111410 5234
rect 114942 5182 114994 5234
rect 115502 5182 115554 5234
rect 116286 5182 116338 5234
rect 116958 5182 117010 5234
rect 119534 5182 119586 5234
rect 124350 5182 124402 5234
rect 131854 5182 131906 5234
rect 132190 5182 132242 5234
rect 134766 5182 134818 5234
rect 135214 5182 135266 5234
rect 138462 5182 138514 5234
rect 139022 5182 139074 5234
rect 139470 5182 139522 5234
rect 139806 5182 139858 5234
rect 140814 5182 140866 5234
rect 7758 5070 7810 5122
rect 8206 5070 8258 5122
rect 10446 5070 10498 5122
rect 16158 5070 16210 5122
rect 17278 5070 17330 5122
rect 17726 5070 17778 5122
rect 21534 5070 21586 5122
rect 25118 5070 25170 5122
rect 25566 5070 25618 5122
rect 41022 5070 41074 5122
rect 41694 5070 41746 5122
rect 44718 5070 44770 5122
rect 45390 5070 45442 5122
rect 46510 5070 46562 5122
rect 52334 5070 52386 5122
rect 55358 5070 55410 5122
rect 55694 5070 55746 5122
rect 62862 5070 62914 5122
rect 67118 5070 67170 5122
rect 72606 5070 72658 5122
rect 77422 5070 77474 5122
rect 77758 5070 77810 5122
rect 86382 5070 86434 5122
rect 86718 5070 86770 5122
rect 89854 5070 89906 5122
rect 90414 5070 90466 5122
rect 93886 5070 93938 5122
rect 94558 5070 94610 5122
rect 94894 5070 94946 5122
rect 102622 5070 102674 5122
rect 106094 5070 106146 5122
rect 106766 5070 106818 5122
rect 110238 5070 110290 5122
rect 116174 5070 116226 5122
rect 120206 5070 120258 5122
rect 120878 5070 120930 5122
rect 121214 5070 121266 5122
rect 124910 5070 124962 5122
rect 128046 5070 128098 5122
rect 128382 5070 128434 5122
rect 129278 5070 129330 5122
rect 130958 5070 131010 5122
rect 133086 5070 133138 5122
rect 134206 5070 134258 5122
rect 137790 5070 137842 5122
rect 12126 4958 12178 5010
rect 29598 4958 29650 5010
rect 54350 4958 54402 5010
rect 54686 4958 54738 5010
rect 59278 4958 59330 5010
rect 60286 4958 60338 5010
rect 60622 4958 60674 5010
rect 85262 4958 85314 5010
rect 85598 4958 85650 5010
rect 107550 4958 107602 5010
rect 110126 4958 110178 5010
rect 117742 4958 117794 5010
rect 118302 4958 118354 5010
rect 129054 4958 129106 5010
rect 130286 4958 130338 5010
rect 133982 4958 134034 5010
rect 135774 4958 135826 5010
rect 136110 4958 136162 5010
rect 136782 4958 136834 5010
rect 137902 4958 137954 5010
rect 6190 4846 6242 4898
rect 11342 4846 11394 4898
rect 12238 4846 12290 4898
rect 12686 4846 12738 4898
rect 20078 4846 20130 4898
rect 22094 4846 22146 4898
rect 28030 4846 28082 4898
rect 30158 4846 30210 4898
rect 44158 4846 44210 4898
rect 58270 4846 58322 4898
rect 59614 4846 59666 4898
rect 69358 4846 69410 4898
rect 80110 4846 80162 4898
rect 84478 4846 84530 4898
rect 89294 4846 89346 4898
rect 90862 4846 90914 4898
rect 97358 4846 97410 4898
rect 103742 4846 103794 4898
rect 107214 4846 107266 4898
rect 108110 4846 108162 4898
rect 118862 4846 118914 4898
rect 123790 4846 123842 4898
rect 125694 4846 125746 4898
rect 129950 4846 130002 4898
rect 38034 4678 38086 4730
rect 38138 4678 38190 4730
rect 38242 4678 38294 4730
rect 74854 4678 74906 4730
rect 74958 4678 75010 4730
rect 75062 4678 75114 4730
rect 111674 4678 111726 4730
rect 111778 4678 111830 4730
rect 111882 4678 111934 4730
rect 148494 4678 148546 4730
rect 148598 4678 148650 4730
rect 148702 4678 148754 4730
rect 8206 4510 8258 4562
rect 12574 4510 12626 4562
rect 13358 4510 13410 4562
rect 13694 4510 13746 4562
rect 15710 4510 15762 4562
rect 16270 4510 16322 4562
rect 18174 4510 18226 4562
rect 21758 4510 21810 4562
rect 26462 4510 26514 4562
rect 28030 4510 28082 4562
rect 28702 4510 28754 4562
rect 29150 4510 29202 4562
rect 46734 4510 46786 4562
rect 48190 4510 48242 4562
rect 54126 4510 54178 4562
rect 57934 4510 57986 4562
rect 58830 4510 58882 4562
rect 65326 4510 65378 4562
rect 66110 4510 66162 4562
rect 69806 4510 69858 4562
rect 70254 4510 70306 4562
rect 79998 4510 80050 4562
rect 85934 4510 85986 4562
rect 86382 4510 86434 4562
rect 88510 4510 88562 4562
rect 89630 4510 89682 4562
rect 90078 4510 90130 4562
rect 103966 4510 104018 4562
rect 104414 4510 104466 4562
rect 108110 4510 108162 4562
rect 110910 4510 110962 4562
rect 114830 4510 114882 4562
rect 115614 4510 115666 4562
rect 118974 4510 119026 4562
rect 121326 4510 121378 4562
rect 125806 4510 125858 4562
rect 128046 4510 128098 4562
rect 131966 4510 132018 4562
rect 133646 4510 133698 4562
rect 137118 4510 137170 4562
rect 138350 4510 138402 4562
rect 138798 4510 138850 4562
rect 142046 4510 142098 4562
rect 145742 4510 145794 4562
rect 7758 4398 7810 4450
rect 16830 4398 16882 4450
rect 27134 4398 27186 4450
rect 27470 4398 27522 4450
rect 28142 4398 28194 4450
rect 29598 4398 29650 4450
rect 54686 4398 54738 4450
rect 55246 4398 55298 4450
rect 56366 4398 56418 4450
rect 58494 4398 58546 4450
rect 61294 4398 61346 4450
rect 78430 4398 78482 4450
rect 79886 4398 79938 4450
rect 80446 4398 80498 4450
rect 89294 4398 89346 4450
rect 111358 4398 111410 4450
rect 119310 4398 119362 4450
rect 127486 4398 127538 4450
rect 128158 4398 128210 4450
rect 137454 4398 137506 4450
rect 5854 4286 5906 4338
rect 6974 4286 7026 4338
rect 7534 4286 7586 4338
rect 8318 4286 8370 4338
rect 8542 4286 8594 4338
rect 8766 4286 8818 4338
rect 8990 4286 9042 4338
rect 9886 4286 9938 4338
rect 10222 4286 10274 4338
rect 15374 4286 15426 4338
rect 17614 4286 17666 4338
rect 20638 4286 20690 4338
rect 21310 4286 21362 4338
rect 22094 4286 22146 4338
rect 22542 4286 22594 4338
rect 26126 4286 26178 4338
rect 52894 4286 52946 4338
rect 53454 4286 53506 4338
rect 54462 4286 54514 4338
rect 56702 4286 56754 4338
rect 57598 4286 57650 4338
rect 63870 4286 63922 4338
rect 68350 4286 68402 4338
rect 68910 4286 68962 4338
rect 69470 4286 69522 4338
rect 70702 4286 70754 4338
rect 72606 4286 72658 4338
rect 74846 4286 74898 4338
rect 79102 4286 79154 4338
rect 105310 4286 105362 4338
rect 105758 4286 105810 4338
rect 110462 4286 110514 4338
rect 114382 4286 114434 4338
rect 117966 4286 118018 4338
rect 118526 4286 118578 4338
rect 122222 4286 122274 4338
rect 122894 4286 122946 4338
rect 123342 4286 123394 4338
rect 127262 4286 127314 4338
rect 128942 4286 128994 4338
rect 129502 4286 129554 4338
rect 133870 4286 133922 4338
rect 138014 4286 138066 4338
rect 141710 4286 141762 4338
rect 145966 4286 146018 4338
rect 4846 4174 4898 4226
rect 6526 4174 6578 4226
rect 14478 4174 14530 4226
rect 14926 4174 14978 4226
rect 16942 4174 16994 4226
rect 25006 4174 25058 4226
rect 25678 4174 25730 4226
rect 31726 4174 31778 4226
rect 32958 4174 33010 4226
rect 33966 4174 34018 4226
rect 36878 4174 36930 4226
rect 37214 4174 37266 4226
rect 38670 4174 38722 4226
rect 40798 4174 40850 4226
rect 42590 4174 42642 4226
rect 44718 4174 44770 4226
rect 45054 4174 45106 4226
rect 47182 4174 47234 4226
rect 48750 4174 48802 4226
rect 51886 4174 51938 4226
rect 55918 4174 55970 4226
rect 81790 4174 81842 4226
rect 93550 4174 93602 4226
rect 97582 4174 97634 4226
rect 101614 4174 101666 4226
rect 109454 4174 109506 4226
rect 113710 4174 113762 4226
rect 121774 4174 121826 4226
rect 126366 4174 126418 4226
rect 132974 4174 133026 4226
rect 134430 4174 134482 4226
rect 141262 4174 141314 4226
rect 145294 4174 145346 4226
rect 108782 4062 108834 4114
rect 132638 4062 132690 4114
rect 19624 3894 19676 3946
rect 19728 3894 19780 3946
rect 19832 3894 19884 3946
rect 56444 3894 56496 3946
rect 56548 3894 56600 3946
rect 56652 3894 56704 3946
rect 93264 3894 93316 3946
rect 93368 3894 93420 3946
rect 93472 3894 93524 3946
rect 130084 3894 130136 3946
rect 130188 3894 130240 3946
rect 130292 3894 130344 3946
rect 8094 3726 8146 3778
rect 12238 3726 12290 3778
rect 17614 3726 17666 3778
rect 17950 3726 18002 3778
rect 18734 3726 18786 3778
rect 54798 3726 54850 3778
rect 55134 3726 55186 3778
rect 108110 3726 108162 3778
rect 108446 3726 108498 3778
rect 127262 3726 127314 3778
rect 12350 3614 12402 3666
rect 12910 3614 12962 3666
rect 19630 3614 19682 3666
rect 21534 3614 21586 3666
rect 35310 3614 35362 3666
rect 43374 3614 43426 3666
rect 47406 3614 47458 3666
rect 75630 3614 75682 3666
rect 78990 3614 79042 3666
rect 94670 3614 94722 3666
rect 102734 3614 102786 3666
rect 110686 3614 110738 3666
rect 112366 3614 112418 3666
rect 115726 3614 115778 3666
rect 119310 3614 119362 3666
rect 123342 3614 123394 3666
rect 123790 3614 123842 3666
rect 127374 3614 127426 3666
rect 131630 3614 131682 3666
rect 135886 3614 135938 3666
rect 138014 3614 138066 3666
rect 139918 3614 139970 3666
rect 143950 3614 144002 3666
rect 5854 3502 5906 3554
rect 7310 3502 7362 3554
rect 8542 3502 8594 3554
rect 8654 3502 8706 3554
rect 8766 3502 8818 3554
rect 15262 3502 15314 3554
rect 16494 3502 16546 3554
rect 17614 3502 17666 3554
rect 20638 3502 20690 3554
rect 22318 3502 22370 3554
rect 26574 3502 26626 3554
rect 31390 3502 31442 3554
rect 36318 3502 36370 3554
rect 40238 3502 40290 3554
rect 41246 3502 41298 3554
rect 42254 3502 42306 3554
rect 44158 3502 44210 3554
rect 46174 3502 46226 3554
rect 48078 3502 48130 3554
rect 51998 3502 52050 3554
rect 55918 3502 55970 3554
rect 57934 3502 57986 3554
rect 58942 3502 58994 3554
rect 59838 3502 59890 3554
rect 61630 3502 61682 3554
rect 62414 3502 62466 3554
rect 63646 3502 63698 3554
rect 65550 3502 65602 3554
rect 66558 3502 66610 3554
rect 67566 3502 67618 3554
rect 69694 3502 69746 3554
rect 70254 3502 70306 3554
rect 70590 3502 70642 3554
rect 71710 3502 71762 3554
rect 73614 3502 73666 3554
rect 77534 3502 77586 3554
rect 81454 3502 81506 3554
rect 82910 3502 82962 3554
rect 85374 3502 85426 3554
rect 89294 3502 89346 3554
rect 93214 3502 93266 3554
rect 97246 3502 97298 3554
rect 98702 3502 98754 3554
rect 101278 3502 101330 3554
rect 105310 3502 105362 3554
rect 109230 3502 109282 3554
rect 113374 3502 113426 3554
rect 117182 3502 117234 3554
rect 118302 3502 118354 3554
rect 121438 3502 121490 3554
rect 125246 3502 125298 3554
rect 126142 3502 126194 3554
rect 129502 3502 129554 3554
rect 131070 3502 131122 3554
rect 133310 3502 133362 3554
rect 137566 3502 137618 3554
rect 140366 3502 140418 3554
rect 144398 3502 144450 3554
rect 6302 3390 6354 3442
rect 9998 3390 10050 3442
rect 10334 3390 10386 3442
rect 10894 3390 10946 3442
rect 11678 3390 11730 3442
rect 14366 3390 14418 3442
rect 15934 3390 15986 3442
rect 18846 3390 18898 3442
rect 22990 3390 23042 3442
rect 23438 3390 23490 3442
rect 25678 3390 25730 3442
rect 27470 3390 27522 3442
rect 28590 3390 28642 3442
rect 29598 3390 29650 3442
rect 30494 3390 30546 3442
rect 31950 3390 32002 3442
rect 33182 3390 33234 3442
rect 34190 3390 34242 3442
rect 37102 3390 37154 3442
rect 38446 3390 38498 3442
rect 39342 3390 39394 3442
rect 44942 3390 44994 3442
rect 48974 3390 49026 3442
rect 49870 3390 49922 3442
rect 50318 3390 50370 3442
rect 51214 3390 51266 3442
rect 53342 3390 53394 3442
rect 54014 3390 54066 3442
rect 54574 3390 54626 3442
rect 57038 3390 57090 3442
rect 60958 3390 61010 3442
rect 62750 3390 62802 3442
rect 63310 3390 63362 3442
rect 64878 3390 64930 3442
rect 68798 3390 68850 3442
rect 72718 3390 72770 3442
rect 74510 3390 74562 3442
rect 74958 3390 75010 3442
rect 76638 3390 76690 3442
rect 78430 3390 78482 3442
rect 79326 3390 79378 3442
rect 80558 3390 80610 3442
rect 82014 3390 82066 3442
rect 82350 3390 82402 3442
rect 84478 3390 84530 3442
rect 86270 3390 86322 3442
rect 86718 3390 86770 3442
rect 88398 3390 88450 3442
rect 90190 3390 90242 3442
rect 90638 3390 90690 3442
rect 92318 3390 92370 3442
rect 93774 3390 93826 3442
rect 96350 3390 96402 3442
rect 97806 3390 97858 3442
rect 100382 3390 100434 3442
rect 101838 3390 101890 3442
rect 104414 3390 104466 3442
rect 106206 3390 106258 3442
rect 106654 3390 106706 3442
rect 109006 3390 109058 3442
rect 109902 3390 109954 3442
rect 111470 3390 111522 3442
rect 113934 3390 113986 3442
rect 116510 3390 116562 3442
rect 120542 3390 120594 3442
rect 121998 3390 122050 3442
rect 124574 3390 124626 3442
rect 128606 3390 128658 3442
rect 130062 3390 130114 3442
rect 132638 3390 132690 3442
rect 136670 3390 136722 3442
rect 141262 3390 141314 3442
rect 145294 3390 145346 3442
rect 6638 3278 6690 3330
rect 7534 3278 7586 3330
rect 11342 3278 11394 3330
rect 16718 3278 16770 3330
rect 22094 3278 22146 3330
rect 23774 3278 23826 3330
rect 27806 3278 27858 3330
rect 29262 3278 29314 3330
rect 32286 3278 32338 3330
rect 33518 3278 33570 3330
rect 34526 3278 34578 3330
rect 37438 3278 37490 3330
rect 38110 3278 38162 3330
rect 41022 3278 41074 3330
rect 42030 3278 42082 3330
rect 45278 3278 45330 3330
rect 45950 3278 46002 3330
rect 49310 3278 49362 3330
rect 50654 3278 50706 3330
rect 51662 3278 51714 3330
rect 53006 3278 53058 3330
rect 58606 3278 58658 3330
rect 59502 3278 59554 3330
rect 66334 3278 66386 3330
rect 67230 3278 67282 3330
rect 74174 3278 74226 3330
rect 78094 3278 78146 3330
rect 85934 3278 85986 3330
rect 89854 3278 89906 3330
rect 94110 3278 94162 3330
rect 98142 3278 98194 3330
rect 102174 3278 102226 3330
rect 105870 3278 105922 3330
rect 110238 3278 110290 3330
rect 114270 3278 114322 3330
rect 117966 3278 118018 3330
rect 122334 3278 122386 3330
rect 126366 3278 126418 3330
rect 130398 3278 130450 3330
rect 38034 3110 38086 3162
rect 38138 3110 38190 3162
rect 38242 3110 38294 3162
rect 74854 3110 74906 3162
rect 74958 3110 75010 3162
rect 75062 3110 75114 3162
rect 111674 3110 111726 3162
rect 111778 3110 111830 3162
rect 111882 3110 111934 3162
rect 148494 3110 148546 3162
rect 148598 3110 148650 3162
rect 148702 3110 148754 3162
rect 105870 2942 105922 2994
rect 106878 2942 106930 2994
<< metal2 >>
rect 4592 39200 4704 40000
rect 5488 39200 5600 40000
rect 6384 39200 6496 40000
rect 7280 39200 7392 40000
rect 7644 39228 8036 39284
rect 4620 36372 4676 39200
rect 5516 37828 5572 39200
rect 5516 37772 6020 37828
rect 5964 36594 6020 37772
rect 5964 36542 5966 36594
rect 6018 36542 6020 36594
rect 5964 36530 6020 36542
rect 4844 36372 4900 36382
rect 4620 36370 4900 36372
rect 4620 36318 4846 36370
rect 4898 36318 4900 36370
rect 4620 36316 4900 36318
rect 4844 36306 4900 36316
rect 6076 35924 6132 35934
rect 6076 35830 6132 35868
rect 6412 35812 6468 39200
rect 7308 39060 7364 39200
rect 7644 39060 7700 39228
rect 7308 39004 7700 39060
rect 7980 36596 8036 39228
rect 8176 39200 8288 40000
rect 9072 39200 9184 40000
rect 9968 39200 10080 40000
rect 10864 39200 10976 40000
rect 11760 39200 11872 40000
rect 12656 39200 12768 40000
rect 13552 39200 13664 40000
rect 13804 39228 14308 39284
rect 8204 36820 8260 39200
rect 8876 37156 8932 37166
rect 8204 36764 8372 36820
rect 8204 36596 8260 36606
rect 7980 36594 8260 36596
rect 7980 36542 8206 36594
rect 8258 36542 8260 36594
rect 7980 36540 8260 36542
rect 8204 36530 8260 36540
rect 6972 36482 7028 36494
rect 6972 36430 6974 36482
rect 7026 36430 7028 36482
rect 6972 35924 7028 36430
rect 6972 35858 7028 35868
rect 7644 36482 7700 36494
rect 7644 36430 7646 36482
rect 7698 36430 7700 36482
rect 6412 35746 6468 35756
rect 7532 35812 7588 35822
rect 7532 35718 7588 35756
rect 6636 35698 6692 35710
rect 6636 35646 6638 35698
rect 6690 35646 6692 35698
rect 6188 34916 6244 34926
rect 6188 34822 6244 34860
rect 6636 34802 6692 35646
rect 6972 34916 7028 34926
rect 6972 34822 7028 34860
rect 6636 34750 6638 34802
rect 6690 34750 6692 34802
rect 6636 34738 6692 34750
rect 7532 34804 7588 34814
rect 7644 34804 7700 36430
rect 7532 34802 7700 34804
rect 7532 34750 7534 34802
rect 7586 34750 7700 34802
rect 7532 34748 7700 34750
rect 7868 35140 7924 35150
rect 7868 34914 7924 35084
rect 7868 34862 7870 34914
rect 7922 34862 7924 34914
rect 7532 34738 7588 34748
rect 7532 34356 7588 34366
rect 7868 34356 7924 34862
rect 7532 34354 7924 34356
rect 7532 34302 7534 34354
rect 7586 34302 7924 34354
rect 7532 34300 7924 34302
rect 7532 34290 7588 34300
rect 7868 7588 7924 34300
rect 7980 34356 8036 34366
rect 8316 34356 8372 36764
rect 8764 35698 8820 35710
rect 8764 35646 8766 35698
rect 8818 35646 8820 35698
rect 8764 35588 8820 35646
rect 8764 35522 8820 35532
rect 8876 35140 8932 37100
rect 8988 36484 9044 36494
rect 8988 35922 9044 36428
rect 8988 35870 8990 35922
rect 9042 35870 9044 35922
rect 8988 35858 9044 35870
rect 8876 35074 8932 35084
rect 9100 35140 9156 39200
rect 9996 36932 10052 39200
rect 9996 36876 10500 36932
rect 10444 36594 10500 36876
rect 10444 36542 10446 36594
rect 10498 36542 10500 36594
rect 10444 36530 10500 36542
rect 9772 36484 9828 36494
rect 9772 36390 9828 36428
rect 10892 36036 10948 39200
rect 11788 36260 11844 39200
rect 12684 37828 12740 39200
rect 13580 39060 13636 39200
rect 13804 39060 13860 39228
rect 13580 39004 13860 39060
rect 12124 37772 12740 37828
rect 12124 36594 12180 37772
rect 12124 36542 12126 36594
rect 12178 36542 12180 36594
rect 12124 36530 12180 36542
rect 14252 36596 14308 39228
rect 14448 39200 14560 40000
rect 15344 39200 15456 40000
rect 16240 39200 16352 40000
rect 17136 39200 17248 40000
rect 18032 39200 18144 40000
rect 18928 39200 19040 40000
rect 19824 39200 19936 40000
rect 20720 39200 20832 40000
rect 21084 39228 21476 39284
rect 14252 36540 14420 36596
rect 12572 36482 12628 36494
rect 12572 36430 12574 36482
rect 12626 36430 12628 36482
rect 11788 36204 11956 36260
rect 10892 35970 10948 35980
rect 11788 36036 11844 36046
rect 10556 35810 10612 35822
rect 10556 35758 10558 35810
rect 10610 35758 10612 35810
rect 10332 35698 10388 35710
rect 10332 35646 10334 35698
rect 10386 35646 10388 35698
rect 9660 35588 9716 35598
rect 9660 35494 9716 35532
rect 9100 35074 9156 35084
rect 10108 35140 10164 35150
rect 10108 35026 10164 35084
rect 10108 34974 10110 35026
rect 10162 34974 10164 35026
rect 10108 34962 10164 34974
rect 10332 35028 10388 35646
rect 10556 35700 10612 35758
rect 11116 35700 11172 35710
rect 10556 35698 11172 35700
rect 10556 35646 11118 35698
rect 11170 35646 11172 35698
rect 10556 35644 11172 35646
rect 11116 35634 11172 35644
rect 11788 35586 11844 35980
rect 11788 35534 11790 35586
rect 11842 35534 11844 35586
rect 11788 35522 11844 35534
rect 10332 34962 10388 34972
rect 11004 35028 11060 35038
rect 8540 34914 8596 34926
rect 9324 34916 9380 34926
rect 8540 34862 8542 34914
rect 8594 34862 8596 34914
rect 8540 34468 8596 34862
rect 8764 34914 9380 34916
rect 8764 34862 9326 34914
rect 9378 34862 9380 34914
rect 8764 34860 9380 34862
rect 8764 34802 8820 34860
rect 9324 34850 9380 34860
rect 8764 34750 8766 34802
rect 8818 34750 8820 34802
rect 8764 34738 8820 34750
rect 8540 34402 8596 34412
rect 8876 34468 8932 34478
rect 7980 34354 8484 34356
rect 7980 34302 7982 34354
rect 8034 34302 8484 34354
rect 7980 34300 8484 34302
rect 7980 34290 8036 34300
rect 8428 34242 8484 34300
rect 8428 34190 8430 34242
rect 8482 34190 8484 34242
rect 8428 34178 8484 34190
rect 8764 34244 8820 34254
rect 8764 34150 8820 34188
rect 7868 7522 7924 7532
rect 8876 5236 8932 34412
rect 9660 34468 9716 34478
rect 9660 34354 9716 34412
rect 9660 34302 9662 34354
rect 9714 34302 9716 34354
rect 9660 34290 9716 34302
rect 11004 34356 11060 34972
rect 11788 34916 11844 34926
rect 11900 34916 11956 36204
rect 11788 34914 11956 34916
rect 11788 34862 11790 34914
rect 11842 34862 11956 34914
rect 11788 34860 11956 34862
rect 11788 34850 11844 34860
rect 11004 34290 11060 34300
rect 11116 34804 11172 34814
rect 11116 20188 11172 34748
rect 11900 34356 11956 34860
rect 12012 35700 12068 35710
rect 12012 34802 12068 35644
rect 12012 34750 12014 34802
rect 12066 34750 12068 34802
rect 12012 34738 12068 34750
rect 12572 34802 12628 36430
rect 13916 36484 13972 36494
rect 13916 36482 14308 36484
rect 13916 36430 13918 36482
rect 13970 36430 14308 36482
rect 13916 36428 14308 36430
rect 13916 36418 13972 36428
rect 13244 35812 13300 35822
rect 13244 35718 13300 35756
rect 13804 35812 13860 35822
rect 13020 35698 13076 35710
rect 13020 35646 13022 35698
rect 13074 35646 13076 35698
rect 12908 34916 12964 34926
rect 12908 34822 12964 34860
rect 12572 34750 12574 34802
rect 12626 34750 12628 34802
rect 12572 34738 12628 34750
rect 12236 34356 12292 34366
rect 11900 34354 12292 34356
rect 11900 34302 12238 34354
rect 12290 34302 12292 34354
rect 11900 34300 12292 34302
rect 12236 34290 12292 34300
rect 13020 34020 13076 35646
rect 13804 35698 13860 35756
rect 13804 35646 13806 35698
rect 13858 35646 13860 35698
rect 13804 35634 13860 35646
rect 13580 34916 13636 34926
rect 13580 34822 13636 34860
rect 14252 34802 14308 36428
rect 14364 35588 14420 36540
rect 14476 36594 14532 39200
rect 14476 36542 14478 36594
rect 14530 36542 14532 36594
rect 14476 36530 14532 36542
rect 14476 35588 14532 35598
rect 14364 35586 14532 35588
rect 14364 35534 14478 35586
rect 14530 35534 14532 35586
rect 14364 35532 14532 35534
rect 14476 35522 14532 35532
rect 14252 34750 14254 34802
rect 14306 34750 14308 34802
rect 14252 34738 14308 34750
rect 14588 34916 14644 34926
rect 13020 33954 13076 33964
rect 13468 34020 13524 34030
rect 13468 33926 13524 33964
rect 14252 31108 14308 31118
rect 11116 20132 11284 20188
rect 8876 5170 8932 5180
rect 9772 5794 9828 5806
rect 9772 5742 9774 5794
rect 9826 5742 9828 5794
rect 7756 5124 7812 5134
rect 7756 5030 7812 5068
rect 8204 5122 8260 5134
rect 8204 5070 8206 5122
rect 8258 5070 8260 5122
rect 6188 4898 6244 4910
rect 6188 4846 6190 4898
rect 6242 4846 6244 4898
rect 5852 4788 5908 4798
rect 5852 4338 5908 4732
rect 6188 4788 6244 4846
rect 6188 4722 6244 4732
rect 8204 4562 8260 5070
rect 8204 4510 8206 4562
rect 8258 4510 8260 4562
rect 8204 4498 8260 4510
rect 7756 4452 7812 4462
rect 7756 4358 7812 4396
rect 5852 4286 5854 4338
rect 5906 4286 5908 4338
rect 5852 4274 5908 4286
rect 6972 4340 7028 4350
rect 6972 4246 7028 4284
rect 7532 4340 7588 4350
rect 7532 4338 7700 4340
rect 7532 4286 7534 4338
rect 7586 4286 7700 4338
rect 7532 4284 7700 4286
rect 7532 4274 7588 4284
rect 4844 4228 4900 4238
rect 4396 4226 4900 4228
rect 4396 4174 4846 4226
rect 4898 4174 4900 4226
rect 4396 4172 4900 4174
rect 4396 800 4452 4172
rect 4844 4162 4900 4172
rect 6524 4226 6580 4238
rect 6524 4174 6526 4226
rect 6578 4174 6580 4226
rect 5852 3556 5908 3566
rect 5852 3462 5908 3500
rect 6300 3444 6356 3454
rect 6300 3350 6356 3388
rect 6524 3444 6580 4174
rect 7644 3892 7700 4284
rect 8316 4338 8372 4350
rect 8316 4286 8318 4338
rect 8370 4286 8372 4338
rect 7644 3836 8148 3892
rect 8092 3778 8148 3836
rect 8092 3726 8094 3778
rect 8146 3726 8148 3778
rect 8092 3714 8148 3726
rect 8316 3668 8372 4286
rect 8540 4340 8596 4350
rect 8764 4340 8820 4350
rect 8988 4340 9044 4350
rect 8540 4338 8708 4340
rect 8540 4286 8542 4338
rect 8594 4286 8708 4338
rect 8540 4284 8708 4286
rect 8540 4274 8596 4284
rect 8316 3602 8372 3612
rect 8540 3892 8596 3902
rect 7308 3556 7364 3566
rect 7308 3462 7364 3500
rect 8428 3556 8484 3566
rect 6524 3378 6580 3388
rect 7084 3444 7140 3454
rect 6636 3332 6692 3342
rect 6636 3238 6692 3276
rect 5740 924 6020 980
rect 5740 800 5796 924
rect 4368 0 4480 800
rect 5712 0 5824 800
rect 5964 196 6020 924
rect 7084 800 7140 3388
rect 7532 3330 7588 3342
rect 7532 3278 7534 3330
rect 7586 3278 7588 3330
rect 7532 2996 7588 3278
rect 7532 2930 7588 2940
rect 8428 800 8484 3500
rect 8540 3554 8596 3836
rect 8540 3502 8542 3554
rect 8594 3502 8596 3554
rect 8540 3490 8596 3502
rect 8652 3554 8708 4284
rect 8764 4338 8932 4340
rect 8764 4286 8766 4338
rect 8818 4286 8932 4338
rect 8764 4284 8932 4286
rect 8764 4274 8820 4284
rect 8652 3502 8654 3554
rect 8706 3502 8708 3554
rect 8652 3332 8708 3502
rect 8764 3668 8820 3678
rect 8764 3554 8820 3612
rect 8764 3502 8766 3554
rect 8818 3502 8820 3554
rect 8764 3490 8820 3502
rect 8652 3266 8708 3276
rect 8876 3332 8932 4284
rect 8988 3892 9044 4284
rect 8988 3826 9044 3836
rect 9772 3892 9828 5742
rect 10108 5794 10164 5806
rect 10108 5742 10110 5794
rect 10162 5742 10164 5794
rect 9884 5124 9940 5134
rect 9884 4338 9940 5068
rect 9884 4286 9886 4338
rect 9938 4286 9940 4338
rect 9884 4274 9940 4286
rect 9772 3826 9828 3836
rect 9996 3668 10052 3678
rect 8876 3266 8932 3276
rect 9772 3444 9828 3454
rect 9772 800 9828 3388
rect 9996 3442 10052 3612
rect 9996 3390 9998 3442
rect 10050 3390 10052 3442
rect 9996 3378 10052 3390
rect 10108 3444 10164 5742
rect 10444 5122 10500 5134
rect 10444 5070 10446 5122
rect 10498 5070 10500 5122
rect 10220 4452 10276 4462
rect 10220 4338 10276 4396
rect 10220 4286 10222 4338
rect 10274 4286 10276 4338
rect 10220 4274 10276 4286
rect 10444 3780 10500 5070
rect 10444 3714 10500 3724
rect 10108 3378 10164 3388
rect 10332 3444 10388 3454
rect 10332 3350 10388 3388
rect 10892 3444 10948 3454
rect 11116 3444 11172 3454
rect 10892 3442 11116 3444
rect 10892 3390 10894 3442
rect 10946 3390 11116 3442
rect 10892 3388 11116 3390
rect 10892 3378 10948 3388
rect 11116 800 11172 3388
rect 11228 3220 11284 20132
rect 11676 5794 11732 5806
rect 11676 5742 11678 5794
rect 11730 5742 11732 5794
rect 11676 5124 11732 5742
rect 11676 5058 11732 5068
rect 12124 5012 12180 5022
rect 12124 4918 12180 4956
rect 12684 5012 12740 5022
rect 11340 4900 11396 4910
rect 11340 4806 11396 4844
rect 12236 4900 12292 4910
rect 12236 4898 12628 4900
rect 12236 4846 12238 4898
rect 12290 4846 12628 4898
rect 12236 4844 12628 4846
rect 12236 4834 12292 4844
rect 12572 4562 12628 4844
rect 12572 4510 12574 4562
rect 12626 4510 12628 4562
rect 12572 4498 12628 4510
rect 12684 4898 12740 4956
rect 12684 4846 12686 4898
rect 12738 4846 12740 4898
rect 12348 4452 12404 4462
rect 12236 3780 12292 3790
rect 12236 3686 12292 3724
rect 12348 3666 12404 4396
rect 12684 4452 12740 4846
rect 13692 5012 13748 5022
rect 13356 4788 13412 4798
rect 13356 4562 13412 4732
rect 13356 4510 13358 4562
rect 13410 4510 13412 4562
rect 13356 4498 13412 4510
rect 13692 4562 13748 4956
rect 14252 4900 14308 31052
rect 14588 9268 14644 34860
rect 14812 34916 14868 34926
rect 14812 34354 14868 34860
rect 15260 34916 15316 34926
rect 15372 34916 15428 39200
rect 15820 37380 15876 37390
rect 15820 34916 15876 37324
rect 16044 36596 16100 36606
rect 16044 36502 16100 36540
rect 15260 34914 15764 34916
rect 15260 34862 15262 34914
rect 15314 34862 15764 34914
rect 15260 34860 15764 34862
rect 15260 34850 15316 34860
rect 15484 34692 15540 34702
rect 15484 34598 15540 34636
rect 14812 34302 14814 34354
rect 14866 34302 14868 34354
rect 14812 34290 14868 34302
rect 15708 34354 15764 34860
rect 15820 34850 15876 34860
rect 15932 35698 15988 35710
rect 15932 35646 15934 35698
rect 15986 35646 15988 35698
rect 15932 34804 15988 35646
rect 16268 35588 16324 39200
rect 17164 36596 17220 39200
rect 18060 37044 18116 39200
rect 18060 36988 18452 37044
rect 17164 36530 17220 36540
rect 16716 36484 16772 36494
rect 16716 36482 16996 36484
rect 16716 36430 16718 36482
rect 16770 36430 16996 36482
rect 16716 36428 16996 36430
rect 16716 36418 16772 36428
rect 16380 35588 16436 35598
rect 16268 35586 16436 35588
rect 16268 35534 16382 35586
rect 16434 35534 16436 35586
rect 16268 35532 16436 35534
rect 16380 35522 16436 35532
rect 16044 34804 16100 34814
rect 15932 34802 16100 34804
rect 15932 34750 16046 34802
rect 16098 34750 16100 34802
rect 15932 34748 16100 34750
rect 16044 34738 16100 34748
rect 16380 34804 16436 34814
rect 16380 34802 16548 34804
rect 16380 34750 16382 34802
rect 16434 34750 16548 34802
rect 16380 34748 16548 34750
rect 16380 34738 16436 34748
rect 15708 34302 15710 34354
rect 15762 34302 15764 34354
rect 15708 34290 15764 34302
rect 16492 34018 16548 34748
rect 16940 34802 16996 36428
rect 18060 36482 18116 36494
rect 18060 36430 18062 36482
rect 18114 36430 18116 36482
rect 17500 36372 17556 36382
rect 17500 36278 17556 36316
rect 17836 35810 17892 35822
rect 17836 35758 17838 35810
rect 17890 35758 17892 35810
rect 16940 34750 16942 34802
rect 16994 34750 16996 34802
rect 16940 34738 16996 34750
rect 17164 34914 17220 34926
rect 17164 34862 17166 34914
rect 17218 34862 17220 34914
rect 16492 33966 16494 34018
rect 16546 33966 16548 34018
rect 16492 29428 16548 33966
rect 17052 34020 17108 34030
rect 17164 34020 17220 34862
rect 17052 34018 17220 34020
rect 17052 33966 17054 34018
rect 17106 33966 17220 34018
rect 17052 33964 17220 33966
rect 17500 34244 17556 34254
rect 17052 33236 17108 33964
rect 17500 33458 17556 34188
rect 17836 34244 17892 35758
rect 18060 35140 18116 36430
rect 18172 36372 18228 36382
rect 18172 35698 18228 36316
rect 18172 35646 18174 35698
rect 18226 35646 18228 35698
rect 18172 35634 18228 35646
rect 18284 36258 18340 36270
rect 18284 36206 18286 36258
rect 18338 36206 18340 36258
rect 18284 35476 18340 36206
rect 18284 35410 18340 35420
rect 18060 35084 18340 35140
rect 18060 34914 18116 34926
rect 18060 34862 18062 34914
rect 18114 34862 18116 34914
rect 18060 34354 18116 34862
rect 18060 34302 18062 34354
rect 18114 34302 18116 34354
rect 18060 34290 18116 34302
rect 17836 34178 17892 34188
rect 17500 33406 17502 33458
rect 17554 33406 17556 33458
rect 17500 33394 17556 33406
rect 17052 33170 17108 33180
rect 18284 33236 18340 35084
rect 18396 35028 18452 36988
rect 18956 36596 19012 39200
rect 19852 37156 19908 39200
rect 20748 39060 20804 39200
rect 21084 39060 21140 39228
rect 20748 39004 21140 39060
rect 19292 37100 19908 37156
rect 18956 36540 19236 36596
rect 18956 36370 19012 36382
rect 18956 36318 18958 36370
rect 19010 36318 19012 36370
rect 18956 35700 19012 36318
rect 18956 35634 19012 35644
rect 18620 35474 18676 35486
rect 18956 35476 19012 35486
rect 18620 35422 18622 35474
rect 18674 35422 18676 35474
rect 18508 35028 18564 35038
rect 18396 35026 18564 35028
rect 18396 34974 18510 35026
rect 18562 34974 18564 35026
rect 18396 34972 18564 34974
rect 18508 34962 18564 34972
rect 18396 34130 18452 34142
rect 18396 34078 18398 34130
rect 18450 34078 18452 34130
rect 18396 33460 18452 34078
rect 18620 33572 18676 35422
rect 18620 33506 18676 33516
rect 18844 35474 19012 35476
rect 18844 35422 18958 35474
rect 19010 35422 19012 35474
rect 18844 35420 19012 35422
rect 18396 33394 18452 33404
rect 18396 33236 18452 33246
rect 18284 33234 18452 33236
rect 18284 33182 18398 33234
rect 18450 33182 18452 33234
rect 18284 33180 18452 33182
rect 18284 32788 18340 33180
rect 18396 33170 18452 33180
rect 18284 31948 18340 32732
rect 16492 29362 16548 29372
rect 18172 31892 18340 31948
rect 18172 9380 18228 31892
rect 18172 9314 18228 9324
rect 14588 9202 14644 9212
rect 15708 7588 15764 7598
rect 14588 6468 14644 6478
rect 14588 6374 14644 6412
rect 15372 6466 15428 6478
rect 15372 6414 15374 6466
rect 15426 6414 15428 6466
rect 14252 4834 14308 4844
rect 15036 5236 15092 5246
rect 13692 4510 13694 4562
rect 13746 4510 13748 4562
rect 13692 4498 13748 4510
rect 12684 4386 12740 4396
rect 12908 4452 12964 4462
rect 12348 3614 12350 3666
rect 12402 3614 12404 3666
rect 12348 3602 12404 3614
rect 12908 3666 12964 4396
rect 14476 4228 14532 4238
rect 14476 4134 14532 4172
rect 14924 4226 14980 4238
rect 14924 4174 14926 4226
rect 14978 4174 14980 4226
rect 14924 4116 14980 4174
rect 14924 4050 14980 4060
rect 12908 3614 12910 3666
rect 12962 3614 12964 3666
rect 12908 3602 12964 3614
rect 11676 3444 11732 3454
rect 11676 3350 11732 3388
rect 13804 3444 13860 3454
rect 11340 3332 11396 3342
rect 11340 3238 11396 3276
rect 11228 3154 11284 3164
rect 13804 800 13860 3388
rect 14364 3444 14420 3454
rect 14364 3350 14420 3388
rect 15036 3332 15092 5180
rect 15372 4564 15428 6414
rect 15372 4498 15428 4508
rect 15484 6468 15540 6478
rect 15372 4340 15428 4350
rect 15036 3266 15092 3276
rect 15148 4338 15428 4340
rect 15148 4286 15374 4338
rect 15426 4286 15428 4338
rect 15148 4284 15428 4286
rect 15148 4228 15204 4284
rect 15372 4274 15428 4284
rect 15148 800 15204 4172
rect 15484 4116 15540 6412
rect 15708 4562 15764 7532
rect 18396 7364 18452 7374
rect 18284 7362 18452 7364
rect 18284 7310 18398 7362
rect 18450 7310 18452 7362
rect 18284 7308 18452 7310
rect 17612 6690 17668 6702
rect 17612 6638 17614 6690
rect 17666 6638 17668 6690
rect 16156 6132 16212 6142
rect 16156 6038 16212 6076
rect 17612 6132 17668 6638
rect 18284 6692 18340 7308
rect 18396 7298 18452 7308
rect 18284 6598 18340 6636
rect 17612 6066 17668 6076
rect 18732 6468 18788 6478
rect 17724 6020 17780 6030
rect 15932 5908 15988 5918
rect 15932 5814 15988 5852
rect 16716 5796 16772 5806
rect 16716 5234 16772 5740
rect 16716 5182 16718 5234
rect 16770 5182 16772 5234
rect 16716 5170 16772 5182
rect 16940 5794 16996 5806
rect 16940 5742 16942 5794
rect 16994 5742 16996 5794
rect 15708 4510 15710 4562
rect 15762 4510 15764 4562
rect 15708 4498 15764 4510
rect 16156 5122 16212 5134
rect 16156 5070 16158 5122
rect 16210 5070 16212 5122
rect 16156 4452 16212 5070
rect 16940 4788 16996 5742
rect 17500 5796 17556 5806
rect 17276 5124 17332 5134
rect 17276 5030 17332 5068
rect 16940 4722 16996 4732
rect 16156 4386 16212 4396
rect 16268 4676 16324 4686
rect 16268 4562 16324 4620
rect 16268 4510 16270 4562
rect 16322 4510 16324 4562
rect 16268 4340 16324 4510
rect 16828 4452 16884 4462
rect 16828 4358 16884 4396
rect 16268 4274 16324 4284
rect 16940 4228 16996 4238
rect 16940 4134 16996 4172
rect 15260 4060 15540 4116
rect 16492 4116 16548 4126
rect 15260 3554 15316 4060
rect 15260 3502 15262 3554
rect 15314 3502 15316 3554
rect 15260 3490 15316 3502
rect 16492 3554 16548 4060
rect 16492 3502 16494 3554
rect 16546 3502 16548 3554
rect 15932 3444 15988 3454
rect 15932 3350 15988 3388
rect 16492 800 16548 3502
rect 17500 3556 17556 5740
rect 17724 5122 17780 5964
rect 18732 6018 18788 6412
rect 18732 5966 18734 6018
rect 18786 5966 18788 6018
rect 18732 5954 18788 5966
rect 17836 5908 17892 5918
rect 17836 5814 17892 5852
rect 18172 5908 18228 5918
rect 18172 5814 18228 5852
rect 18844 5908 18900 35420
rect 18956 35410 19012 35420
rect 19180 34242 19236 36540
rect 19292 34916 19348 37100
rect 19622 36876 19886 36886
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19622 36810 19886 36820
rect 19740 36482 19796 36494
rect 19740 36430 19742 36482
rect 19794 36430 19796 36482
rect 19516 36372 19572 36382
rect 19516 36278 19572 36316
rect 19740 36148 19796 36430
rect 20188 36372 20244 36382
rect 20076 36260 20132 36270
rect 19516 35924 19572 35934
rect 19740 35924 19796 36092
rect 19516 35922 19796 35924
rect 19516 35870 19518 35922
rect 19570 35870 19796 35922
rect 19516 35868 19796 35870
rect 19964 36258 20132 36260
rect 19964 36206 20078 36258
rect 20130 36206 20132 36258
rect 19964 36204 20132 36206
rect 19516 35858 19572 35868
rect 19404 35476 19460 35486
rect 19404 35140 19460 35420
rect 19622 35308 19886 35318
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19622 35242 19886 35252
rect 19404 35084 19684 35140
rect 19292 34850 19348 34860
rect 19628 34914 19684 35084
rect 19628 34862 19630 34914
rect 19682 34862 19684 34914
rect 19628 34850 19684 34862
rect 19516 34804 19572 34814
rect 19516 34354 19572 34748
rect 19516 34302 19518 34354
rect 19570 34302 19572 34354
rect 19516 34290 19572 34302
rect 19180 34190 19182 34242
rect 19234 34190 19236 34242
rect 18956 33460 19012 33470
rect 19180 33460 19236 34190
rect 19622 33740 19886 33750
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19622 33674 19886 33684
rect 19852 33572 19908 33582
rect 18956 33458 19236 33460
rect 18956 33406 18958 33458
rect 19010 33406 19236 33458
rect 18956 33404 19236 33406
rect 19292 33460 19348 33470
rect 18956 33394 19012 33404
rect 19292 31220 19348 33404
rect 19852 33458 19908 33516
rect 19852 33406 19854 33458
rect 19906 33406 19908 33458
rect 19852 33124 19908 33406
rect 19852 33058 19908 33068
rect 19622 32172 19886 32182
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19622 32106 19886 32116
rect 19292 31154 19348 31164
rect 19622 30604 19886 30614
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19622 30538 19886 30548
rect 19622 29036 19886 29046
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19622 28970 19886 28980
rect 19622 27468 19886 27478
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19622 27402 19886 27412
rect 19622 25900 19886 25910
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19622 25834 19886 25844
rect 19622 24332 19886 24342
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19622 24266 19886 24276
rect 19622 22764 19886 22774
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19622 22698 19886 22708
rect 19622 21196 19886 21206
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19622 21130 19886 21140
rect 19622 19628 19886 19638
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19622 19562 19886 19572
rect 19622 18060 19886 18070
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19622 17994 19886 18004
rect 19622 16492 19886 16502
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19622 16426 19886 16436
rect 19622 14924 19886 14934
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19622 14858 19886 14868
rect 19622 13356 19886 13366
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19622 13290 19886 13300
rect 19622 11788 19886 11798
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19622 11722 19886 11732
rect 19622 10220 19886 10230
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19622 10154 19886 10164
rect 19622 8652 19886 8662
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19622 8586 19886 8596
rect 19292 7364 19348 7374
rect 19292 6804 19348 7308
rect 19622 7084 19886 7094
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19622 7018 19886 7028
rect 19628 6916 19684 6926
rect 19628 6822 19684 6860
rect 19964 6916 20020 36204
rect 20076 36194 20132 36204
rect 20076 35698 20132 35710
rect 20076 35646 20078 35698
rect 20130 35646 20132 35698
rect 20076 35364 20132 35646
rect 20076 35298 20132 35308
rect 20076 34356 20132 34366
rect 20076 34242 20132 34300
rect 20076 34190 20078 34242
rect 20130 34190 20132 34242
rect 20076 33684 20132 34190
rect 20076 33618 20132 33628
rect 20188 33124 20244 36316
rect 20748 36258 20804 36270
rect 20748 36206 20750 36258
rect 20802 36206 20804 36258
rect 20412 35812 20468 35822
rect 20412 35718 20468 35756
rect 20748 35364 20804 36206
rect 20748 35298 20804 35308
rect 20972 35698 21028 35710
rect 20972 35646 20974 35698
rect 21026 35646 21028 35698
rect 20300 35026 20356 35038
rect 20300 34974 20302 35026
rect 20354 34974 20356 35026
rect 20300 34916 20356 34974
rect 20300 34850 20356 34860
rect 20972 34354 21028 35646
rect 21420 35588 21476 39228
rect 21616 39200 21728 40000
rect 22512 39200 22624 40000
rect 23408 39200 23520 40000
rect 24304 39200 24416 40000
rect 25200 39200 25312 40000
rect 26096 39200 26208 40000
rect 26992 39200 27104 40000
rect 27888 39200 28000 40000
rect 28784 39200 28896 40000
rect 29680 39200 29792 40000
rect 30576 39200 30688 40000
rect 31472 39200 31584 40000
rect 32368 39200 32480 40000
rect 33264 39200 33376 40000
rect 34160 39200 34272 40000
rect 35056 39200 35168 40000
rect 35952 39200 36064 40000
rect 36848 39200 36960 40000
rect 37744 39200 37856 40000
rect 38640 39200 38752 40000
rect 39536 39200 39648 40000
rect 40432 39200 40544 40000
rect 41328 39200 41440 40000
rect 42224 39200 42336 40000
rect 43120 39200 43232 40000
rect 44016 39200 44128 40000
rect 44912 39200 45024 40000
rect 45808 39200 45920 40000
rect 46704 39200 46816 40000
rect 47600 39200 47712 40000
rect 48496 39200 48608 40000
rect 49392 39200 49504 40000
rect 50288 39200 50400 40000
rect 51184 39200 51296 40000
rect 52080 39200 52192 40000
rect 52976 39200 53088 40000
rect 53228 39228 53620 39284
rect 21644 36596 21700 39200
rect 21644 36530 21700 36540
rect 22204 36596 22260 36606
rect 22204 36502 22260 36540
rect 21756 36482 21812 36494
rect 21756 36430 21758 36482
rect 21810 36430 21812 36482
rect 21644 35588 21700 35598
rect 21420 35586 21700 35588
rect 21420 35534 21646 35586
rect 21698 35534 21700 35586
rect 21420 35532 21700 35534
rect 21644 35522 21700 35532
rect 21756 35364 21812 36430
rect 22092 35364 22148 35374
rect 21756 35308 21924 35364
rect 21868 34802 21924 35308
rect 21868 34750 21870 34802
rect 21922 34750 21924 34802
rect 21868 34738 21924 34750
rect 20972 34302 20974 34354
rect 21026 34302 21028 34354
rect 20972 34290 21028 34302
rect 20412 34244 20468 34254
rect 20412 34150 20468 34188
rect 21308 34130 21364 34142
rect 21308 34078 21310 34130
rect 21362 34078 21364 34130
rect 21308 33908 21364 34078
rect 21308 33842 21364 33852
rect 21756 34018 21812 34030
rect 21756 33966 21758 34018
rect 21810 33966 21812 34018
rect 21756 33908 21812 33966
rect 21756 33842 21812 33852
rect 20636 33684 20692 33694
rect 20636 33458 20692 33628
rect 20636 33406 20638 33458
rect 20690 33406 20692 33458
rect 20636 33394 20692 33406
rect 21756 33684 21812 33694
rect 20300 33124 20356 33134
rect 20188 33122 20356 33124
rect 20188 33070 20302 33122
rect 20354 33070 20356 33122
rect 20188 33068 20356 33070
rect 20300 32452 20356 33068
rect 20300 32386 20356 32396
rect 20300 7364 20356 7374
rect 20300 7270 20356 7308
rect 19964 6850 20020 6860
rect 20524 6916 20580 6926
rect 18844 5842 18900 5852
rect 18956 6748 19348 6804
rect 18956 5906 19012 6748
rect 18956 5854 18958 5906
rect 19010 5854 19012 5906
rect 18956 5842 19012 5854
rect 19068 6578 19124 6590
rect 19068 6526 19070 6578
rect 19122 6526 19124 6578
rect 19068 5348 19124 6526
rect 19292 6578 19348 6748
rect 20524 6690 20580 6860
rect 20524 6638 20526 6690
rect 20578 6638 20580 6690
rect 20524 6626 20580 6638
rect 19292 6526 19294 6578
rect 19346 6526 19348 6578
rect 19292 6514 19348 6526
rect 19964 6466 20020 6478
rect 19964 6414 19966 6466
rect 20018 6414 20020 6466
rect 19628 6020 19684 6030
rect 19628 5926 19684 5964
rect 19964 6018 20020 6414
rect 19964 5966 19966 6018
rect 20018 5966 20020 6018
rect 19964 5954 20020 5966
rect 21532 5908 21588 5918
rect 21532 5814 21588 5852
rect 20636 5796 20692 5806
rect 21196 5796 21252 5806
rect 20636 5794 21252 5796
rect 20636 5742 20638 5794
rect 20690 5742 21198 5794
rect 21250 5742 21252 5794
rect 20636 5740 21252 5742
rect 20524 5684 20580 5694
rect 20076 5682 20580 5684
rect 20076 5630 20526 5682
rect 20578 5630 20580 5682
rect 20076 5628 20580 5630
rect 19622 5516 19886 5526
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19622 5450 19886 5460
rect 19068 5282 19124 5292
rect 17724 5070 17726 5122
rect 17778 5070 17780 5122
rect 17724 5058 17780 5070
rect 20076 4898 20132 5628
rect 20524 5618 20580 5628
rect 20076 4846 20078 4898
rect 20130 4846 20132 4898
rect 20076 4834 20132 4846
rect 20300 5460 20356 5470
rect 20300 4900 20356 5404
rect 18172 4562 18228 4574
rect 18172 4510 18174 4562
rect 18226 4510 18228 4562
rect 17612 4340 17668 4350
rect 17612 4246 17668 4284
rect 17948 4340 18004 4350
rect 17612 3892 17668 3902
rect 17612 3778 17668 3836
rect 17612 3726 17614 3778
rect 17666 3726 17668 3778
rect 17612 3714 17668 3726
rect 17948 3778 18004 4284
rect 18172 4228 18228 4510
rect 18172 4162 18228 4172
rect 18732 4564 18788 4574
rect 17948 3726 17950 3778
rect 18002 3726 18004 3778
rect 17948 3714 18004 3726
rect 18732 3778 18788 4508
rect 20300 4228 20356 4844
rect 20636 4788 20692 5740
rect 21196 5730 21252 5740
rect 20300 4162 20356 4172
rect 20412 4732 20692 4788
rect 20748 5348 20804 5358
rect 20412 4452 20468 4732
rect 19622 3948 19886 3958
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19622 3882 19886 3892
rect 18732 3726 18734 3778
rect 18786 3726 18788 3778
rect 18732 3714 18788 3726
rect 19628 3668 19684 3678
rect 19180 3666 19684 3668
rect 19180 3614 19630 3666
rect 19682 3614 19684 3666
rect 19180 3612 19684 3614
rect 17612 3556 17668 3566
rect 17500 3554 17668 3556
rect 17500 3502 17614 3554
rect 17666 3502 17668 3554
rect 17500 3500 17668 3502
rect 17612 3490 17668 3500
rect 18844 3444 18900 3454
rect 18844 3350 18900 3388
rect 16716 3332 16772 3342
rect 16716 3238 16772 3276
rect 19180 800 19236 3612
rect 19628 3602 19684 3612
rect 20412 3668 20468 4396
rect 20412 3602 20468 3612
rect 20524 4340 20580 4350
rect 20524 800 20580 4284
rect 20636 4338 20692 4350
rect 20636 4286 20638 4338
rect 20690 4286 20692 4338
rect 20636 4228 20692 4286
rect 20636 4162 20692 4172
rect 20636 3556 20692 3566
rect 20748 3556 20804 5292
rect 21532 5124 21588 5134
rect 21308 5068 21532 5124
rect 21308 4340 21364 5068
rect 21532 5030 21588 5068
rect 21756 4562 21812 33628
rect 22092 31948 22148 35308
rect 22540 34916 22596 39200
rect 23100 38500 23156 38510
rect 23100 35922 23156 38444
rect 23100 35870 23102 35922
rect 23154 35870 23156 35922
rect 23100 35858 23156 35870
rect 22876 35698 22932 35710
rect 22876 35646 22878 35698
rect 22930 35646 22932 35698
rect 22764 34916 22820 34926
rect 22540 34914 22820 34916
rect 22540 34862 22766 34914
rect 22818 34862 22820 34914
rect 22540 34860 22820 34862
rect 22204 34802 22260 34814
rect 22204 34750 22206 34802
rect 22258 34750 22260 34802
rect 22204 34020 22260 34750
rect 22764 34356 22820 34860
rect 22876 34580 22932 35646
rect 23436 35588 23492 39200
rect 24332 37828 24388 39200
rect 23884 37772 24388 37828
rect 23884 36594 23940 37772
rect 23884 36542 23886 36594
rect 23938 36542 23940 36594
rect 23884 36530 23940 36542
rect 24444 36482 24500 36494
rect 24444 36430 24446 36482
rect 24498 36430 24500 36482
rect 24220 36148 24276 36158
rect 23436 35522 23492 35532
rect 23660 35698 23716 35710
rect 23660 35646 23662 35698
rect 23714 35646 23716 35698
rect 23100 35252 23156 35262
rect 23100 34802 23156 35196
rect 23100 34750 23102 34802
rect 23154 34750 23156 34802
rect 23100 34738 23156 34750
rect 23660 34802 23716 35646
rect 23996 35364 24052 35374
rect 24220 35364 24276 36092
rect 24332 35588 24388 35598
rect 24332 35494 24388 35532
rect 24220 35308 24388 35364
rect 23996 34916 24052 35308
rect 23996 34914 24276 34916
rect 23996 34862 23998 34914
rect 24050 34862 24276 34914
rect 23996 34860 24276 34862
rect 23996 34850 24052 34860
rect 23660 34750 23662 34802
rect 23714 34750 23716 34802
rect 23660 34738 23716 34750
rect 22876 34514 22932 34524
rect 23324 34468 23380 34478
rect 22876 34356 22932 34366
rect 22764 34354 22932 34356
rect 22764 34302 22878 34354
rect 22930 34302 22932 34354
rect 22764 34300 22932 34302
rect 22876 34290 22932 34300
rect 23324 34354 23380 34412
rect 23324 34302 23326 34354
rect 23378 34302 23380 34354
rect 23324 34290 23380 34302
rect 24220 34354 24276 34860
rect 24220 34302 24222 34354
rect 24274 34302 24276 34354
rect 24220 34290 24276 34302
rect 22428 34020 22484 34030
rect 22204 34018 22484 34020
rect 22204 33966 22430 34018
rect 22482 33966 22484 34018
rect 22204 33964 22484 33966
rect 22428 33796 22484 33964
rect 22428 33730 22484 33740
rect 22092 31892 22260 31948
rect 22204 8428 22260 31892
rect 24332 25732 24388 35308
rect 24444 34804 24500 36430
rect 25228 34916 25284 39200
rect 25788 36820 25844 36830
rect 25676 35586 25732 35598
rect 25676 35534 25678 35586
rect 25730 35534 25732 35586
rect 25676 35476 25732 35534
rect 25676 35410 25732 35420
rect 25452 34916 25508 34926
rect 25228 34914 25508 34916
rect 25228 34862 25454 34914
rect 25506 34862 25508 34914
rect 25228 34860 25508 34862
rect 24556 34804 24612 34814
rect 24444 34802 24612 34804
rect 24444 34750 24558 34802
rect 24610 34750 24612 34802
rect 24444 34748 24612 34750
rect 24556 34738 24612 34748
rect 24892 34802 24948 34814
rect 24892 34750 24894 34802
rect 24946 34750 24948 34802
rect 24892 34132 24948 34750
rect 25452 34356 25508 34860
rect 25788 34802 25844 36764
rect 26012 36596 26068 36606
rect 26124 36596 26180 39200
rect 26012 36594 26180 36596
rect 26012 36542 26014 36594
rect 26066 36542 26180 36594
rect 26012 36540 26180 36542
rect 26572 37604 26628 37614
rect 26012 36530 26068 36540
rect 26460 36482 26516 36494
rect 26460 36430 26462 36482
rect 26514 36430 26516 36482
rect 26236 35698 26292 35710
rect 26236 35646 26238 35698
rect 26290 35646 26292 35698
rect 25788 34750 25790 34802
rect 25842 34750 25844 34802
rect 25788 34738 25844 34750
rect 25900 35476 25956 35486
rect 25452 34290 25508 34300
rect 24892 34066 24948 34076
rect 25004 34244 25060 34254
rect 25004 30996 25060 34188
rect 25564 34132 25620 34142
rect 25564 34038 25620 34076
rect 25004 30930 25060 30940
rect 25116 31220 25172 31230
rect 24332 25666 24388 25676
rect 25116 25620 25172 31164
rect 25116 8428 25172 25564
rect 25900 20188 25956 35420
rect 26236 35476 26292 35646
rect 26236 35410 26292 35420
rect 26460 34804 26516 36430
rect 26572 35922 26628 37548
rect 26572 35870 26574 35922
rect 26626 35870 26628 35922
rect 26572 35858 26628 35870
rect 27020 35588 27076 39200
rect 27804 36596 27860 36606
rect 27804 36502 27860 36540
rect 27916 35812 27972 39200
rect 27692 35756 27972 35812
rect 28364 37268 28420 37278
rect 27356 35588 27412 35598
rect 27020 35586 27412 35588
rect 27020 35534 27358 35586
rect 27410 35534 27412 35586
rect 27020 35532 27412 35534
rect 27356 35522 27412 35532
rect 26572 34804 26628 34814
rect 26460 34802 26628 34804
rect 26460 34750 26574 34802
rect 26626 34750 26628 34802
rect 26460 34748 26628 34750
rect 26572 34738 26628 34748
rect 26908 34802 26964 34814
rect 26908 34750 26910 34802
rect 26962 34750 26964 34802
rect 26012 34356 26068 34366
rect 26012 34262 26068 34300
rect 26908 34020 26964 34750
rect 27692 34356 27748 35756
rect 28140 35700 28196 35710
rect 27804 35698 28196 35700
rect 27804 35646 28142 35698
rect 28194 35646 28196 35698
rect 27804 35644 28196 35646
rect 27804 34802 27860 35644
rect 28140 35634 28196 35644
rect 27804 34750 27806 34802
rect 27858 34750 27860 34802
rect 27804 34738 27860 34750
rect 28140 34804 28196 34814
rect 28140 34710 28196 34748
rect 28364 34356 28420 37212
rect 28812 36596 28868 39200
rect 28812 36530 28868 36540
rect 28476 36484 28532 36494
rect 28476 36390 28532 36428
rect 29596 36484 29652 36494
rect 29484 36370 29540 36382
rect 29484 36318 29486 36370
rect 29538 36318 29540 36370
rect 29372 35700 29428 35710
rect 29372 35606 29428 35644
rect 29036 35476 29092 35486
rect 28924 35474 29092 35476
rect 28924 35422 29038 35474
rect 29090 35422 29092 35474
rect 28924 35420 29092 35422
rect 28700 34804 28756 34814
rect 28700 34690 28756 34748
rect 28700 34638 28702 34690
rect 28754 34638 28756 34690
rect 28476 34356 28532 34366
rect 27692 34354 28196 34356
rect 27692 34302 27694 34354
rect 27746 34302 28196 34354
rect 27692 34300 28196 34302
rect 28364 34354 28532 34356
rect 28364 34302 28478 34354
rect 28530 34302 28532 34354
rect 28364 34300 28532 34302
rect 27692 34290 27748 34300
rect 28140 34242 28196 34300
rect 28476 34290 28532 34300
rect 28700 34356 28756 34638
rect 28700 34290 28756 34300
rect 28140 34190 28142 34242
rect 28194 34190 28196 34242
rect 28140 34178 28196 34190
rect 27132 34020 27188 34030
rect 26908 34018 27188 34020
rect 26908 33966 27134 34018
rect 27186 33966 27188 34018
rect 26908 33964 27188 33966
rect 27132 33572 27188 33964
rect 27132 33506 27188 33516
rect 28364 33124 28420 33134
rect 26908 29428 26964 29438
rect 26908 26516 26964 29372
rect 28364 27636 28420 33068
rect 28364 27570 28420 27580
rect 26908 26450 26964 26460
rect 27804 26516 27860 26526
rect 25900 20132 26292 20188
rect 21756 4510 21758 4562
rect 21810 4510 21812 4562
rect 21756 4498 21812 4510
rect 21980 8372 22260 8428
rect 25004 8372 25172 8428
rect 21308 4338 21588 4340
rect 21308 4286 21310 4338
rect 21362 4286 21588 4338
rect 21308 4284 21588 4286
rect 21308 4274 21364 4284
rect 21532 3666 21588 4284
rect 21532 3614 21534 3666
rect 21586 3614 21588 3666
rect 21532 3602 21588 3614
rect 20636 3554 20804 3556
rect 20636 3502 20638 3554
rect 20690 3502 20804 3554
rect 20636 3500 20804 3502
rect 20636 3490 20692 3500
rect 21980 3332 22036 8372
rect 22092 4900 22148 4910
rect 25004 4900 25060 8372
rect 26124 6468 26180 6478
rect 25564 6466 26180 6468
rect 25564 6414 26126 6466
rect 26178 6414 26180 6466
rect 25564 6412 26180 6414
rect 25116 5124 25172 5134
rect 25116 5030 25172 5068
rect 25564 5122 25620 6412
rect 26124 6402 26180 6412
rect 25564 5070 25566 5122
rect 25618 5070 25620 5122
rect 25564 5058 25620 5070
rect 22092 4898 22260 4900
rect 22092 4846 22094 4898
rect 22146 4846 22260 4898
rect 22092 4844 22260 4846
rect 25004 4844 25172 4900
rect 22092 4834 22148 4844
rect 22092 4340 22148 4350
rect 22092 4246 22148 4284
rect 22204 3556 22260 4844
rect 22540 4340 22596 4350
rect 22540 4246 22596 4284
rect 25004 4228 25060 4238
rect 25004 4134 25060 4172
rect 22316 3556 22372 3566
rect 22204 3554 22372 3556
rect 22204 3502 22318 3554
rect 22370 3502 22372 3554
rect 22204 3500 22372 3502
rect 22092 3332 22148 3342
rect 21980 3330 22148 3332
rect 21980 3278 22094 3330
rect 22146 3278 22148 3330
rect 21980 3276 22148 3278
rect 22092 3266 22148 3276
rect 22316 2772 22372 3500
rect 22988 3444 23044 3454
rect 23436 3444 23492 3454
rect 22988 3442 23492 3444
rect 22988 3390 22990 3442
rect 23042 3390 23438 3442
rect 23490 3390 23492 3442
rect 22988 3388 23492 3390
rect 22988 3378 23044 3388
rect 21868 2716 22372 2772
rect 21868 800 21924 2716
rect 23212 800 23268 3388
rect 23436 3378 23492 3388
rect 24556 3444 24612 3454
rect 23772 3330 23828 3342
rect 23772 3278 23774 3330
rect 23826 3278 23828 3330
rect 23772 3220 23828 3278
rect 23772 3154 23828 3164
rect 24556 800 24612 3388
rect 25116 3220 25172 4844
rect 26124 4340 26180 4350
rect 25900 4338 26180 4340
rect 25900 4286 26126 4338
rect 26178 4286 26180 4338
rect 25900 4284 26180 4286
rect 25676 4226 25732 4238
rect 25676 4174 25678 4226
rect 25730 4174 25732 4226
rect 25676 4116 25732 4174
rect 25676 4050 25732 4060
rect 25900 4228 25956 4284
rect 26124 4274 26180 4284
rect 25676 3444 25732 3454
rect 25676 3350 25732 3388
rect 25116 3154 25172 3164
rect 25900 800 25956 4172
rect 26236 3332 26292 20132
rect 26460 9268 26516 9278
rect 26348 7250 26404 7262
rect 26348 7198 26350 7250
rect 26402 7198 26404 7250
rect 26348 6690 26404 7198
rect 26348 6638 26350 6690
rect 26402 6638 26404 6690
rect 26348 6626 26404 6638
rect 26460 4562 26516 9212
rect 26460 4510 26462 4562
rect 26514 4510 26516 4562
rect 26460 4498 26516 4510
rect 26572 7588 26628 7598
rect 26572 5236 26628 7532
rect 26908 7586 26964 7598
rect 26908 7534 26910 7586
rect 26962 7534 26964 7586
rect 26684 7476 26740 7486
rect 26684 7382 26740 7420
rect 26908 7364 26964 7534
rect 27244 7588 27300 7598
rect 27244 7494 27300 7532
rect 26908 7298 26964 7308
rect 27132 7252 27188 7262
rect 27132 6690 27188 7196
rect 27132 6638 27134 6690
rect 27186 6638 27188 6690
rect 27132 6626 27188 6638
rect 27692 6692 27748 6702
rect 27356 6468 27412 6478
rect 27356 6374 27412 6412
rect 27692 6020 27748 6636
rect 27692 5906 27748 5964
rect 27692 5854 27694 5906
rect 27746 5854 27748 5906
rect 27692 5842 27748 5854
rect 26572 3554 26628 5180
rect 27132 4564 27188 4574
rect 27132 4450 27188 4508
rect 27132 4398 27134 4450
rect 27186 4398 27188 4450
rect 27132 4386 27188 4398
rect 27468 4452 27524 4462
rect 27468 4358 27524 4396
rect 26572 3502 26574 3554
rect 26626 3502 26628 3554
rect 26572 3490 26628 3502
rect 27244 4116 27300 4126
rect 26236 3266 26292 3276
rect 27244 3444 27300 4060
rect 27468 3444 27524 3454
rect 27244 3442 27524 3444
rect 27244 3390 27470 3442
rect 27522 3390 27524 3442
rect 27244 3388 27524 3390
rect 27244 800 27300 3388
rect 27468 3378 27524 3388
rect 27804 3330 27860 26460
rect 28028 8036 28084 8046
rect 28028 7476 28084 7980
rect 28588 8036 28644 8046
rect 28924 8036 28980 35420
rect 29036 35410 29092 35420
rect 29372 34916 29428 34926
rect 29484 34916 29540 36318
rect 29428 34860 29540 34916
rect 29036 34692 29092 34702
rect 29036 34354 29092 34636
rect 29036 34302 29038 34354
rect 29090 34302 29092 34354
rect 29036 34290 29092 34302
rect 29372 34354 29428 34860
rect 29596 34802 29652 36428
rect 29708 35588 29764 39200
rect 30156 37828 30212 37838
rect 30156 36708 30212 37772
rect 30156 36576 30212 36652
rect 29708 35522 29764 35532
rect 29820 36370 29876 36382
rect 29820 36318 29822 36370
rect 29874 36318 29876 36370
rect 29820 35698 29876 36318
rect 30492 36260 30548 36270
rect 30268 36258 30548 36260
rect 30268 36206 30494 36258
rect 30546 36206 30548 36258
rect 30268 36204 30548 36206
rect 29820 35646 29822 35698
rect 29874 35646 29876 35698
rect 29820 35140 29876 35646
rect 30156 35810 30212 35822
rect 30156 35758 30158 35810
rect 30210 35758 30212 35810
rect 29820 35084 30100 35140
rect 29596 34750 29598 34802
rect 29650 34750 29652 34802
rect 29596 34738 29652 34750
rect 29932 34916 29988 34926
rect 29372 34302 29374 34354
rect 29426 34302 29428 34354
rect 29372 34290 29428 34302
rect 29820 34356 29876 34366
rect 29932 34356 29988 34860
rect 29820 34354 29988 34356
rect 29820 34302 29822 34354
rect 29874 34302 29988 34354
rect 29820 34300 29988 34302
rect 29820 34290 29876 34300
rect 30044 33460 30100 35084
rect 30156 34692 30212 35758
rect 30156 34626 30212 34636
rect 30044 33394 30100 33404
rect 30268 31948 30324 36204
rect 30492 36194 30548 36204
rect 30604 35812 30660 39200
rect 31500 36594 31556 39200
rect 31500 36542 31502 36594
rect 31554 36542 31556 36594
rect 31500 36530 31556 36542
rect 31724 36708 31780 36718
rect 30380 35756 30660 35812
rect 30380 34356 30436 35756
rect 30828 35698 30884 35710
rect 30828 35646 30830 35698
rect 30882 35646 30884 35698
rect 30604 35140 30660 35150
rect 30604 34914 30660 35084
rect 30604 34862 30606 34914
rect 30658 34862 30660 34914
rect 30604 34850 30660 34862
rect 30828 34802 30884 35646
rect 31500 35588 31556 35598
rect 31500 35494 31556 35532
rect 31388 35140 31444 35150
rect 31388 35026 31444 35084
rect 31388 34974 31390 35026
rect 31442 34974 31444 35026
rect 31388 34962 31444 34974
rect 30828 34750 30830 34802
rect 30882 34750 30884 34802
rect 30828 34738 30884 34750
rect 30380 34354 30884 34356
rect 30380 34302 30382 34354
rect 30434 34302 30884 34354
rect 30380 34300 30884 34302
rect 30380 34290 30436 34300
rect 30828 34242 30884 34300
rect 31724 34354 31780 36652
rect 31836 36484 31892 36494
rect 31836 34802 31892 36428
rect 32172 36484 32228 36494
rect 32172 36390 32228 36428
rect 32396 35812 32452 39200
rect 32396 35746 32452 35756
rect 32620 35700 32676 35710
rect 32620 35586 32676 35644
rect 32620 35534 32622 35586
rect 32674 35534 32676 35586
rect 31836 34750 31838 34802
rect 31890 34750 31892 34802
rect 31836 34738 31892 34750
rect 32172 34802 32228 34814
rect 32172 34750 32174 34802
rect 32226 34750 32228 34802
rect 31724 34302 31726 34354
rect 31778 34302 31780 34354
rect 31724 34290 31780 34302
rect 30828 34190 30830 34242
rect 30882 34190 30884 34242
rect 30828 34178 30884 34190
rect 31164 34242 31220 34254
rect 31164 34190 31166 34242
rect 31218 34190 31220 34242
rect 30604 33460 30660 33470
rect 30604 33366 30660 33404
rect 31052 33460 31108 33470
rect 31052 33366 31108 33404
rect 31164 33348 31220 34190
rect 32172 34020 32228 34750
rect 32396 34020 32452 34030
rect 32172 34018 32452 34020
rect 32172 33966 32398 34018
rect 32450 33966 32452 34018
rect 32172 33964 32452 33966
rect 31164 33282 31220 33292
rect 30268 31892 30436 31948
rect 28588 8034 28756 8036
rect 28588 7982 28590 8034
rect 28642 7982 28756 8034
rect 28588 7980 28756 7982
rect 28588 7970 28644 7980
rect 28700 7588 28756 7980
rect 28924 7970 28980 7980
rect 28812 7588 28868 7598
rect 28700 7586 28868 7588
rect 28700 7534 28814 7586
rect 28866 7534 28868 7586
rect 28700 7532 28868 7534
rect 28028 7410 28084 7420
rect 28588 7476 28644 7486
rect 28588 7382 28644 7420
rect 28364 7364 28420 7374
rect 28252 7252 28308 7262
rect 28252 7158 28308 7196
rect 28364 6802 28420 7308
rect 28812 7364 28868 7532
rect 28812 7298 28868 7308
rect 29372 7586 29428 7598
rect 29372 7534 29374 7586
rect 29426 7534 29428 7586
rect 28364 6750 28366 6802
rect 28418 6750 28420 6802
rect 28364 6738 28420 6750
rect 27916 6580 27972 6590
rect 27916 6466 27972 6524
rect 27916 6414 27918 6466
rect 27970 6414 27972 6466
rect 27916 5460 27972 6414
rect 28252 6468 28308 6478
rect 28252 5906 28308 6412
rect 29372 6244 29428 7534
rect 30380 7476 30436 31892
rect 32396 9268 32452 33964
rect 32620 26404 32676 35534
rect 32844 34916 32900 34926
rect 32844 34822 32900 34860
rect 33292 34916 33348 39200
rect 34188 37828 34244 39200
rect 34188 37772 34692 37828
rect 33852 37044 33908 37054
rect 33516 36596 33572 36606
rect 33516 36482 33572 36540
rect 33516 36430 33518 36482
rect 33570 36430 33572 36482
rect 33516 36418 33572 36430
rect 33852 36370 33908 36988
rect 34636 36594 34692 37772
rect 34636 36542 34638 36594
rect 34690 36542 34692 36594
rect 34636 36530 34692 36542
rect 35084 36596 35140 39200
rect 35980 36706 36036 39200
rect 35980 36654 35982 36706
rect 36034 36654 36036 36706
rect 35980 36642 36036 36654
rect 36540 36706 36596 36718
rect 36540 36654 36542 36706
rect 36594 36654 36596 36706
rect 35084 36530 35140 36540
rect 36092 36596 36148 36606
rect 36092 36502 36148 36540
rect 33852 36318 33854 36370
rect 33906 36318 33908 36370
rect 33852 36306 33908 36318
rect 35532 36482 35588 36494
rect 35532 36430 35534 36482
rect 35586 36430 35588 36482
rect 34524 35812 34580 35822
rect 34524 35718 34580 35756
rect 33068 34690 33124 34702
rect 33068 34638 33070 34690
rect 33122 34638 33124 34690
rect 33068 31892 33124 34638
rect 33292 34356 33348 34860
rect 33628 35698 33684 35710
rect 33628 35646 33630 35698
rect 33682 35646 33684 35698
rect 33628 34802 33684 35646
rect 33628 34750 33630 34802
rect 33682 34750 33684 34802
rect 33628 34738 33684 34750
rect 33964 34802 34020 34814
rect 33964 34750 33966 34802
rect 34018 34750 34020 34802
rect 33516 34356 33572 34366
rect 33292 34354 33572 34356
rect 33292 34302 33518 34354
rect 33570 34302 33572 34354
rect 33292 34300 33572 34302
rect 33516 34290 33572 34300
rect 33964 34020 34020 34750
rect 34524 34802 34580 34814
rect 34524 34750 34526 34802
rect 34578 34750 34580 34802
rect 34188 34020 34244 34030
rect 33964 34018 34244 34020
rect 33964 33966 34190 34018
rect 34242 33966 34244 34018
rect 33964 33964 34244 33966
rect 34188 33684 34244 33964
rect 34188 33618 34244 33628
rect 34524 34020 34580 34750
rect 35532 34802 35588 36430
rect 36316 35924 36372 35934
rect 35532 34750 35534 34802
rect 35586 34750 35588 34802
rect 35532 34738 35588 34750
rect 35868 34802 35924 34814
rect 35868 34750 35870 34802
rect 35922 34750 35924 34802
rect 33068 31826 33124 31836
rect 32620 26338 32676 26348
rect 32396 9202 32452 9212
rect 33516 9380 33572 9390
rect 30380 7382 30436 7420
rect 29932 7364 29988 7374
rect 29932 7270 29988 7308
rect 29596 6580 29652 6590
rect 29596 6486 29652 6524
rect 29372 6178 29428 6188
rect 31388 6244 31444 6254
rect 31388 6130 31444 6188
rect 31388 6078 31390 6130
rect 31442 6078 31444 6130
rect 28252 5854 28254 5906
rect 28306 5854 28308 5906
rect 28252 5842 28308 5854
rect 30604 6018 30660 6030
rect 30604 5966 30606 6018
rect 30658 5966 30660 6018
rect 27916 5394 27972 5404
rect 29708 5348 29764 5358
rect 29708 5254 29764 5292
rect 30604 5348 30660 5966
rect 30604 5282 30660 5292
rect 28588 5236 28644 5246
rect 28588 5142 28644 5180
rect 28700 5124 28756 5134
rect 28028 4898 28084 4910
rect 28028 4846 28030 4898
rect 28082 4846 28084 4898
rect 28028 4562 28084 4846
rect 28028 4510 28030 4562
rect 28082 4510 28084 4562
rect 28028 4498 28084 4510
rect 28700 4562 28756 5068
rect 29596 5010 29652 5022
rect 29596 4958 29598 5010
rect 29650 4958 29652 5010
rect 29596 4900 29652 4958
rect 28700 4510 28702 4562
rect 28754 4510 28756 4562
rect 28700 4498 28756 4510
rect 29148 4564 29204 4574
rect 28140 4452 28196 4462
rect 28140 4358 28196 4396
rect 29148 4116 29204 4508
rect 29596 4452 29652 4844
rect 30156 4900 30212 4910
rect 30156 4806 30212 4844
rect 29596 4358 29652 4396
rect 29148 4050 29204 4060
rect 31388 3554 31444 6078
rect 31724 6020 31780 6030
rect 31724 5926 31780 5964
rect 31724 4228 31780 4238
rect 31724 4226 31892 4228
rect 31724 4174 31726 4226
rect 31778 4174 31892 4226
rect 31724 4172 31892 4174
rect 31724 4162 31780 4172
rect 31388 3502 31390 3554
rect 31442 3502 31444 3554
rect 31388 3490 31444 3502
rect 27804 3278 27806 3330
rect 27858 3278 27860 3330
rect 27804 3266 27860 3278
rect 28588 3444 28644 3454
rect 28588 800 28644 3388
rect 29596 3444 29652 3454
rect 29596 3350 29652 3388
rect 29932 3444 29988 3454
rect 29260 3332 29316 3342
rect 29260 3238 29316 3276
rect 29932 800 29988 3388
rect 30492 3444 30548 3454
rect 30492 3350 30548 3388
rect 31276 3444 31332 3454
rect 31276 800 31332 3388
rect 31836 3444 31892 4172
rect 32956 4226 33012 4238
rect 32956 4174 32958 4226
rect 33010 4174 33012 4226
rect 31948 3444 32004 3454
rect 31892 3442 32004 3444
rect 31892 3390 31950 3442
rect 32002 3390 32004 3442
rect 31892 3388 32004 3390
rect 31836 3378 31892 3388
rect 31948 3378 32004 3388
rect 32620 3444 32676 3454
rect 32284 3330 32340 3342
rect 32284 3278 32286 3330
rect 32338 3278 32340 3330
rect 32284 3220 32340 3278
rect 32284 3154 32340 3164
rect 32620 800 32676 3388
rect 32956 3444 33012 4174
rect 32956 3378 33012 3388
rect 33180 3444 33236 3454
rect 33180 3350 33236 3388
rect 33516 3330 33572 9324
rect 33516 3278 33518 3330
rect 33570 3278 33572 3330
rect 33516 3266 33572 3278
rect 33964 4226 34020 4238
rect 33964 4174 33966 4226
rect 34018 4174 34020 4226
rect 33964 3444 34020 4174
rect 34188 3444 34244 3454
rect 33964 3442 34244 3444
rect 33964 3390 34190 3442
rect 34242 3390 34244 3442
rect 33964 3388 34244 3390
rect 33964 800 34020 3388
rect 34188 3378 34244 3388
rect 34524 3330 34580 33964
rect 34860 34690 34916 34702
rect 34860 34638 34862 34690
rect 34914 34638 34916 34690
rect 34860 29204 34916 34638
rect 35084 34020 35140 34030
rect 35868 34020 35924 34750
rect 36092 34020 36148 34030
rect 35868 34018 36148 34020
rect 35868 33966 36094 34018
rect 36146 33966 36148 34018
rect 35868 33964 36148 33966
rect 35084 33926 35140 33964
rect 34860 29138 34916 29148
rect 36092 11620 36148 33964
rect 36316 29316 36372 35868
rect 36540 35810 36596 36654
rect 36540 35758 36542 35810
rect 36594 35758 36596 35810
rect 36540 35746 36596 35758
rect 36540 34916 36596 34926
rect 36876 34916 36932 39200
rect 37772 36594 37828 39200
rect 37772 36542 37774 36594
rect 37826 36542 37828 36594
rect 37772 36530 37828 36542
rect 38444 36484 38500 36494
rect 38444 36390 38500 36428
rect 38032 36092 38296 36102
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38032 36026 38296 36036
rect 38668 35924 38724 39200
rect 38556 35868 38724 35924
rect 39004 38388 39060 38398
rect 39004 35922 39060 38332
rect 39564 36594 39620 39200
rect 39564 36542 39566 36594
rect 39618 36542 39620 36594
rect 39564 36530 39620 36542
rect 39004 35870 39006 35922
rect 39058 35870 39060 35922
rect 36540 34914 36932 34916
rect 36540 34862 36542 34914
rect 36594 34862 36932 34914
rect 36540 34860 36932 34862
rect 36540 34850 36596 34860
rect 36764 34690 36820 34702
rect 36764 34638 36766 34690
rect 36818 34638 36820 34690
rect 36764 32564 36820 34638
rect 36876 34354 36932 34860
rect 36876 34302 36878 34354
rect 36930 34302 36932 34354
rect 36876 34290 36932 34302
rect 37436 35698 37492 35710
rect 37436 35646 37438 35698
rect 37490 35646 37492 35698
rect 37436 34354 37492 35646
rect 37436 34302 37438 34354
rect 37490 34302 37492 34354
rect 37436 34290 37492 34302
rect 37548 35588 37604 35598
rect 37548 34132 37604 35532
rect 38108 35588 38164 35598
rect 38108 35494 38164 35532
rect 37772 34916 37828 34926
rect 37772 34822 37828 34860
rect 38332 34916 38388 34926
rect 38556 34916 38612 35868
rect 39004 35858 39060 35870
rect 39116 36484 39172 36494
rect 38388 34860 38612 34916
rect 38668 35698 38724 35710
rect 38668 35646 38670 35698
rect 38722 35646 38724 35698
rect 38332 34784 38388 34860
rect 38556 34692 38612 34702
rect 38444 34690 38612 34692
rect 38444 34638 38558 34690
rect 38610 34638 38612 34690
rect 38444 34636 38612 34638
rect 38032 34524 38296 34534
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38032 34458 38296 34468
rect 37548 34066 37604 34076
rect 37772 34132 37828 34142
rect 37772 34130 37940 34132
rect 37772 34078 37774 34130
rect 37826 34078 37940 34130
rect 37772 34076 37940 34078
rect 37772 34066 37828 34076
rect 36764 32498 36820 32508
rect 37436 33796 37492 33806
rect 36316 29250 36372 29260
rect 36092 11554 36148 11564
rect 36316 4228 36372 4238
rect 34524 3278 34526 3330
rect 34578 3278 34580 3330
rect 34524 3266 34580 3278
rect 35308 3666 35364 3678
rect 35308 3614 35310 3666
rect 35362 3614 35364 3666
rect 35308 800 35364 3614
rect 36316 3554 36372 4172
rect 36316 3502 36318 3554
rect 36370 3502 36372 3554
rect 36316 3490 36372 3502
rect 36876 4226 36932 4238
rect 36876 4174 36878 4226
rect 36930 4174 36932 4226
rect 36876 3444 36932 4174
rect 37212 4228 37268 4238
rect 37212 4134 37268 4172
rect 37100 3444 37156 3454
rect 36652 3442 37156 3444
rect 36652 3390 37102 3442
rect 37154 3390 37156 3442
rect 36652 3388 37156 3390
rect 36652 800 36708 3388
rect 37100 3378 37156 3388
rect 37436 3330 37492 33740
rect 37436 3278 37438 3330
rect 37490 3278 37492 3330
rect 37436 3266 37492 3278
rect 37772 33236 37828 33246
rect 37772 3332 37828 33180
rect 37884 33124 37940 34076
rect 38444 33348 38500 34636
rect 38556 34626 38612 34636
rect 38556 34018 38612 34030
rect 38556 33966 38558 34018
rect 38610 33966 38612 34018
rect 38556 33796 38612 33966
rect 38556 33730 38612 33740
rect 38444 33292 38612 33348
rect 38332 33236 38388 33246
rect 38388 33180 38500 33236
rect 38332 33170 38388 33180
rect 37996 33124 38052 33162
rect 37884 33068 37996 33124
rect 37996 33058 38052 33068
rect 38444 33122 38500 33180
rect 38444 33070 38446 33122
rect 38498 33070 38500 33122
rect 38444 33058 38500 33070
rect 38032 32956 38296 32966
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38032 32890 38296 32900
rect 38556 32900 38612 33292
rect 38668 33236 38724 35646
rect 39116 34802 39172 36428
rect 40236 36484 40292 36494
rect 40236 36390 40292 36428
rect 40460 35924 40516 39200
rect 41356 36594 41412 39200
rect 41356 36542 41358 36594
rect 41410 36542 41412 36594
rect 41356 36530 41412 36542
rect 41804 36820 41860 36830
rect 40348 35868 40516 35924
rect 40908 36484 40964 36494
rect 39900 35812 39956 35822
rect 39900 35718 39956 35756
rect 39564 35698 39620 35710
rect 39564 35646 39566 35698
rect 39618 35646 39620 35698
rect 39116 34750 39118 34802
rect 39170 34750 39172 34802
rect 39116 34738 39172 34750
rect 39340 35588 39396 35598
rect 39116 34130 39172 34142
rect 39116 34078 39118 34130
rect 39170 34078 39172 34130
rect 39116 33796 39172 34078
rect 39116 33730 39172 33740
rect 38668 33170 38724 33180
rect 38556 32834 38612 32844
rect 38032 31388 38296 31398
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38032 31322 38296 31332
rect 38032 29820 38296 29830
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38032 29754 38296 29764
rect 38032 28252 38296 28262
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38032 28186 38296 28196
rect 38032 26684 38296 26694
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38032 26618 38296 26628
rect 38032 25116 38296 25126
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38032 25050 38296 25060
rect 38032 23548 38296 23558
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38032 23482 38296 23492
rect 38032 21980 38296 21990
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38032 21914 38296 21924
rect 38032 20412 38296 20422
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38032 20346 38296 20356
rect 39340 20188 39396 35532
rect 39564 35588 39620 35646
rect 39564 35522 39620 35532
rect 40348 35252 40404 35868
rect 40796 35810 40852 35822
rect 40796 35758 40798 35810
rect 40850 35758 40852 35810
rect 40572 35700 40628 35710
rect 40572 35698 40740 35700
rect 40572 35646 40574 35698
rect 40626 35646 40740 35698
rect 40572 35644 40740 35646
rect 40572 35634 40628 35644
rect 40124 35196 40628 35252
rect 40124 34914 40180 35196
rect 40124 34862 40126 34914
rect 40178 34862 40180 34914
rect 40124 34850 40180 34862
rect 39452 34804 39508 34814
rect 39452 34802 39620 34804
rect 39452 34750 39454 34802
rect 39506 34750 39620 34802
rect 39452 34748 39620 34750
rect 39452 34738 39508 34748
rect 39452 34242 39508 34254
rect 39452 34190 39454 34242
rect 39506 34190 39508 34242
rect 39452 27300 39508 34190
rect 39564 34020 39620 34748
rect 40348 34690 40404 34702
rect 40348 34638 40350 34690
rect 40402 34638 40404 34690
rect 39900 34020 39956 34030
rect 39564 34018 39956 34020
rect 39564 33966 39902 34018
rect 39954 33966 39956 34018
rect 39564 33964 39956 33966
rect 39452 27234 39508 27244
rect 39900 22932 39956 33964
rect 40348 32340 40404 34638
rect 40572 34354 40628 35196
rect 40572 34302 40574 34354
rect 40626 34302 40628 34354
rect 40572 34290 40628 34302
rect 40684 33908 40740 35644
rect 40796 35476 40852 35758
rect 40796 35410 40852 35420
rect 40908 34802 40964 36428
rect 41804 35922 41860 36764
rect 41804 35870 41806 35922
rect 41858 35870 41860 35922
rect 40908 34750 40910 34802
rect 40962 34750 40964 34802
rect 40908 34738 40964 34750
rect 41132 35812 41188 35822
rect 40684 33842 40740 33852
rect 40348 32274 40404 32284
rect 41132 28420 41188 35756
rect 41804 35812 41860 35870
rect 41804 35746 41860 35756
rect 42028 35028 42084 35038
rect 42252 35028 42308 39200
rect 43148 36594 43204 39200
rect 43148 36542 43150 36594
rect 43202 36542 43204 36594
rect 43148 36530 43204 36542
rect 42364 36482 42420 36494
rect 42364 36430 42366 36482
rect 42418 36430 42420 36482
rect 42364 35922 42420 36430
rect 43372 36484 43428 36494
rect 43260 36372 43316 36382
rect 42364 35870 42366 35922
rect 42418 35870 42420 35922
rect 42364 35858 42420 35870
rect 42588 35924 42644 35934
rect 42028 35026 42532 35028
rect 42028 34974 42030 35026
rect 42082 34974 42532 35026
rect 42028 34972 42532 34974
rect 42028 34962 42084 34972
rect 42476 34914 42532 34972
rect 42476 34862 42478 34914
rect 42530 34862 42532 34914
rect 42476 34850 42532 34862
rect 41132 28354 41188 28364
rect 41244 34802 41300 34814
rect 41244 34750 41246 34802
rect 41298 34750 41300 34802
rect 41244 34020 41300 34750
rect 42588 34468 42644 35868
rect 43260 35922 43316 36316
rect 43260 35870 43262 35922
rect 43314 35870 43316 35922
rect 43260 35858 43316 35870
rect 42588 34402 42644 34412
rect 42700 35698 42756 35710
rect 42700 35646 42702 35698
rect 42754 35646 42756 35698
rect 41468 34020 41524 34030
rect 41244 34018 41524 34020
rect 41244 33966 41470 34018
rect 41522 33966 41524 34018
rect 41244 33964 41524 33966
rect 39900 22866 39956 22876
rect 41244 21028 41300 33964
rect 41468 33954 41524 33964
rect 41916 34018 41972 34030
rect 41916 33966 41918 34018
rect 41970 33966 41972 34018
rect 41244 20962 41300 20972
rect 41916 33908 41972 33966
rect 42700 34020 42756 35646
rect 43372 35026 43428 36428
rect 43932 35812 43988 35822
rect 43932 35718 43988 35756
rect 43372 34974 43374 35026
rect 43426 34974 43428 35026
rect 43372 34962 43428 34974
rect 43820 35028 43876 35038
rect 44044 35028 44100 39200
rect 44156 36484 44212 36494
rect 44156 36390 44212 36428
rect 44380 35810 44436 35822
rect 44380 35758 44382 35810
rect 44434 35758 44436 35810
rect 44380 35700 44436 35758
rect 44940 35700 44996 39200
rect 45724 36932 45780 36942
rect 45724 36482 45780 36876
rect 45724 36430 45726 36482
rect 45778 36430 45780 36482
rect 45724 36372 45780 36430
rect 45724 36306 45780 36316
rect 45276 36260 45332 36270
rect 45276 36166 45332 36204
rect 44380 35644 44772 35700
rect 44940 35644 45108 35700
rect 44380 35476 44436 35486
rect 44604 35476 44660 35486
rect 43820 35026 44324 35028
rect 43820 34974 43822 35026
rect 43874 34974 44324 35026
rect 43820 34972 44324 34974
rect 43820 34962 43876 34972
rect 44268 34914 44324 34972
rect 44268 34862 44270 34914
rect 44322 34862 44324 34914
rect 44268 34850 44324 34862
rect 42812 34692 42868 34702
rect 42812 34690 43092 34692
rect 42812 34638 42814 34690
rect 42866 34638 43092 34690
rect 42812 34636 43092 34638
rect 42812 34626 42868 34636
rect 42924 34020 42980 34030
rect 42700 34018 42980 34020
rect 42700 33966 42926 34018
rect 42978 33966 42980 34018
rect 42700 33964 42980 33966
rect 39340 20132 39620 20188
rect 38032 18844 38296 18854
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38032 18778 38296 18788
rect 38032 17276 38296 17286
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38032 17210 38296 17220
rect 38032 15708 38296 15718
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38032 15642 38296 15652
rect 38032 14140 38296 14150
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38032 14074 38296 14084
rect 38032 12572 38296 12582
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38032 12506 38296 12516
rect 38032 11004 38296 11014
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38032 10938 38296 10948
rect 38032 9436 38296 9446
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38032 9370 38296 9380
rect 38032 7868 38296 7878
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38032 7802 38296 7812
rect 38892 6580 38948 6590
rect 38032 6300 38296 6310
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38032 6234 38296 6244
rect 38892 6130 38948 6524
rect 38892 6078 38894 6130
rect 38946 6078 38948 6130
rect 38892 6066 38948 6078
rect 39452 6580 39508 6590
rect 39452 6130 39508 6524
rect 39452 6078 39454 6130
rect 39506 6078 39508 6130
rect 39452 5684 39508 6078
rect 39452 5618 39508 5628
rect 38032 4732 38296 4742
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38032 4666 38296 4676
rect 38668 4228 38724 4238
rect 38444 4226 38724 4228
rect 38444 4174 38670 4226
rect 38722 4174 38724 4226
rect 38444 4172 38724 4174
rect 38444 3442 38500 4172
rect 38668 4162 38724 4172
rect 38444 3390 38446 3442
rect 38498 3390 38500 3442
rect 38108 3332 38164 3342
rect 37772 3330 38164 3332
rect 37772 3278 38110 3330
rect 38162 3278 38164 3330
rect 37772 3276 38164 3278
rect 38108 3266 38164 3276
rect 38032 3164 38296 3174
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38032 3098 38296 3108
rect 38444 2548 38500 3390
rect 37996 2492 38500 2548
rect 39340 3442 39396 3454
rect 39340 3390 39342 3442
rect 39394 3390 39396 3442
rect 37996 800 38052 2492
rect 39340 800 39396 3390
rect 39564 3332 39620 20132
rect 41916 8428 41972 33852
rect 42924 19460 42980 33964
rect 43036 32676 43092 34636
rect 43596 34020 43652 34030
rect 43036 32610 43092 32620
rect 43148 33124 43204 33134
rect 43148 31948 43204 33068
rect 43036 31892 43204 31948
rect 43036 20188 43092 31892
rect 43596 27188 43652 33964
rect 44380 31948 44436 35420
rect 44492 35474 44660 35476
rect 44492 35422 44606 35474
rect 44658 35422 44660 35474
rect 44492 35420 44660 35422
rect 44492 34020 44548 35420
rect 44604 35410 44660 35420
rect 44492 33954 44548 33964
rect 44604 34690 44660 34702
rect 44604 34638 44606 34690
rect 44658 34638 44660 34690
rect 44380 31892 44548 31948
rect 44492 28868 44548 31892
rect 44492 28802 44548 28812
rect 43596 27122 43652 27132
rect 44604 26180 44660 34638
rect 44716 34132 44772 35644
rect 44716 33460 44772 34076
rect 44716 33394 44772 33404
rect 44940 35474 44996 35486
rect 44940 35422 44942 35474
rect 44994 35422 44996 35474
rect 44604 26114 44660 26124
rect 43036 20132 43204 20188
rect 42924 19394 42980 19404
rect 41916 8372 42084 8428
rect 41916 6468 41972 6478
rect 41692 6466 41972 6468
rect 41692 6414 41918 6466
rect 41970 6414 41972 6466
rect 41692 6412 41972 6414
rect 39788 6132 39844 6142
rect 39788 5348 39844 6076
rect 39788 5282 39844 5292
rect 41020 5124 41076 5134
rect 41020 5030 41076 5068
rect 41692 5122 41748 6412
rect 41916 6402 41972 6412
rect 41692 5070 41694 5122
rect 41746 5070 41748 5122
rect 41692 5058 41748 5070
rect 40236 4900 40292 4910
rect 40236 3554 40292 4844
rect 40796 4228 40852 4238
rect 40236 3502 40238 3554
rect 40290 3502 40292 3554
rect 40236 3490 40292 3502
rect 40684 4226 40852 4228
rect 40684 4174 40798 4226
rect 40850 4174 40852 4226
rect 40684 4172 40852 4174
rect 40684 3556 40740 4172
rect 40796 4162 40852 4172
rect 39564 3266 39620 3276
rect 40684 800 40740 3500
rect 41244 3556 41300 3566
rect 41244 3462 41300 3500
rect 41020 3332 41076 3342
rect 41020 3238 41076 3276
rect 42028 3330 42084 8372
rect 42252 6580 42308 6590
rect 43036 6580 43092 6590
rect 42252 6578 43092 6580
rect 42252 6526 42254 6578
rect 42306 6526 43038 6578
rect 43090 6526 43092 6578
rect 42252 6524 43092 6526
rect 42252 6514 42308 6524
rect 43036 6514 43092 6524
rect 42588 4226 42644 4238
rect 42588 4174 42590 4226
rect 42642 4174 42644 4226
rect 42028 3278 42030 3330
rect 42082 3278 42084 3330
rect 42028 3266 42084 3278
rect 42252 3556 42308 3566
rect 42588 3556 42644 4174
rect 42252 3554 42644 3556
rect 42252 3502 42254 3554
rect 42306 3502 42644 3554
rect 42252 3500 42644 3502
rect 42252 2548 42308 3500
rect 43148 3220 43204 20132
rect 44268 7586 44324 7598
rect 44268 7534 44270 7586
rect 44322 7534 44324 7586
rect 44156 7364 44212 7374
rect 43372 6916 43428 6926
rect 43372 6822 43428 6860
rect 44156 6690 44212 7308
rect 44156 6638 44158 6690
rect 44210 6638 44212 6690
rect 44156 6626 44212 6638
rect 44044 6578 44100 6590
rect 44044 6526 44046 6578
rect 44098 6526 44100 6578
rect 43820 5908 43876 5918
rect 43820 5814 43876 5852
rect 44044 4900 44100 6526
rect 44268 5906 44324 7534
rect 44604 7474 44660 7486
rect 44604 7422 44606 7474
rect 44658 7422 44660 7474
rect 44604 6692 44660 7422
rect 44940 6916 44996 35422
rect 45052 35140 45108 35644
rect 45612 35588 45668 35598
rect 45612 35494 45668 35532
rect 45052 35074 45108 35084
rect 45724 35140 45780 35150
rect 45724 35026 45780 35084
rect 45724 34974 45726 35026
rect 45778 34974 45780 35026
rect 45724 34962 45780 34974
rect 45836 34130 45892 39200
rect 46732 36708 46788 39200
rect 47628 36932 47684 39200
rect 47628 36866 47684 36876
rect 46732 36642 46788 36652
rect 47628 36708 47684 36718
rect 47516 36482 47572 36494
rect 47516 36430 47518 36482
rect 47570 36430 47572 36482
rect 46844 36370 46900 36382
rect 46844 36318 46846 36370
rect 46898 36318 46900 36370
rect 46060 36258 46116 36270
rect 46060 36206 46062 36258
rect 46114 36206 46116 36258
rect 46060 36036 46116 36206
rect 46060 35970 46116 35980
rect 46396 35812 46452 35822
rect 46396 35718 46452 35756
rect 46172 35698 46228 35710
rect 46172 35646 46174 35698
rect 46226 35646 46228 35698
rect 46172 35588 46228 35646
rect 46060 34244 46116 34254
rect 46060 34150 46116 34188
rect 45836 34078 45838 34130
rect 45890 34078 45892 34130
rect 45276 34020 45332 34030
rect 45276 33926 45332 33964
rect 45836 33460 45892 34078
rect 45836 33394 45892 33404
rect 46172 31948 46228 35532
rect 46620 34914 46676 34926
rect 46620 34862 46622 34914
rect 46674 34862 46676 34914
rect 46620 34354 46676 34862
rect 46620 34302 46622 34354
rect 46674 34302 46676 34354
rect 46620 34290 46676 34302
rect 46844 34692 46900 36318
rect 47180 36370 47236 36382
rect 47180 36318 47182 36370
rect 47234 36318 47236 36370
rect 46956 35812 47012 35822
rect 46956 35698 47012 35756
rect 46956 35646 46958 35698
rect 47010 35646 47012 35698
rect 46956 35634 47012 35646
rect 46284 33460 46340 33470
rect 46284 33366 46340 33404
rect 46844 33458 46900 34636
rect 47068 34356 47124 34366
rect 46956 34130 47012 34142
rect 46956 34078 46958 34130
rect 47010 34078 47012 34130
rect 46956 34020 47012 34078
rect 46956 33954 47012 33964
rect 46844 33406 46846 33458
rect 46898 33406 46900 33458
rect 46844 33394 46900 33406
rect 46060 31892 46228 31948
rect 45276 26964 45332 26974
rect 45164 7364 45220 7374
rect 45164 7270 45220 7308
rect 44604 6626 44660 6636
rect 44828 6692 44884 6702
rect 44940 6692 44996 6860
rect 44828 6690 44996 6692
rect 44828 6638 44830 6690
rect 44882 6638 44996 6690
rect 44828 6636 44996 6638
rect 44828 6626 44884 6636
rect 44268 5854 44270 5906
rect 44322 5854 44324 5906
rect 44268 5842 44324 5854
rect 44044 4834 44100 4844
rect 44156 5236 44212 5246
rect 44156 4898 44212 5180
rect 44156 4846 44158 4898
rect 44210 4846 44212 4898
rect 44156 4834 44212 4846
rect 44716 5122 44772 5134
rect 44716 5070 44718 5122
rect 44770 5070 44772 5122
rect 44716 4900 44772 5070
rect 44716 4834 44772 4844
rect 45052 4340 45108 4350
rect 44716 4226 44772 4238
rect 44716 4174 44718 4226
rect 44770 4174 44772 4226
rect 43148 3154 43204 3164
rect 43372 3666 43428 3678
rect 43372 3614 43374 3666
rect 43426 3614 43428 3666
rect 42028 2492 42308 2548
rect 42028 800 42084 2492
rect 43372 800 43428 3614
rect 44156 3556 44212 3566
rect 44156 3462 44212 3500
rect 44716 3444 44772 4174
rect 45052 4226 45108 4284
rect 45052 4174 45054 4226
rect 45106 4174 45108 4226
rect 45052 3556 45108 4174
rect 45052 3490 45108 3500
rect 44940 3444 44996 3454
rect 44716 3442 44996 3444
rect 44716 3390 44942 3442
rect 44994 3390 44996 3442
rect 44716 3388 44996 3390
rect 44716 800 44772 3388
rect 44940 3378 44996 3388
rect 45276 3330 45332 26908
rect 46060 17668 46116 31892
rect 47068 26964 47124 34300
rect 47180 34132 47236 36318
rect 47516 36260 47572 36430
rect 47516 36194 47572 36204
rect 47628 35586 47684 36652
rect 48524 36596 48580 39200
rect 48524 36530 48580 36540
rect 49308 37268 49364 37278
rect 48972 36482 49028 36494
rect 48972 36430 48974 36482
rect 49026 36430 49028 36482
rect 47852 36260 47908 36270
rect 47852 36258 48020 36260
rect 47852 36206 47854 36258
rect 47906 36206 48020 36258
rect 47852 36204 48020 36206
rect 47852 36194 47908 36204
rect 47628 35534 47630 35586
rect 47682 35534 47684 35586
rect 47628 35522 47684 35534
rect 47740 34802 47796 34814
rect 47740 34750 47742 34802
rect 47794 34750 47796 34802
rect 47292 34690 47348 34702
rect 47292 34638 47294 34690
rect 47346 34638 47348 34690
rect 47292 34356 47348 34638
rect 47292 34290 47348 34300
rect 47740 34356 47796 34750
rect 47740 34290 47796 34300
rect 47180 34066 47236 34076
rect 47404 34020 47460 34030
rect 47404 33926 47460 33964
rect 47964 31948 48020 36204
rect 48748 35588 48804 35598
rect 48636 35586 48804 35588
rect 48636 35534 48750 35586
rect 48802 35534 48804 35586
rect 48636 35532 48804 35534
rect 48636 34802 48692 35532
rect 48748 35522 48804 35532
rect 48636 34750 48638 34802
rect 48690 34750 48692 34802
rect 48076 34692 48132 34702
rect 48076 34598 48132 34636
rect 48524 34244 48580 34254
rect 48188 34132 48244 34142
rect 48188 34038 48244 34076
rect 47068 26898 47124 26908
rect 47852 31892 48020 31948
rect 48412 34020 48468 34030
rect 46060 17602 46116 17612
rect 46172 7364 46228 7374
rect 45948 6916 46004 6926
rect 45948 6822 46004 6860
rect 45612 6692 45668 6702
rect 45612 6598 45668 6636
rect 46172 6578 46228 7308
rect 47180 7364 47236 7374
rect 47180 7270 47236 7308
rect 47852 6916 47908 31892
rect 48412 24500 48468 33964
rect 48524 33236 48580 34188
rect 48524 33170 48580 33180
rect 48412 24434 48468 24444
rect 48636 11284 48692 34750
rect 48972 34802 49028 36430
rect 49308 35588 49364 37212
rect 49420 35812 49476 39200
rect 49532 36596 49588 36606
rect 49532 36502 49588 36540
rect 49420 35756 49700 35812
rect 49420 35588 49476 35598
rect 49308 35586 49476 35588
rect 49308 35534 49422 35586
rect 49474 35534 49476 35586
rect 49308 35532 49476 35534
rect 49420 35522 49476 35532
rect 48972 34750 48974 34802
rect 49026 34750 49028 34802
rect 48972 34738 49028 34750
rect 49196 35252 49252 35262
rect 48860 34356 48916 34366
rect 48860 34262 48916 34300
rect 49196 33458 49252 35196
rect 49532 35252 49588 35262
rect 49532 34914 49588 35196
rect 49532 34862 49534 34914
rect 49586 34862 49588 34914
rect 49532 34850 49588 34862
rect 49644 34356 49700 35756
rect 50316 35810 50372 39200
rect 51212 36036 51268 39200
rect 51324 36596 51380 36606
rect 51324 36502 51380 36540
rect 52108 36596 52164 39200
rect 53004 39060 53060 39200
rect 53228 39060 53284 39228
rect 53004 39004 53284 39060
rect 52892 37268 52948 37278
rect 52108 36530 52164 36540
rect 52668 36708 52724 36718
rect 51996 36482 52052 36494
rect 51996 36430 51998 36482
rect 52050 36430 52052 36482
rect 51996 36148 52052 36430
rect 51996 36082 52052 36092
rect 50316 35758 50318 35810
rect 50370 35758 50372 35810
rect 50316 35746 50372 35758
rect 50652 35980 51268 36036
rect 49980 35140 50036 35150
rect 49644 34242 49700 34300
rect 49644 34190 49646 34242
rect 49698 34190 49700 34242
rect 49644 34178 49700 34190
rect 49868 34690 49924 34702
rect 49868 34638 49870 34690
rect 49922 34638 49924 34690
rect 49196 33406 49198 33458
rect 49250 33406 49252 33458
rect 49196 31948 49252 33406
rect 49196 31892 49364 31948
rect 48636 11218 48692 11228
rect 47852 6692 47908 6860
rect 47964 6692 48020 6702
rect 47852 6690 48020 6692
rect 47852 6638 47966 6690
rect 48018 6638 48020 6690
rect 47852 6636 48020 6638
rect 47964 6626 48020 6636
rect 46172 6526 46174 6578
rect 46226 6526 46228 6578
rect 46172 6514 46228 6526
rect 46508 6578 46564 6590
rect 46508 6526 46510 6578
rect 46562 6526 46564 6578
rect 45948 5572 46004 5582
rect 45388 5124 45444 5134
rect 45388 5030 45444 5068
rect 45948 4228 46004 5516
rect 46508 5572 46564 6526
rect 47516 6466 47572 6478
rect 47516 6414 47518 6466
rect 47570 6414 47572 6466
rect 46732 6132 46788 6142
rect 46732 6130 47124 6132
rect 46732 6078 46734 6130
rect 46786 6078 47124 6130
rect 46732 6076 47124 6078
rect 46732 6066 46788 6076
rect 46508 5506 46564 5516
rect 47068 5346 47124 6076
rect 47292 5684 47348 5694
rect 47516 5684 47572 6414
rect 47628 5908 47684 5918
rect 47628 5814 47684 5852
rect 47292 5682 47572 5684
rect 47292 5630 47294 5682
rect 47346 5630 47572 5682
rect 47292 5628 47572 5630
rect 47740 5796 47796 5806
rect 47292 5572 47348 5628
rect 47292 5506 47348 5516
rect 47068 5294 47070 5346
rect 47122 5294 47124 5346
rect 47068 5282 47124 5294
rect 46396 5236 46452 5246
rect 46620 5236 46676 5246
rect 46396 5142 46452 5180
rect 46508 5180 46620 5236
rect 46508 5122 46564 5180
rect 46508 5070 46510 5122
rect 46562 5070 46564 5122
rect 46508 5058 46564 5070
rect 46620 4564 46676 5180
rect 47180 5236 47236 5246
rect 47628 5236 47684 5246
rect 47740 5236 47796 5740
rect 47236 5234 47796 5236
rect 47236 5182 47630 5234
rect 47682 5182 47796 5234
rect 47236 5180 47796 5182
rect 47180 5104 47236 5180
rect 47628 5170 47684 5180
rect 46732 4564 46788 4574
rect 46620 4562 46788 4564
rect 46620 4510 46734 4562
rect 46786 4510 46788 4562
rect 46620 4508 46788 4510
rect 46732 4498 46788 4508
rect 48188 4564 48244 4574
rect 45948 4162 46004 4172
rect 46172 4228 46228 4238
rect 46172 3556 46228 4172
rect 47180 4228 47236 4238
rect 47180 4134 47236 4172
rect 46060 3554 46228 3556
rect 46060 3502 46174 3554
rect 46226 3502 46228 3554
rect 46060 3500 46228 3502
rect 45276 3278 45278 3330
rect 45330 3278 45332 3330
rect 45276 3266 45332 3278
rect 45948 3332 46004 3342
rect 45948 3238 46004 3276
rect 46060 800 46116 3500
rect 46172 3490 46228 3500
rect 47404 3666 47460 3678
rect 47404 3614 47406 3666
rect 47458 3614 47460 3666
rect 47404 800 47460 3614
rect 48076 3556 48132 3566
rect 48188 3556 48244 4508
rect 48076 3554 48244 3556
rect 48076 3502 48078 3554
rect 48130 3502 48244 3554
rect 48076 3500 48244 3502
rect 48748 4226 48804 4238
rect 48748 4174 48750 4226
rect 48802 4174 48804 4226
rect 48076 3490 48132 3500
rect 48748 3444 48804 4174
rect 48972 3444 49028 3454
rect 48748 3442 49028 3444
rect 48748 3390 48974 3442
rect 49026 3390 49028 3442
rect 48748 3388 49028 3390
rect 48748 800 48804 3388
rect 48972 3378 49028 3388
rect 49308 3330 49364 31892
rect 49868 28084 49924 34638
rect 49980 34354 50036 35084
rect 50652 34916 50708 35980
rect 51884 35812 51940 35822
rect 51548 35810 51940 35812
rect 51548 35758 51886 35810
rect 51938 35758 51940 35810
rect 51548 35756 51940 35758
rect 51212 35700 51268 35710
rect 51212 35698 51492 35700
rect 51212 35646 51214 35698
rect 51266 35646 51492 35698
rect 51212 35644 51492 35646
rect 51212 35634 51268 35644
rect 50652 34914 50820 34916
rect 50652 34862 50654 34914
rect 50706 34862 50820 34914
rect 50652 34860 50820 34862
rect 50652 34850 50708 34860
rect 49980 34302 49982 34354
rect 50034 34302 50036 34354
rect 49980 34290 50036 34302
rect 50316 34692 50372 34702
rect 49868 28018 49924 28028
rect 50316 26292 50372 34636
rect 50764 34356 50820 34860
rect 51436 34802 51492 35644
rect 51436 34750 51438 34802
rect 51490 34750 51492 34802
rect 51436 34738 51492 34750
rect 50876 34692 50932 34702
rect 50876 34690 51044 34692
rect 50876 34638 50878 34690
rect 50930 34638 51044 34690
rect 50876 34636 51044 34638
rect 50876 34626 50932 34636
rect 50876 34356 50932 34366
rect 50764 34354 50932 34356
rect 50764 34302 50878 34354
rect 50930 34302 50932 34354
rect 50764 34300 50932 34302
rect 50876 34290 50932 34300
rect 50988 34356 51044 34636
rect 50988 34290 51044 34300
rect 51212 34020 51268 34030
rect 50316 26226 50372 26236
rect 50652 33572 50708 33582
rect 49308 3278 49310 3330
rect 49362 3278 49364 3330
rect 49308 3266 49364 3278
rect 49532 26068 49588 26078
rect 49532 3332 49588 26012
rect 50540 6468 50596 6478
rect 50540 5684 50596 6412
rect 50540 5618 50596 5628
rect 49868 3444 49924 3454
rect 50316 3444 50372 3454
rect 49868 3442 50372 3444
rect 49868 3390 49870 3442
rect 49922 3390 50318 3442
rect 50370 3390 50372 3442
rect 49868 3388 50372 3390
rect 49868 3378 49924 3388
rect 49532 3266 49588 3276
rect 50092 800 50148 3388
rect 50316 3378 50372 3388
rect 50652 3330 50708 33516
rect 51212 33572 51268 33964
rect 51212 33506 51268 33516
rect 51548 33348 51604 35756
rect 51884 35746 51940 35756
rect 52444 35810 52500 35822
rect 52444 35758 52446 35810
rect 52498 35758 52500 35810
rect 52444 35476 52500 35758
rect 52668 35698 52724 36652
rect 52892 36370 52948 37212
rect 52892 36318 52894 36370
rect 52946 36318 52948 36370
rect 52892 36306 52948 36318
rect 53004 36482 53060 36494
rect 53004 36430 53006 36482
rect 53058 36430 53060 36482
rect 53004 35700 53060 36430
rect 52668 35646 52670 35698
rect 52722 35646 52724 35698
rect 52668 35634 52724 35646
rect 52892 35644 53060 35700
rect 53564 35812 53620 39228
rect 53872 39200 53984 40000
rect 54236 39228 54628 39284
rect 53900 39060 53956 39200
rect 54236 39060 54292 39228
rect 53900 39004 54292 39060
rect 54572 37604 54628 39228
rect 54768 39200 54880 40000
rect 55664 39200 55776 40000
rect 56560 39200 56672 40000
rect 57456 39200 57568 40000
rect 58352 39200 58464 40000
rect 59248 39200 59360 40000
rect 60144 39200 60256 40000
rect 61040 39200 61152 40000
rect 61936 39200 62048 40000
rect 62832 39200 62944 40000
rect 63728 39200 63840 40000
rect 64624 39200 64736 40000
rect 65520 39200 65632 40000
rect 66416 39200 66528 40000
rect 67312 39200 67424 40000
rect 68208 39200 68320 40000
rect 69104 39200 69216 40000
rect 70000 39200 70112 40000
rect 70896 39200 71008 40000
rect 71792 39200 71904 40000
rect 72688 39200 72800 40000
rect 73584 39200 73696 40000
rect 74480 39200 74592 40000
rect 75376 39200 75488 40000
rect 76272 39200 76384 40000
rect 77168 39200 77280 40000
rect 78064 39200 78176 40000
rect 78960 39200 79072 40000
rect 79856 39200 79968 40000
rect 80752 39200 80864 40000
rect 81648 39200 81760 40000
rect 82544 39200 82656 40000
rect 83440 39200 83552 40000
rect 84336 39200 84448 40000
rect 84700 39228 85092 39284
rect 54796 38052 54852 39200
rect 54796 37996 55076 38052
rect 54572 37548 54964 37604
rect 53900 36708 53956 36718
rect 53676 36484 53732 36494
rect 53676 36482 53844 36484
rect 53676 36430 53678 36482
rect 53730 36430 53844 36482
rect 53676 36428 53844 36430
rect 53676 36418 53732 36428
rect 53788 35924 53844 36428
rect 53788 35858 53844 35868
rect 53676 35812 53732 35822
rect 53564 35810 53732 35812
rect 53564 35758 53678 35810
rect 53730 35758 53732 35810
rect 53564 35756 53732 35758
rect 52892 35476 52948 35644
rect 52444 35420 52948 35476
rect 53004 35476 53060 35486
rect 51548 33254 51604 33292
rect 51660 35364 51716 35374
rect 51660 34354 51716 35308
rect 51660 34302 51662 34354
rect 51714 34302 51716 34354
rect 51660 34244 51716 34302
rect 51660 26068 51716 34188
rect 51772 34802 51828 34814
rect 51772 34750 51774 34802
rect 51826 34750 51828 34802
rect 51772 33460 51828 34750
rect 52332 34802 52388 34814
rect 52332 34750 52334 34802
rect 52386 34750 52388 34802
rect 52220 34468 52276 34478
rect 52220 34354 52276 34412
rect 52220 34302 52222 34354
rect 52274 34302 52276 34354
rect 52220 34290 52276 34302
rect 52332 34020 52388 34750
rect 52332 33954 52388 33964
rect 51996 33460 52052 33470
rect 51772 33458 52052 33460
rect 51772 33406 51998 33458
rect 52050 33406 52052 33458
rect 51772 33404 52052 33406
rect 51996 30212 52052 33404
rect 52444 33348 52500 35420
rect 53004 35382 53060 35420
rect 53452 35028 53508 35038
rect 52556 35026 53508 35028
rect 52556 34974 53454 35026
rect 53506 34974 53508 35026
rect 52556 34972 53508 34974
rect 52556 34242 52612 34972
rect 53452 34962 53508 34972
rect 52556 34190 52558 34242
rect 52610 34190 52612 34242
rect 52556 34178 52612 34190
rect 52668 34690 52724 34702
rect 52668 34638 52670 34690
rect 52722 34638 52724 34690
rect 52444 33282 52500 33292
rect 52668 31948 52724 34638
rect 53116 34244 53172 34254
rect 53116 34150 53172 34188
rect 53452 34244 53508 34254
rect 53452 34150 53508 34188
rect 53340 33460 53396 33470
rect 52780 33348 52836 33358
rect 52780 33254 52836 33292
rect 51996 30146 52052 30156
rect 52444 31892 52724 31948
rect 52444 29652 52500 31892
rect 53340 31108 53396 33404
rect 53452 32788 53508 32798
rect 53564 32788 53620 35756
rect 53676 35746 53732 35756
rect 53788 35588 53844 35598
rect 53452 32786 53620 32788
rect 53452 32734 53454 32786
rect 53506 32734 53620 32786
rect 53452 32732 53620 32734
rect 53676 35476 53732 35486
rect 53452 32722 53508 32732
rect 53340 31042 53396 31052
rect 52444 29586 52500 29596
rect 51660 26002 51716 26012
rect 53004 14308 53060 14318
rect 51660 7364 51716 7374
rect 50988 6468 51044 6478
rect 50988 6374 51044 6412
rect 51324 6466 51380 6478
rect 51324 6414 51326 6466
rect 51378 6414 51380 6466
rect 51324 6356 51380 6414
rect 51324 6290 51380 6300
rect 51436 4228 51492 4238
rect 51212 3444 51268 3454
rect 51212 3350 51268 3388
rect 50652 3278 50654 3330
rect 50706 3278 50708 3330
rect 50652 3266 50708 3278
rect 51436 800 51492 4172
rect 51660 3330 51716 7308
rect 52556 7252 52612 7262
rect 52556 5236 52612 7196
rect 52668 6466 52724 6478
rect 52668 6414 52670 6466
rect 52722 6414 52724 6466
rect 52668 6356 52724 6414
rect 52668 6290 52724 6300
rect 52892 6020 52948 6030
rect 52668 5236 52724 5246
rect 52556 5234 52724 5236
rect 52556 5182 52670 5234
rect 52722 5182 52724 5234
rect 52556 5180 52724 5182
rect 52668 5170 52724 5180
rect 52332 5122 52388 5134
rect 52332 5070 52334 5122
rect 52386 5070 52388 5122
rect 51884 4228 51940 4238
rect 51884 4134 51940 4172
rect 51996 3556 52052 3566
rect 51996 3462 52052 3500
rect 52332 3556 52388 5070
rect 52892 4338 52948 5964
rect 52892 4286 52894 4338
rect 52946 4286 52948 4338
rect 52892 4274 52948 4286
rect 52332 3490 52388 3500
rect 52780 3556 52836 3566
rect 51660 3278 51662 3330
rect 51714 3278 51716 3330
rect 51660 3266 51716 3278
rect 52780 800 52836 3500
rect 53004 3330 53060 14252
rect 53452 7252 53508 7262
rect 53452 6690 53508 7196
rect 53452 6638 53454 6690
rect 53506 6638 53508 6690
rect 53452 6132 53508 6638
rect 53564 6132 53620 6142
rect 53452 6130 53620 6132
rect 53452 6078 53566 6130
rect 53618 6078 53620 6130
rect 53452 6076 53620 6078
rect 53564 6066 53620 6076
rect 53116 6020 53172 6030
rect 53116 5926 53172 5964
rect 53676 5236 53732 35420
rect 53788 35138 53844 35532
rect 53788 35086 53790 35138
rect 53842 35086 53844 35138
rect 53788 35074 53844 35086
rect 53900 33458 53956 36652
rect 54908 36594 54964 37548
rect 54908 36542 54910 36594
rect 54962 36542 54964 36594
rect 54908 36530 54964 36542
rect 54012 36260 54068 36270
rect 54012 36258 54516 36260
rect 54012 36206 54014 36258
rect 54066 36206 54516 36258
rect 54012 36204 54516 36206
rect 54012 36194 54068 36204
rect 54012 35812 54068 35822
rect 54012 35810 54404 35812
rect 54012 35758 54014 35810
rect 54066 35758 54404 35810
rect 54012 35756 54404 35758
rect 54012 35746 54068 35756
rect 54236 35588 54292 35598
rect 53900 33406 53902 33458
rect 53954 33406 53956 33458
rect 53900 33394 53956 33406
rect 54012 34802 54068 34814
rect 54012 34750 54014 34802
rect 54066 34750 54068 34802
rect 54012 34580 54068 34750
rect 54012 33460 54068 34524
rect 54236 34354 54292 35532
rect 54236 34302 54238 34354
rect 54290 34302 54292 34354
rect 54236 34290 54292 34302
rect 54012 33394 54068 33404
rect 54348 31108 54404 35756
rect 54460 33684 54516 36204
rect 54572 36148 54628 36158
rect 54572 35922 54628 36092
rect 54572 35870 54574 35922
rect 54626 35870 54628 35922
rect 54572 35858 54628 35870
rect 54796 35924 54852 35934
rect 54796 35140 54852 35868
rect 54908 35700 54964 35710
rect 54908 35606 54964 35644
rect 54796 35084 54964 35140
rect 54572 34916 54628 34926
rect 54572 34822 54628 34860
rect 54796 34356 54852 34366
rect 54908 34356 54964 35084
rect 55020 34916 55076 37996
rect 55692 37380 55748 39200
rect 55692 37324 55860 37380
rect 55804 35810 55860 37324
rect 56588 37044 56644 39200
rect 56028 36988 56644 37044
rect 56924 38276 56980 38286
rect 55804 35758 55806 35810
rect 55858 35758 55860 35810
rect 55804 35746 55860 35758
rect 55916 36482 55972 36494
rect 55916 36430 55918 36482
rect 55970 36430 55972 36482
rect 55020 34784 55076 34860
rect 55244 35700 55300 35710
rect 54796 34354 54964 34356
rect 54796 34302 54798 34354
rect 54850 34302 54964 34354
rect 54796 34300 54964 34302
rect 54796 34290 54852 34300
rect 55132 34020 55188 34030
rect 55244 34020 55300 35644
rect 55132 34018 55300 34020
rect 55132 33966 55134 34018
rect 55186 33966 55300 34018
rect 55132 33964 55300 33966
rect 55132 33954 55188 33964
rect 54460 33628 54964 33684
rect 54460 33348 54516 33358
rect 54460 33254 54516 33292
rect 54348 31042 54404 31052
rect 54908 20188 54964 33628
rect 54908 20132 55188 20188
rect 54572 7252 54628 7262
rect 54012 6466 54068 6478
rect 54012 6414 54014 6466
rect 54066 6414 54068 6466
rect 54012 6356 54068 6414
rect 54012 6290 54068 6300
rect 53676 5104 53732 5180
rect 54460 5236 54516 5246
rect 54348 5012 54404 5022
rect 54124 5010 54404 5012
rect 54124 4958 54350 5010
rect 54402 4958 54404 5010
rect 54124 4956 54404 4958
rect 54124 4562 54180 4956
rect 54348 4946 54404 4956
rect 54124 4510 54126 4562
rect 54178 4510 54180 4562
rect 54124 4498 54180 4510
rect 53452 4340 53508 4350
rect 53452 4246 53508 4284
rect 54012 4340 54068 4350
rect 54012 3668 54068 4284
rect 54460 4338 54516 5180
rect 54460 4286 54462 4338
rect 54514 4286 54516 4338
rect 54460 4274 54516 4286
rect 54572 4452 54628 7196
rect 55132 6132 55188 20132
rect 55244 19348 55300 33964
rect 55356 34690 55412 34702
rect 55356 34638 55358 34690
rect 55410 34638 55412 34690
rect 55356 29988 55412 34638
rect 55804 34020 55860 34030
rect 55916 34020 55972 36430
rect 56028 35026 56084 36988
rect 56442 36876 56706 36886
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56442 36810 56706 36820
rect 56812 36370 56868 36382
rect 56812 36318 56814 36370
rect 56866 36318 56868 36370
rect 56700 35700 56756 35710
rect 56700 35606 56756 35644
rect 56442 35308 56706 35318
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56442 35242 56706 35252
rect 56028 34974 56030 35026
rect 56082 34974 56084 35026
rect 56028 34916 56084 34974
rect 56812 34916 56868 36318
rect 56028 34850 56084 34860
rect 56588 34860 56868 34916
rect 56476 34804 56532 34814
rect 55804 34018 55972 34020
rect 55804 33966 55806 34018
rect 55858 33966 55972 34018
rect 55804 33964 55972 33966
rect 56028 34244 56084 34254
rect 55804 33572 55860 33964
rect 55804 33506 55860 33516
rect 56028 31220 56084 34188
rect 56140 34020 56196 34030
rect 56140 33926 56196 33964
rect 56476 34020 56532 34748
rect 56476 33954 56532 33964
rect 56588 34354 56644 34860
rect 56812 34692 56868 34702
rect 56924 34692 56980 38220
rect 57148 38052 57204 38062
rect 57148 36370 57204 37996
rect 57484 37828 57540 39200
rect 57484 37772 57988 37828
rect 57932 36594 57988 37772
rect 57932 36542 57934 36594
rect 57986 36542 57988 36594
rect 57932 36530 57988 36542
rect 57148 36318 57150 36370
rect 57202 36318 57204 36370
rect 57148 36306 57204 36318
rect 57596 36484 57652 36494
rect 57596 35922 57652 36428
rect 57596 35870 57598 35922
rect 57650 35870 57652 35922
rect 57596 35858 57652 35870
rect 57484 35700 57540 35710
rect 57372 34916 57428 34926
rect 57372 34822 57428 34860
rect 56812 34690 56980 34692
rect 56812 34638 56814 34690
rect 56866 34638 56980 34690
rect 56812 34636 56980 34638
rect 56812 34626 56868 34636
rect 56588 34302 56590 34354
rect 56642 34302 56644 34354
rect 56588 33908 56644 34302
rect 56588 33842 56644 33852
rect 57484 34354 57540 35644
rect 57820 35698 57876 35710
rect 57820 35646 57822 35698
rect 57874 35646 57876 35698
rect 57484 34302 57486 34354
rect 57538 34302 57540 34354
rect 56442 33740 56706 33750
rect 56028 31154 56084 31164
rect 56252 33684 56308 33694
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56442 33674 56706 33684
rect 55356 29922 55412 29932
rect 55244 19282 55300 19292
rect 56252 7364 56308 33628
rect 56442 32172 56706 32182
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56442 32106 56706 32116
rect 56442 30604 56706 30614
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56442 30538 56706 30548
rect 57484 29540 57540 34302
rect 57708 34690 57764 34702
rect 57708 34638 57710 34690
rect 57762 34638 57764 34690
rect 57708 31556 57764 34638
rect 57708 31490 57764 31500
rect 57820 34018 57876 35646
rect 58380 34916 58436 39200
rect 58940 38612 58996 38622
rect 58828 36484 58884 36494
rect 58828 36390 58884 36428
rect 58716 36260 58772 36270
rect 58604 35812 58660 35822
rect 58604 35718 58660 35756
rect 58604 34916 58660 34926
rect 58380 34914 58660 34916
rect 58380 34862 58606 34914
rect 58658 34862 58660 34914
rect 58380 34860 58660 34862
rect 58380 34354 58436 34860
rect 58604 34850 58660 34860
rect 58380 34302 58382 34354
rect 58434 34302 58436 34354
rect 58380 34290 58436 34302
rect 57820 33966 57822 34018
rect 57874 33966 57876 34018
rect 57484 29474 57540 29484
rect 56442 29036 56706 29046
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56442 28970 56706 28980
rect 56442 27468 56706 27478
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56442 27402 56706 27412
rect 56442 25900 56706 25910
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56442 25834 56706 25844
rect 56442 24332 56706 24342
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56442 24266 56706 24276
rect 56442 22764 56706 22774
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56442 22698 56706 22708
rect 56442 21196 56706 21206
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56442 21130 56706 21140
rect 56442 19628 56706 19638
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56442 19562 56706 19572
rect 56442 18060 56706 18070
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56442 17994 56706 18004
rect 56442 16492 56706 16502
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56442 16426 56706 16436
rect 56442 14924 56706 14934
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56442 14858 56706 14868
rect 56442 13356 56706 13366
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56442 13290 56706 13300
rect 57820 12740 57876 33966
rect 58716 34018 58772 36204
rect 58940 35922 58996 38556
rect 59276 37604 59332 39200
rect 59276 37548 59780 37604
rect 59612 37380 59668 37390
rect 58940 35870 58942 35922
rect 58994 35870 58996 35922
rect 58940 35858 58996 35870
rect 59164 36484 59220 36494
rect 58716 33966 58718 34018
rect 58770 33966 58772 34018
rect 58716 32788 58772 33966
rect 58716 32722 58772 32732
rect 58940 34690 58996 34702
rect 58940 34638 58942 34690
rect 58994 34638 58996 34690
rect 58156 30212 58212 30222
rect 58156 20188 58212 30156
rect 58940 30100 58996 34638
rect 58940 30034 58996 30044
rect 59052 34020 59108 34030
rect 58156 20132 58436 20188
rect 57820 12674 57876 12684
rect 56442 11788 56706 11798
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56442 11722 56706 11732
rect 56442 10220 56706 10230
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56442 10154 56706 10164
rect 56442 8652 56706 8662
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56442 8586 56706 8596
rect 58156 8148 58212 8158
rect 56252 7298 56308 7308
rect 57708 7588 57764 7598
rect 56442 7084 56706 7094
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56442 7018 56706 7028
rect 57148 6690 57204 6702
rect 57148 6638 57150 6690
rect 57202 6638 57204 6690
rect 54796 6130 55188 6132
rect 54796 6078 55134 6130
rect 55186 6078 55188 6130
rect 54796 6076 55188 6078
rect 54684 5236 54740 5246
rect 54684 5010 54740 5180
rect 54684 4958 54686 5010
rect 54738 4958 54740 5010
rect 54684 4946 54740 4958
rect 54684 4452 54740 4462
rect 54572 4450 54740 4452
rect 54572 4398 54686 4450
rect 54738 4398 54740 4450
rect 54572 4396 54740 4398
rect 53788 3556 53844 3566
rect 53340 3444 53396 3454
rect 53340 3350 53396 3388
rect 53004 3278 53006 3330
rect 53058 3278 53060 3330
rect 53004 3266 53060 3278
rect 53788 2996 53844 3500
rect 54012 3442 54068 3612
rect 54012 3390 54014 3442
rect 54066 3390 54068 3442
rect 54012 3378 54068 3390
rect 54124 3444 54180 3454
rect 53788 2930 53844 2940
rect 54124 800 54180 3388
rect 54572 3442 54628 4396
rect 54684 4386 54740 4396
rect 54796 3778 54852 6076
rect 55132 6066 55188 6076
rect 55244 6132 55300 6142
rect 55244 4564 55300 6076
rect 55692 6132 55748 6142
rect 55356 5908 55412 5918
rect 55356 5122 55412 5852
rect 55692 5794 55748 6076
rect 57148 5908 57204 6638
rect 57708 6690 57764 7532
rect 58156 7364 58212 8092
rect 57708 6638 57710 6690
rect 57762 6638 57764 6690
rect 57708 6626 57764 6638
rect 58044 7362 58212 7364
rect 58044 7310 58158 7362
rect 58210 7310 58212 7362
rect 58044 7308 58212 7310
rect 57148 5842 57204 5852
rect 57820 5908 57876 5918
rect 57820 5814 57876 5852
rect 55692 5742 55694 5794
rect 55746 5742 55748 5794
rect 55692 5684 55748 5742
rect 55692 5618 55748 5628
rect 56364 5794 56420 5806
rect 56364 5742 56366 5794
rect 56418 5742 56420 5794
rect 56364 5682 56420 5742
rect 56364 5630 56366 5682
rect 56418 5630 56420 5682
rect 56364 5618 56420 5630
rect 56812 5794 56868 5806
rect 56812 5742 56814 5794
rect 56866 5742 56868 5794
rect 56442 5516 56706 5526
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56442 5450 56706 5460
rect 55356 5070 55358 5122
rect 55410 5070 55412 5122
rect 55356 5058 55412 5070
rect 55692 5236 55748 5246
rect 55692 5122 55748 5180
rect 55692 5070 55694 5122
rect 55746 5070 55748 5122
rect 55692 5058 55748 5070
rect 56812 4564 56868 5742
rect 57484 5794 57540 5806
rect 57484 5742 57486 5794
rect 57538 5742 57540 5794
rect 55244 4450 55300 4508
rect 56588 4508 56812 4564
rect 55244 4398 55246 4450
rect 55298 4398 55300 4450
rect 55244 4386 55300 4398
rect 56364 4450 56420 4462
rect 56364 4398 56366 4450
rect 56418 4398 56420 4450
rect 55916 4226 55972 4238
rect 55916 4174 55918 4226
rect 55970 4174 55972 4226
rect 54796 3726 54798 3778
rect 54850 3726 54852 3778
rect 54796 3714 54852 3726
rect 55132 3780 55188 3790
rect 55132 3686 55188 3724
rect 55916 3556 55972 4174
rect 56364 4116 56420 4398
rect 56588 4116 56644 4508
rect 56812 4498 56868 4508
rect 56924 5682 56980 5694
rect 56924 5630 56926 5682
rect 56978 5630 56980 5682
rect 56700 4340 56756 4350
rect 56924 4340 56980 5630
rect 57484 5012 57540 5742
rect 57484 4946 57540 4956
rect 57932 5460 57988 5470
rect 57932 4562 57988 5404
rect 57932 4510 57934 4562
rect 57986 4510 57988 4562
rect 57932 4498 57988 4510
rect 56700 4338 56980 4340
rect 56700 4286 56702 4338
rect 56754 4286 56980 4338
rect 56700 4284 56980 4286
rect 56700 4274 56756 4284
rect 56588 4060 56868 4116
rect 56364 4050 56420 4060
rect 56442 3948 56706 3958
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56442 3882 56706 3892
rect 55916 3462 55972 3500
rect 54572 3390 54574 3442
rect 54626 3390 54628 3442
rect 54572 3378 54628 3390
rect 55468 3444 55524 3454
rect 55468 800 55524 3388
rect 56812 800 56868 4060
rect 56924 2996 56980 4284
rect 57596 4338 57652 4350
rect 57596 4286 57598 4338
rect 57650 4286 57652 4338
rect 57596 3780 57652 4286
rect 57596 3714 57652 3724
rect 57932 3556 57988 3566
rect 58044 3556 58100 7308
rect 58156 7298 58212 7308
rect 58268 5796 58324 5806
rect 58268 5702 58324 5740
rect 58268 5236 58324 5246
rect 57932 3554 58100 3556
rect 57932 3502 57934 3554
rect 57986 3502 58100 3554
rect 57932 3500 58100 3502
rect 58156 5012 58212 5022
rect 57932 3490 57988 3500
rect 57036 3444 57092 3454
rect 57036 3350 57092 3388
rect 56924 2930 56980 2940
rect 58156 800 58212 4956
rect 58268 4898 58324 5180
rect 58268 4846 58270 4898
rect 58322 4846 58324 4898
rect 58268 4834 58324 4846
rect 58380 2660 58436 20132
rect 59052 14308 59108 33964
rect 59164 33460 59220 36428
rect 59500 36370 59556 36382
rect 59500 36318 59502 36370
rect 59554 36318 59556 36370
rect 59500 36260 59556 36318
rect 59500 36194 59556 36204
rect 59276 35812 59332 35822
rect 59276 34354 59332 35756
rect 59612 35026 59668 37324
rect 59724 35586 59780 37548
rect 59836 36260 59892 36270
rect 59836 36258 60004 36260
rect 59836 36206 59838 36258
rect 59890 36206 60004 36258
rect 59836 36204 60004 36206
rect 59836 36194 59892 36204
rect 59724 35534 59726 35586
rect 59778 35534 59780 35586
rect 59724 35522 59780 35534
rect 59612 34974 59614 35026
rect 59666 34974 59668 35026
rect 59612 34916 59668 34974
rect 59612 34850 59668 34860
rect 59276 34302 59278 34354
rect 59330 34302 59332 34354
rect 59276 34290 59332 34302
rect 59836 34020 59892 34030
rect 59836 33926 59892 33964
rect 59276 33460 59332 33470
rect 59164 33458 59332 33460
rect 59164 33406 59278 33458
rect 59330 33406 59332 33458
rect 59164 33404 59332 33406
rect 59276 33394 59332 33404
rect 59948 27860 60004 36204
rect 60172 35812 60228 39200
rect 60172 35746 60228 35756
rect 60732 37716 60788 37726
rect 60732 35698 60788 37660
rect 61068 36594 61124 39200
rect 61404 37940 61460 37950
rect 61068 36542 61070 36594
rect 61122 36542 61124 36594
rect 61068 36530 61124 36542
rect 61292 36820 61348 36830
rect 60732 35646 60734 35698
rect 60786 35646 60788 35698
rect 60060 34802 60116 34814
rect 60060 34750 60062 34802
rect 60114 34750 60116 34802
rect 60060 34132 60116 34750
rect 60060 34066 60116 34076
rect 60620 34690 60676 34702
rect 60620 34638 60622 34690
rect 60674 34638 60676 34690
rect 60620 34132 60676 34638
rect 60172 34020 60228 34030
rect 60620 34020 60676 34076
rect 60228 34018 60676 34020
rect 60228 33966 60622 34018
rect 60674 33966 60676 34018
rect 60228 33964 60676 33966
rect 60172 33888 60228 33964
rect 60284 33460 60340 33470
rect 60284 33366 60340 33404
rect 60620 33124 60676 33964
rect 60732 33460 60788 35646
rect 61292 35922 61348 36764
rect 61404 36484 61460 37884
rect 61404 36418 61460 36428
rect 61740 36482 61796 36494
rect 61740 36430 61742 36482
rect 61794 36430 61796 36482
rect 61292 35870 61294 35922
rect 61346 35870 61348 35922
rect 61292 35588 61348 35870
rect 61292 35522 61348 35532
rect 61516 35698 61572 35710
rect 61516 35646 61518 35698
rect 61570 35646 61572 35698
rect 61516 34692 61572 35646
rect 61180 34636 61572 34692
rect 61628 34690 61684 34702
rect 61628 34638 61630 34690
rect 61682 34638 61684 34690
rect 61180 34132 61236 34636
rect 61628 34580 61684 34638
rect 61180 34038 61236 34076
rect 61292 34524 61684 34580
rect 60732 33394 60788 33404
rect 61292 33348 61348 34524
rect 61740 34244 61796 36430
rect 61628 34188 61796 34244
rect 61292 33282 61348 33292
rect 61404 33684 61460 33694
rect 60396 33122 60676 33124
rect 60396 33070 60622 33122
rect 60674 33070 60676 33122
rect 60396 33068 60676 33070
rect 59948 27794 60004 27804
rect 60284 32452 60340 32462
rect 60284 26852 60340 32396
rect 60284 26786 60340 26796
rect 59052 14242 59108 14252
rect 60284 14308 60340 14318
rect 59052 11620 59108 11630
rect 58716 7362 58772 7374
rect 58716 7310 58718 7362
rect 58770 7310 58772 7362
rect 58492 4564 58548 4574
rect 58492 4450 58548 4508
rect 58492 4398 58494 4450
rect 58546 4398 58548 4450
rect 58492 4386 58548 4398
rect 58716 3668 58772 7310
rect 59052 5908 59108 11564
rect 60284 11620 60340 14252
rect 60284 11554 60340 11564
rect 59612 9268 59668 9278
rect 59164 7588 59220 7598
rect 59164 7494 59220 7532
rect 59500 7476 59556 7486
rect 59500 7382 59556 7420
rect 59052 5852 59220 5908
rect 58828 5796 58884 5806
rect 58828 5794 59108 5796
rect 58828 5742 58830 5794
rect 58882 5742 59108 5794
rect 58828 5740 59108 5742
rect 58828 5730 58884 5740
rect 58828 5572 58884 5582
rect 58828 5346 58884 5516
rect 58828 5294 58830 5346
rect 58882 5294 58884 5346
rect 58828 5282 58884 5294
rect 59052 4900 59108 5740
rect 59052 4834 59108 4844
rect 59164 4676 59220 5852
rect 59388 5796 59444 5806
rect 59388 5702 59444 5740
rect 59276 5682 59332 5694
rect 59276 5630 59278 5682
rect 59330 5630 59332 5682
rect 59276 5236 59332 5630
rect 59276 5170 59332 5180
rect 59276 5012 59332 5022
rect 59276 4918 59332 4956
rect 59612 4898 59668 9212
rect 60396 8428 60452 33068
rect 60620 33058 60676 33068
rect 61404 20188 61460 33628
rect 61628 32788 61684 34188
rect 61740 34020 61796 34030
rect 61740 34018 61908 34020
rect 61740 33966 61742 34018
rect 61794 33966 61908 34018
rect 61740 33964 61908 33966
rect 61740 33954 61796 33964
rect 61740 33460 61796 33470
rect 61740 33366 61796 33404
rect 61628 32722 61684 32732
rect 61852 32452 61908 33964
rect 61964 33460 62020 39200
rect 62636 37380 62692 37390
rect 62524 37044 62580 37054
rect 62524 36372 62580 36988
rect 62300 36370 62580 36372
rect 62300 36318 62526 36370
rect 62578 36318 62580 36370
rect 62300 36316 62580 36318
rect 62188 34916 62244 34926
rect 62188 34822 62244 34860
rect 62300 34356 62356 36316
rect 62524 36306 62580 36316
rect 62188 34300 62356 34356
rect 62412 35810 62468 35822
rect 62412 35758 62414 35810
rect 62466 35758 62468 35810
rect 62188 33572 62244 34300
rect 62300 34132 62356 34142
rect 62300 34038 62356 34076
rect 62188 33516 62356 33572
rect 62020 33404 62244 33460
rect 61964 33394 62020 33404
rect 62188 33346 62244 33404
rect 62188 33294 62190 33346
rect 62242 33294 62244 33346
rect 62188 33282 62244 33294
rect 61852 32386 61908 32396
rect 62076 33124 62132 33134
rect 62076 32786 62132 33068
rect 62300 32900 62356 33516
rect 62412 33124 62468 35758
rect 62524 34692 62580 34702
rect 62636 34692 62692 37324
rect 62524 34690 62692 34692
rect 62524 34638 62526 34690
rect 62578 34638 62692 34690
rect 62524 34636 62692 34638
rect 62748 36482 62804 36494
rect 62748 36430 62750 36482
rect 62802 36430 62804 36482
rect 62748 35698 62804 36430
rect 62748 35646 62750 35698
rect 62802 35646 62804 35698
rect 62524 34626 62580 34636
rect 62636 34356 62692 34366
rect 62636 34262 62692 34300
rect 62748 33348 62804 35646
rect 62860 35028 62916 39200
rect 63308 36482 63364 36494
rect 63308 36430 63310 36482
rect 63362 36430 63364 36482
rect 62860 34962 62916 34972
rect 63196 35474 63252 35486
rect 63196 35422 63198 35474
rect 63250 35422 63252 35474
rect 63084 34356 63140 34366
rect 63084 33458 63140 34300
rect 63084 33406 63086 33458
rect 63138 33406 63140 33458
rect 63084 33394 63140 33406
rect 62748 33282 62804 33292
rect 62412 33058 62468 33068
rect 62524 33124 62580 33134
rect 62524 33122 62692 33124
rect 62524 33070 62526 33122
rect 62578 33070 62692 33122
rect 62524 33068 62692 33070
rect 62524 33058 62580 33068
rect 62300 32844 62580 32900
rect 62076 32734 62078 32786
rect 62130 32734 62132 32786
rect 62076 31892 62132 32734
rect 62524 32786 62580 32844
rect 62524 32734 62526 32786
rect 62578 32734 62580 32786
rect 62524 32722 62580 32734
rect 62636 32004 62692 33068
rect 62636 31938 62692 31948
rect 62972 32788 63028 32798
rect 62076 31826 62132 31836
rect 62972 27972 63028 32732
rect 63196 32788 63252 35422
rect 63308 34244 63364 36430
rect 63644 36258 63700 36270
rect 63644 36206 63646 36258
rect 63698 36206 63700 36258
rect 63532 35474 63588 35486
rect 63532 35422 63534 35474
rect 63586 35422 63588 35474
rect 63420 35028 63476 35038
rect 63420 34934 63476 34972
rect 63308 34188 63476 34244
rect 63308 34018 63364 34030
rect 63308 33966 63310 34018
rect 63362 33966 63364 34018
rect 63308 33348 63364 33966
rect 63420 33460 63476 34188
rect 63532 33684 63588 35422
rect 63532 33618 63588 33628
rect 63420 33394 63476 33404
rect 63308 33282 63364 33292
rect 63196 32722 63252 32732
rect 62972 27906 63028 27916
rect 61404 20132 61684 20188
rect 60172 8372 60452 8428
rect 59948 6580 60004 6590
rect 59948 6486 60004 6524
rect 59836 5908 59892 5918
rect 59836 5814 59892 5852
rect 60172 5012 60228 8372
rect 60732 8034 60788 8046
rect 60732 7982 60734 8034
rect 60786 7982 60788 8034
rect 60284 7364 60340 7374
rect 60732 7364 60788 7982
rect 61628 8034 61684 20132
rect 62188 8930 62244 8942
rect 62188 8878 62190 8930
rect 62242 8878 62244 8930
rect 62188 8484 62244 8878
rect 63084 8930 63140 8942
rect 63084 8878 63086 8930
rect 63138 8878 63140 8930
rect 63084 8428 63140 8878
rect 63532 8930 63588 8942
rect 63532 8878 63534 8930
rect 63586 8878 63588 8930
rect 62076 8036 62132 8046
rect 61628 7982 61630 8034
rect 61682 7982 61684 8034
rect 60956 7476 61012 7486
rect 60956 7382 61012 7420
rect 61292 7476 61348 7486
rect 61628 7476 61684 7982
rect 61852 8034 62132 8036
rect 61852 7982 62078 8034
rect 62130 7982 62132 8034
rect 61852 7980 62132 7982
rect 61852 7588 61908 7980
rect 62076 7970 62132 7980
rect 61292 7474 61684 7476
rect 61292 7422 61294 7474
rect 61346 7422 61684 7474
rect 61292 7420 61684 7422
rect 61740 7586 61908 7588
rect 61740 7534 61854 7586
rect 61906 7534 61908 7586
rect 61740 7532 61908 7534
rect 61292 7410 61348 7420
rect 60284 7362 60788 7364
rect 60284 7310 60286 7362
rect 60338 7310 60788 7362
rect 60284 7308 60788 7310
rect 60284 6468 60340 7308
rect 61628 7252 61684 7262
rect 60284 5908 60340 6412
rect 60732 6466 60788 6478
rect 60732 6414 60734 6466
rect 60786 6414 60788 6466
rect 60732 6020 60788 6414
rect 60732 5954 60788 5964
rect 61292 6468 61348 6478
rect 60284 5842 60340 5852
rect 60508 5906 60564 5918
rect 60508 5854 60510 5906
rect 60562 5854 60564 5906
rect 60508 5460 60564 5854
rect 60508 5394 60564 5404
rect 60284 5012 60340 5022
rect 60172 5010 60340 5012
rect 60172 4958 60286 5010
rect 60338 4958 60340 5010
rect 60172 4956 60340 4958
rect 60284 4946 60340 4956
rect 60620 5012 60676 5022
rect 60620 4918 60676 4956
rect 59612 4846 59614 4898
rect 59666 4846 59668 4898
rect 59612 4788 59668 4846
rect 59612 4722 59668 4732
rect 58828 4620 59220 4676
rect 58828 4562 58884 4620
rect 58828 4510 58830 4562
rect 58882 4510 58884 4562
rect 58828 4498 58884 4510
rect 61292 4450 61348 6412
rect 61292 4398 61294 4450
rect 61346 4398 61348 4450
rect 61292 4386 61348 4398
rect 58940 3668 58996 3678
rect 58716 3612 58940 3668
rect 58940 3554 58996 3612
rect 60844 3668 60900 3678
rect 58940 3502 58942 3554
rect 58994 3502 58996 3554
rect 58940 3490 58996 3502
rect 59836 3556 59892 3566
rect 59836 3462 59892 3500
rect 59612 3444 59668 3454
rect 58604 3330 58660 3342
rect 58604 3278 58606 3330
rect 58658 3278 58660 3330
rect 58604 3220 58660 3278
rect 58604 2772 58660 3164
rect 59500 3330 59556 3342
rect 59500 3278 59502 3330
rect 59554 3278 59556 3330
rect 59500 2996 59556 3278
rect 59500 2930 59556 2940
rect 58604 2706 58660 2716
rect 58380 2594 58436 2604
rect 59612 1764 59668 3388
rect 59500 1708 59668 1764
rect 59500 800 59556 1708
rect 60844 800 60900 3612
rect 61628 3554 61684 7196
rect 61740 6020 61796 7532
rect 61852 7522 61908 7532
rect 62076 7476 62132 7486
rect 62076 7382 62132 7420
rect 61964 6692 62020 6702
rect 62188 6692 62244 8428
rect 62636 8372 63364 8428
rect 62636 8370 62692 8372
rect 62636 8318 62638 8370
rect 62690 8318 62692 8370
rect 62636 8306 62692 8318
rect 62748 8034 62804 8046
rect 62748 7982 62750 8034
rect 62802 7982 62804 8034
rect 61964 6690 62244 6692
rect 61964 6638 61966 6690
rect 62018 6638 62244 6690
rect 61964 6636 62244 6638
rect 62412 6690 62468 6702
rect 62412 6638 62414 6690
rect 62466 6638 62468 6690
rect 61964 6626 62020 6636
rect 61852 6580 61908 6590
rect 61852 6486 61908 6524
rect 62412 6468 62468 6638
rect 62412 6402 62468 6412
rect 62748 6130 62804 7982
rect 62860 7588 62916 7598
rect 62860 7494 62916 7532
rect 62748 6078 62750 6130
rect 62802 6078 62804 6130
rect 62748 6066 62804 6078
rect 63084 6690 63140 6702
rect 63084 6638 63086 6690
rect 63138 6638 63140 6690
rect 63084 6132 63140 6638
rect 63084 6066 63140 6076
rect 61740 5954 61796 5964
rect 63308 5796 63364 8372
rect 63532 7812 63588 8878
rect 63644 8260 63700 36206
rect 63756 36036 63812 39200
rect 64316 37492 64372 37502
rect 64652 37492 64708 39200
rect 64652 37436 65156 37492
rect 63756 35980 64260 36036
rect 64204 35810 64260 35980
rect 64204 35758 64206 35810
rect 64258 35758 64260 35810
rect 63868 34804 63924 34814
rect 63868 34356 63924 34748
rect 63868 34224 63924 34300
rect 64204 33460 64260 35758
rect 64316 34916 64372 37436
rect 64652 37268 64708 37278
rect 64540 36596 64596 36606
rect 64540 36502 64596 36540
rect 64540 35924 64596 35934
rect 64652 35924 64708 37212
rect 64988 36484 65044 36494
rect 64988 36390 65044 36428
rect 64540 35922 64708 35924
rect 64540 35870 64542 35922
rect 64594 35870 64708 35922
rect 64540 35868 64708 35870
rect 64540 35858 64596 35868
rect 65100 35026 65156 37436
rect 65548 36484 65604 39200
rect 65324 36372 65380 36382
rect 65324 36278 65380 36316
rect 65100 34974 65102 35026
rect 65154 34974 65156 35026
rect 65100 34962 65156 34974
rect 64316 34914 64708 34916
rect 64316 34862 64318 34914
rect 64370 34862 64708 34914
rect 64316 34860 64708 34862
rect 64316 34850 64372 34860
rect 64652 34354 64708 34860
rect 64652 34302 64654 34354
rect 64706 34302 64708 34354
rect 64652 34290 64708 34302
rect 65436 34468 65492 34478
rect 65436 34354 65492 34412
rect 65436 34302 65438 34354
rect 65490 34302 65492 34354
rect 65436 34290 65492 34302
rect 64764 34244 64820 34254
rect 64540 33460 64596 33470
rect 64204 33458 64596 33460
rect 64204 33406 64542 33458
rect 64594 33406 64596 33458
rect 64204 33404 64596 33406
rect 64540 33394 64596 33404
rect 63756 33348 63812 33358
rect 63756 33254 63812 33292
rect 64204 33122 64260 33134
rect 64204 33070 64206 33122
rect 64258 33070 64260 33122
rect 64204 32788 64260 33070
rect 64204 32722 64260 32732
rect 64764 30884 64820 34188
rect 65100 33460 65156 33470
rect 65100 33366 65156 33404
rect 65548 33458 65604 36428
rect 65660 38164 65716 38174
rect 65660 36372 65716 38108
rect 66108 36596 66164 36606
rect 66108 36482 66164 36540
rect 66444 36596 66500 39200
rect 66444 36530 66500 36540
rect 66108 36430 66110 36482
rect 66162 36430 66164 36482
rect 65996 36372 66052 36382
rect 65660 36306 65716 36316
rect 65884 36370 66052 36372
rect 65884 36318 65998 36370
rect 66050 36318 66052 36370
rect 65884 36316 66052 36318
rect 65772 35810 65828 35822
rect 65772 35758 65774 35810
rect 65826 35758 65828 35810
rect 65772 34468 65828 35758
rect 65772 34402 65828 34412
rect 65548 33406 65550 33458
rect 65602 33406 65604 33458
rect 65548 33394 65604 33406
rect 65884 34018 65940 36316
rect 65996 36306 66052 36316
rect 66108 35700 66164 36430
rect 66780 36484 66836 36494
rect 66780 36390 66836 36428
rect 67116 36260 67172 36270
rect 67004 36258 67172 36260
rect 67004 36206 67118 36258
rect 67170 36206 67172 36258
rect 67004 36204 67172 36206
rect 66108 35568 66164 35644
rect 66668 35700 66724 35710
rect 66556 35476 66612 35486
rect 66556 35382 66612 35420
rect 66668 35028 66724 35644
rect 66108 34916 66164 34926
rect 66108 34914 66500 34916
rect 66108 34862 66110 34914
rect 66162 34862 66500 34914
rect 66668 34896 66724 34972
rect 66892 35474 66948 35486
rect 66892 35422 66894 35474
rect 66946 35422 66948 35474
rect 66108 34860 66500 34862
rect 66108 34850 66164 34860
rect 65884 33966 65886 34018
rect 65938 33966 65940 34018
rect 65884 32900 65940 33966
rect 65884 32834 65940 32844
rect 66332 34132 66388 34142
rect 64764 30818 64820 30828
rect 66332 20188 66388 34076
rect 66444 34018 66500 34860
rect 66444 33966 66446 34018
rect 66498 33966 66500 34018
rect 66444 31668 66500 33966
rect 66444 31602 66500 31612
rect 66332 20132 66500 20188
rect 64988 9604 65044 9614
rect 64540 9602 65044 9604
rect 64540 9550 64990 9602
rect 65042 9550 65044 9602
rect 64540 9548 65044 9550
rect 64540 9154 64596 9548
rect 64988 9538 65044 9548
rect 64540 9102 64542 9154
rect 64594 9102 64596 9154
rect 64540 8484 64596 9102
rect 65772 9154 65828 9166
rect 65772 9102 65774 9154
rect 65826 9102 65828 9154
rect 65436 9044 65492 9054
rect 64876 9042 65492 9044
rect 64876 8990 65438 9042
rect 65490 8990 65492 9042
rect 64876 8988 65492 8990
rect 64652 8820 64708 8830
rect 64652 8818 64820 8820
rect 64652 8766 64654 8818
rect 64706 8766 64820 8818
rect 64652 8764 64820 8766
rect 64652 8754 64708 8764
rect 64540 8372 64708 8428
rect 63644 8194 63700 8204
rect 63868 8258 63924 8270
rect 63868 8206 63870 8258
rect 63922 8206 63924 8258
rect 63532 7756 63700 7812
rect 63532 7586 63588 7598
rect 63532 7534 63534 7586
rect 63586 7534 63588 7586
rect 63420 7476 63476 7486
rect 63420 7382 63476 7420
rect 63532 7252 63588 7534
rect 63532 7186 63588 7196
rect 62860 5124 62916 5134
rect 62860 5030 62916 5068
rect 61628 3502 61630 3554
rect 61682 3502 61684 3554
rect 61628 3490 61684 3502
rect 62188 5012 62244 5022
rect 60956 3444 61012 3454
rect 60956 3350 61012 3388
rect 62188 800 62244 4956
rect 62412 3556 62468 3566
rect 62412 3462 62468 3500
rect 62748 3556 62804 3566
rect 62748 3442 62804 3500
rect 62748 3390 62750 3442
rect 62802 3390 62804 3442
rect 62748 3378 62804 3390
rect 63308 3442 63364 5740
rect 63532 5682 63588 5694
rect 63532 5630 63534 5682
rect 63586 5630 63588 5682
rect 63532 3780 63588 5630
rect 63532 3714 63588 3724
rect 63644 3556 63700 7756
rect 63868 7476 63924 8206
rect 64540 8260 64596 8270
rect 64540 8166 64596 8204
rect 63980 8148 64036 8158
rect 63980 8054 64036 8092
rect 63868 7410 63924 7420
rect 64204 7588 64260 7598
rect 64204 7474 64260 7532
rect 64204 7422 64206 7474
rect 64258 7422 64260 7474
rect 64204 7410 64260 7422
rect 64540 7252 64596 7262
rect 64316 7250 64596 7252
rect 64316 7198 64542 7250
rect 64594 7198 64596 7250
rect 64316 7196 64596 7198
rect 63980 6132 64036 6142
rect 63980 6038 64036 6076
rect 64316 6018 64372 7196
rect 64540 7186 64596 7196
rect 64652 6692 64708 8372
rect 64652 6626 64708 6636
rect 64764 6580 64820 8764
rect 64876 8482 64932 8988
rect 65436 8978 65492 8988
rect 64876 8430 64878 8482
rect 64930 8430 64932 8482
rect 64876 8418 64932 8430
rect 65772 8372 65828 9102
rect 66332 8930 66388 8942
rect 66332 8878 66334 8930
rect 66386 8878 66388 8930
rect 66332 8428 66388 8878
rect 65772 8306 65828 8316
rect 65996 8372 66388 8428
rect 65996 8258 66052 8372
rect 65996 8206 65998 8258
rect 66050 8206 66052 8258
rect 65436 8148 65492 8158
rect 65324 6580 65380 6590
rect 64764 6578 65380 6580
rect 64764 6526 65326 6578
rect 65378 6526 65380 6578
rect 64764 6524 65380 6526
rect 65324 6514 65380 6524
rect 65324 6132 65380 6142
rect 65436 6132 65492 8092
rect 65548 8146 65604 8158
rect 65548 8094 65550 8146
rect 65602 8094 65604 8146
rect 65548 7476 65604 8094
rect 65996 8036 66052 8206
rect 65548 7382 65604 7420
rect 65660 7586 65716 7598
rect 65660 7534 65662 7586
rect 65714 7534 65716 7586
rect 65324 6130 65492 6132
rect 65324 6078 65326 6130
rect 65378 6078 65492 6130
rect 65324 6076 65492 6078
rect 65324 6066 65380 6076
rect 64316 5966 64318 6018
rect 64370 5966 64372 6018
rect 64316 5954 64372 5966
rect 63980 5236 64036 5246
rect 63980 5142 64036 5180
rect 63868 5124 63924 5134
rect 63868 4338 63924 5068
rect 65660 5012 65716 7534
rect 65996 6356 66052 7980
rect 66444 7700 66500 20132
rect 66556 8148 66612 8158
rect 66556 8054 66612 8092
rect 66332 7476 66388 7486
rect 66444 7476 66500 7644
rect 66892 7588 66948 35422
rect 67004 34132 67060 36204
rect 67116 36194 67172 36204
rect 67116 34916 67172 34926
rect 67116 34822 67172 34860
rect 67340 34916 67396 39200
rect 68236 36932 68292 39200
rect 68236 36866 68292 36876
rect 68796 37828 68852 37838
rect 67900 36596 67956 36606
rect 67676 36484 67732 36494
rect 67340 34850 67396 34860
rect 67452 35476 67508 35486
rect 67004 34066 67060 34076
rect 67452 34018 67508 35420
rect 67564 34916 67620 34926
rect 67564 34822 67620 34860
rect 67676 34356 67732 36428
rect 67788 36372 67844 36382
rect 67788 36278 67844 36316
rect 67900 35810 67956 36540
rect 68796 36596 68852 37772
rect 68796 36530 68852 36540
rect 68908 36932 68964 36942
rect 68908 36594 68964 36876
rect 68908 36542 68910 36594
rect 68962 36542 68964 36594
rect 68908 36530 68964 36542
rect 67900 35758 67902 35810
rect 67954 35758 67956 35810
rect 67900 35746 67956 35758
rect 68572 36148 68628 36158
rect 67900 34692 67956 34702
rect 67900 34690 68068 34692
rect 67900 34638 67902 34690
rect 67954 34638 68068 34690
rect 67900 34636 68068 34638
rect 67900 34626 67956 34636
rect 67900 34356 67956 34366
rect 67676 34354 67956 34356
rect 67676 34302 67902 34354
rect 67954 34302 67956 34354
rect 67676 34300 67956 34302
rect 67452 33966 67454 34018
rect 67506 33966 67508 34018
rect 67452 32564 67508 33966
rect 67452 32498 67508 32508
rect 67900 25508 67956 34300
rect 68012 30212 68068 34636
rect 68572 33796 68628 36092
rect 68796 35700 68852 35710
rect 68796 35698 69076 35700
rect 68796 35646 68798 35698
rect 68850 35646 69076 35698
rect 68796 35644 69076 35646
rect 68796 35634 68852 35644
rect 68684 35028 68740 35038
rect 68684 34934 68740 34972
rect 68572 33730 68628 33740
rect 69020 34018 69076 35644
rect 69132 35028 69188 39200
rect 69692 37828 69748 37838
rect 69692 36482 69748 37772
rect 70028 36932 70084 39200
rect 70028 36866 70084 36876
rect 70588 36932 70644 36942
rect 70588 36594 70644 36876
rect 70588 36542 70590 36594
rect 70642 36542 70644 36594
rect 70588 36530 70644 36542
rect 69692 36430 69694 36482
rect 69746 36430 69748 36482
rect 69692 36372 69748 36430
rect 69692 36306 69748 36316
rect 70812 36148 70868 36158
rect 70812 35922 70868 36092
rect 70812 35870 70814 35922
rect 70866 35870 70868 35922
rect 70812 35858 70868 35870
rect 69916 35810 69972 35822
rect 69916 35758 69918 35810
rect 69970 35758 69972 35810
rect 69580 35698 69636 35710
rect 69580 35646 69582 35698
rect 69634 35646 69636 35698
rect 69580 35252 69636 35646
rect 69916 35700 69972 35758
rect 70476 35812 70532 35822
rect 70476 35718 70532 35756
rect 70924 35812 70980 39200
rect 71484 36484 71540 36494
rect 71484 36482 71652 36484
rect 71484 36430 71486 36482
rect 71538 36430 71652 36482
rect 71484 36428 71652 36430
rect 71484 36418 71540 36428
rect 69916 35634 69972 35644
rect 69580 35186 69636 35196
rect 70140 35252 70196 35262
rect 69132 34916 69188 34972
rect 70140 35026 70196 35196
rect 70140 34974 70142 35026
rect 70194 34974 70196 35026
rect 70140 34962 70196 34974
rect 70924 35028 70980 35756
rect 71596 35252 71652 36428
rect 71820 35586 71876 39200
rect 72492 37156 72548 37166
rect 71820 35534 71822 35586
rect 71874 35534 71876 35586
rect 71820 35522 71876 35534
rect 72380 36482 72436 36494
rect 72380 36430 72382 36482
rect 72434 36430 72436 36482
rect 71036 35028 71092 35038
rect 70924 35026 71092 35028
rect 70924 34974 71038 35026
rect 71090 34974 71092 35026
rect 70924 34972 71092 34974
rect 71036 34962 71092 34972
rect 71596 35026 71652 35196
rect 71596 34974 71598 35026
rect 71650 34974 71652 35026
rect 71596 34962 71652 34974
rect 72044 35028 72100 35038
rect 72044 34934 72100 34972
rect 69356 34916 69412 34926
rect 69132 34914 69412 34916
rect 69132 34862 69358 34914
rect 69410 34862 69412 34914
rect 69132 34860 69412 34862
rect 69356 34850 69412 34860
rect 69020 33966 69022 34018
rect 69074 33966 69076 34018
rect 68012 30146 68068 30156
rect 69020 28532 69076 33966
rect 69692 34690 69748 34702
rect 69692 34638 69694 34690
rect 69746 34638 69748 34690
rect 69692 31892 69748 34638
rect 72156 34020 72212 34030
rect 72380 34020 72436 36430
rect 72492 35026 72548 37100
rect 72604 36260 72660 36270
rect 72604 35698 72660 36204
rect 72604 35646 72606 35698
rect 72658 35646 72660 35698
rect 72604 35634 72660 35646
rect 72492 34974 72494 35026
rect 72546 34974 72548 35026
rect 72492 34962 72548 34974
rect 72716 35028 72772 39200
rect 72828 38724 72884 38734
rect 72828 36148 72884 38668
rect 73612 37828 73668 39200
rect 73388 37772 73668 37828
rect 73388 36594 73444 37772
rect 73388 36542 73390 36594
rect 73442 36542 73444 36594
rect 73388 36530 73444 36542
rect 73836 37156 73892 37166
rect 72828 36082 72884 36092
rect 73724 36148 73780 36158
rect 73724 35698 73780 36092
rect 73724 35646 73726 35698
rect 73778 35646 73780 35698
rect 73724 35634 73780 35646
rect 72716 34916 72772 34972
rect 73276 35364 73332 35374
rect 72940 34916 72996 34926
rect 72716 34914 72996 34916
rect 72716 34862 72942 34914
rect 72994 34862 72996 34914
rect 72716 34860 72996 34862
rect 72940 34850 72996 34860
rect 73276 34802 73332 35308
rect 73836 34914 73892 37100
rect 74396 36820 74452 36830
rect 74396 36482 74452 36764
rect 74396 36430 74398 36482
rect 74450 36430 74452 36482
rect 74396 36418 74452 36430
rect 74284 36372 74340 36382
rect 73948 36370 74340 36372
rect 73948 36318 74286 36370
rect 74338 36318 74340 36370
rect 73948 36316 74340 36318
rect 73948 35922 74004 36316
rect 74284 36306 74340 36316
rect 73948 35870 73950 35922
rect 74002 35870 74004 35922
rect 73948 35858 74004 35870
rect 74508 36148 74564 39200
rect 75068 36932 75124 36942
rect 73836 34862 73838 34914
rect 73890 34862 73892 34914
rect 73836 34850 73892 34862
rect 74284 35588 74340 35598
rect 73276 34750 73278 34802
rect 73330 34750 73332 34802
rect 73276 34738 73332 34750
rect 74172 34690 74228 34702
rect 74172 34638 74174 34690
rect 74226 34638 74228 34690
rect 73164 34580 73220 34590
rect 73164 34356 73220 34524
rect 73836 34580 73892 34590
rect 73276 34356 73332 34366
rect 73164 34354 73332 34356
rect 73164 34302 73278 34354
rect 73330 34302 73332 34354
rect 73164 34300 73332 34302
rect 73276 34290 73332 34300
rect 73836 34242 73892 34524
rect 73948 34356 74004 34366
rect 73948 34262 74004 34300
rect 73836 34190 73838 34242
rect 73890 34190 73892 34242
rect 73836 34178 73892 34190
rect 74172 34244 74228 34638
rect 74172 34178 74228 34188
rect 72716 34020 72772 34030
rect 72380 34018 72772 34020
rect 72380 33966 72718 34018
rect 72770 33966 72772 34018
rect 72380 33964 72772 33966
rect 72156 32340 72212 33964
rect 72716 33460 72772 33964
rect 72716 33394 72772 33404
rect 73836 33460 73892 33470
rect 74284 33460 74340 35532
rect 74396 34804 74452 34814
rect 74396 34354 74452 34748
rect 74396 34302 74398 34354
rect 74450 34302 74452 34354
rect 74396 34290 74452 34302
rect 73836 33458 74340 33460
rect 73836 33406 73838 33458
rect 73890 33406 74286 33458
rect 74338 33406 74340 33458
rect 73836 33404 74340 33406
rect 74508 33460 74564 36092
rect 74620 36820 74676 36830
rect 74620 35698 74676 36764
rect 75068 36708 75124 36876
rect 75068 36706 75236 36708
rect 75068 36654 75070 36706
rect 75122 36654 75236 36706
rect 75068 36652 75236 36654
rect 75068 36642 75124 36652
rect 74852 36092 75116 36102
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 74852 36026 75116 36036
rect 74620 35646 74622 35698
rect 74674 35646 74676 35698
rect 74620 35588 74676 35646
rect 74620 35522 74676 35532
rect 74732 35810 74788 35822
rect 74732 35758 74734 35810
rect 74786 35758 74788 35810
rect 74732 35364 74788 35758
rect 74732 35298 74788 35308
rect 75180 35140 75236 36652
rect 75404 36596 75460 39200
rect 75068 35084 75236 35140
rect 75292 36540 75460 36596
rect 74732 34916 74788 34926
rect 74732 34692 74788 34860
rect 75068 34692 75124 35084
rect 75292 34916 75348 36540
rect 75404 36260 75460 36270
rect 75404 36258 75572 36260
rect 75404 36206 75406 36258
rect 75458 36206 75572 36258
rect 75404 36204 75572 36206
rect 75404 36194 75460 36204
rect 75404 35476 75460 35486
rect 75404 35382 75460 35420
rect 75292 34850 75348 34860
rect 75404 34804 75460 34814
rect 75292 34692 75348 34702
rect 75404 34692 75460 34748
rect 75068 34636 75236 34692
rect 74732 34626 74788 34636
rect 74852 34524 75116 34534
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 74852 34458 75116 34468
rect 75180 34354 75236 34636
rect 75292 34690 75460 34692
rect 75292 34638 75294 34690
rect 75346 34638 75460 34690
rect 75292 34636 75460 34638
rect 75292 34626 75348 34636
rect 75404 34580 75460 34636
rect 75404 34514 75460 34524
rect 75180 34302 75182 34354
rect 75234 34302 75236 34354
rect 75180 34290 75236 34302
rect 74620 33460 74676 33470
rect 74508 33458 74676 33460
rect 74508 33406 74622 33458
rect 74674 33406 74676 33458
rect 74508 33404 74676 33406
rect 73836 33394 73892 33404
rect 74284 33394 74340 33404
rect 74620 33394 74676 33404
rect 74852 32956 75116 32966
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 74852 32890 75116 32900
rect 72156 32274 72212 32284
rect 69692 31826 69748 31836
rect 74852 31388 75116 31398
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 74852 31322 75116 31332
rect 74852 29820 75116 29830
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 74852 29754 75116 29764
rect 69020 28466 69076 28476
rect 74852 28252 75116 28262
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 74852 28186 75116 28196
rect 74852 26684 75116 26694
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 74852 26618 75116 26628
rect 67900 25442 67956 25452
rect 74852 25116 75116 25126
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 74852 25050 75116 25060
rect 75516 24724 75572 36204
rect 75852 35588 75908 35598
rect 75740 35474 75796 35486
rect 75740 35422 75742 35474
rect 75794 35422 75796 35474
rect 75628 34916 75684 34926
rect 75628 34354 75684 34860
rect 75628 34302 75630 34354
rect 75682 34302 75684 34354
rect 75628 34290 75684 34302
rect 75516 24658 75572 24668
rect 73052 24612 73108 24622
rect 68796 22932 68852 22942
rect 68796 17780 68852 22876
rect 69804 21028 69860 21038
rect 68908 17780 68964 17790
rect 68796 17724 68908 17780
rect 67340 15428 67396 15438
rect 67004 8260 67060 8270
rect 67004 8166 67060 8204
rect 67228 7700 67284 7710
rect 67228 7606 67284 7644
rect 66892 7522 66948 7532
rect 66332 7474 66500 7476
rect 66332 7422 66334 7474
rect 66386 7422 66500 7474
rect 66332 7420 66500 7422
rect 66332 7410 66388 7420
rect 66108 7252 66164 7262
rect 66108 6690 66164 7196
rect 66668 7250 66724 7262
rect 66668 7198 66670 7250
rect 66722 7198 66724 7250
rect 66108 6638 66110 6690
rect 66162 6638 66164 6690
rect 66108 6626 66164 6638
rect 66332 6692 66388 6702
rect 65996 6290 66052 6300
rect 66108 6132 66164 6142
rect 66108 6038 66164 6076
rect 65324 4956 65716 5012
rect 66108 5460 66164 5470
rect 65324 4562 65380 4956
rect 65324 4510 65326 4562
rect 65378 4510 65380 4562
rect 65324 4498 65380 4510
rect 63868 4286 63870 4338
rect 63922 4286 63924 4338
rect 63868 4274 63924 4286
rect 63308 3390 63310 3442
rect 63362 3390 63364 3442
rect 63308 3378 63364 3390
rect 63532 3444 63588 3454
rect 63644 3424 63700 3500
rect 64988 3556 65044 3566
rect 64876 3444 64932 3454
rect 63532 800 63588 3388
rect 64876 3350 64932 3388
rect 64988 1764 65044 3500
rect 65548 3554 65604 4956
rect 66108 4562 66164 5404
rect 66108 4510 66110 4562
rect 66162 4510 66164 4562
rect 66108 4498 66164 4510
rect 65548 3502 65550 3554
rect 65602 3502 65604 3554
rect 65548 3490 65604 3502
rect 66332 3330 66388 6636
rect 66668 6690 66724 7198
rect 66668 6638 66670 6690
rect 66722 6638 66724 6690
rect 66668 6626 66724 6638
rect 66892 6466 66948 6478
rect 66892 6414 66894 6466
rect 66946 6414 66948 6466
rect 66892 4340 66948 6414
rect 67116 5124 67172 5134
rect 67116 5030 67172 5068
rect 66892 4274 66948 4284
rect 66556 4228 66612 4238
rect 66556 3668 66612 4172
rect 66556 3554 66612 3612
rect 66556 3502 66558 3554
rect 66610 3502 66612 3554
rect 66556 3490 66612 3502
rect 66332 3278 66334 3330
rect 66386 3278 66388 3330
rect 66332 3266 66388 3278
rect 67228 3332 67284 3342
rect 67340 3332 67396 15372
rect 68796 15428 68852 17724
rect 68908 17714 68964 17724
rect 68796 15362 68852 15372
rect 68348 8372 68404 8382
rect 67676 6692 67732 6702
rect 68124 6692 68180 6702
rect 67732 6636 67844 6692
rect 67676 6598 67732 6636
rect 67564 6466 67620 6478
rect 67564 6414 67566 6466
rect 67618 6414 67620 6466
rect 67564 6132 67620 6414
rect 67564 6066 67620 6076
rect 67676 5460 67732 5470
rect 67676 5346 67732 5404
rect 67676 5294 67678 5346
rect 67730 5294 67732 5346
rect 67676 5282 67732 5294
rect 67788 5236 67844 6636
rect 68124 6598 68180 6636
rect 68348 5906 68404 8316
rect 68348 5854 68350 5906
rect 68402 5854 68404 5906
rect 68348 5842 68404 5854
rect 68572 6692 68628 6702
rect 68572 6466 68628 6636
rect 69356 6692 69412 6702
rect 69356 6598 69412 6636
rect 68572 6414 68574 6466
rect 68626 6414 68628 6466
rect 68236 5236 68292 5246
rect 67788 5234 68292 5236
rect 67788 5182 67790 5234
rect 67842 5182 68238 5234
rect 68290 5182 68292 5234
rect 67788 5180 68292 5182
rect 67788 5170 67844 5180
rect 68236 5170 68292 5180
rect 68348 4340 68404 4350
rect 68348 4246 68404 4284
rect 67564 3556 67620 3566
rect 67564 3462 67620 3500
rect 67228 3330 67396 3332
rect 67228 3278 67230 3330
rect 67282 3278 67396 3330
rect 67228 3276 67396 3278
rect 67676 3444 67732 3454
rect 67228 3266 67284 3276
rect 67676 1764 67732 3388
rect 64876 1708 65044 1764
rect 67564 1708 67732 1764
rect 64876 800 64932 1708
rect 67564 800 67620 1708
rect 5964 140 6468 196
rect 6412 84 6468 140
rect 6412 18 6468 28
rect 7056 0 7168 800
rect 8400 0 8512 800
rect 9744 0 9856 800
rect 11088 0 11200 800
rect 12432 0 12544 800
rect 13776 0 13888 800
rect 15120 0 15232 800
rect 16464 0 16576 800
rect 17808 0 17920 800
rect 19152 0 19264 800
rect 20496 0 20608 800
rect 21840 0 21952 800
rect 23184 0 23296 800
rect 24528 0 24640 800
rect 25872 0 25984 800
rect 27216 0 27328 800
rect 28560 0 28672 800
rect 29904 0 30016 800
rect 31248 0 31360 800
rect 32592 0 32704 800
rect 33936 0 34048 800
rect 35280 0 35392 800
rect 36624 0 36736 800
rect 37968 0 38080 800
rect 39312 0 39424 800
rect 40656 0 40768 800
rect 42000 0 42112 800
rect 43344 0 43456 800
rect 44688 0 44800 800
rect 46032 0 46144 800
rect 47376 0 47488 800
rect 48720 0 48832 800
rect 50064 0 50176 800
rect 51408 0 51520 800
rect 52752 0 52864 800
rect 54096 0 54208 800
rect 55440 0 55552 800
rect 56784 0 56896 800
rect 58128 0 58240 800
rect 59472 0 59584 800
rect 60816 0 60928 800
rect 62160 0 62272 800
rect 63504 0 63616 800
rect 64848 0 64960 800
rect 66192 0 66304 800
rect 67536 0 67648 800
rect 68572 84 68628 6414
rect 69020 5906 69076 5918
rect 69020 5854 69022 5906
rect 69074 5854 69076 5906
rect 69020 5796 69076 5854
rect 69356 5796 69412 5806
rect 69020 5794 69412 5796
rect 69020 5742 69358 5794
rect 69410 5742 69412 5794
rect 69020 5740 69412 5742
rect 69356 5348 69412 5740
rect 69356 5282 69412 5292
rect 68908 5236 68964 5246
rect 68908 4338 68964 5180
rect 69692 5236 69748 5246
rect 69692 5142 69748 5180
rect 69804 5012 69860 20972
rect 71372 21028 71428 21038
rect 69356 4900 69412 4910
rect 69356 4898 69524 4900
rect 69356 4846 69358 4898
rect 69410 4846 69524 4898
rect 69356 4844 69524 4846
rect 69356 4834 69412 4844
rect 68908 4286 68910 4338
rect 68962 4286 68964 4338
rect 68908 4274 68964 4286
rect 69468 4338 69524 4844
rect 69804 4562 69860 4956
rect 69804 4510 69806 4562
rect 69858 4510 69860 4562
rect 69804 4498 69860 4510
rect 70140 5684 70196 5694
rect 69468 4286 69470 4338
rect 69522 4286 69524 4338
rect 68796 3444 68852 3454
rect 68796 3350 68852 3388
rect 68908 924 69188 980
rect 68908 800 68964 924
rect 68572 18 68628 28
rect 68880 0 68992 800
rect 69132 756 69188 924
rect 69468 756 69524 4286
rect 69692 3556 69748 3566
rect 70140 3556 70196 5628
rect 70700 5124 70756 5134
rect 70252 4564 70308 4574
rect 70252 4228 70308 4508
rect 70700 4340 70756 5068
rect 71372 4788 71428 20972
rect 71372 4722 71428 4732
rect 72604 6578 72660 6590
rect 72604 6526 72606 6578
rect 72658 6526 72660 6578
rect 72604 5122 72660 6526
rect 72604 5070 72606 5122
rect 72658 5070 72660 5122
rect 70700 4246 70756 4284
rect 72604 4340 72660 5070
rect 73052 5012 73108 24556
rect 74852 23548 75116 23558
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 74852 23482 75116 23492
rect 74852 21980 75116 21990
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 74852 21914 75116 21924
rect 74852 20412 75116 20422
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 74852 20346 75116 20356
rect 73052 4946 73108 4956
rect 74172 19460 74228 19470
rect 72604 4246 72660 4284
rect 70252 4162 70308 4172
rect 70252 3556 70308 3566
rect 69692 3554 70308 3556
rect 69692 3502 69694 3554
rect 69746 3502 70254 3554
rect 70306 3502 70308 3554
rect 69692 3500 70308 3502
rect 69692 3490 69748 3500
rect 70252 3490 70308 3500
rect 70588 3556 70644 3566
rect 70588 3462 70644 3500
rect 71708 3556 71764 3566
rect 71708 3462 71764 3500
rect 73612 3556 73668 3566
rect 73612 3462 73668 3500
rect 71596 3444 71652 3454
rect 71596 800 71652 3388
rect 72716 3444 72772 3454
rect 72716 3350 72772 3388
rect 72940 3444 72996 3454
rect 72940 800 72996 3388
rect 74172 3330 74228 19404
rect 74852 18844 75116 18854
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 74852 18778 75116 18788
rect 74852 17276 75116 17286
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 74852 17210 75116 17220
rect 74852 15708 75116 15718
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 74852 15642 75116 15652
rect 74852 14140 75116 14150
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 74852 14074 75116 14084
rect 74852 12572 75116 12582
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 74852 12506 75116 12516
rect 75740 11172 75796 35422
rect 75852 34916 75908 35532
rect 76300 35028 76356 39200
rect 76748 36482 76804 36494
rect 76748 36430 76750 36482
rect 76802 36430 76804 36482
rect 76636 36372 76692 36382
rect 76300 34962 76356 34972
rect 76412 36370 76692 36372
rect 76412 36318 76638 36370
rect 76690 36318 76692 36370
rect 76412 36316 76692 36318
rect 76188 34916 76244 34926
rect 75852 34914 76132 34916
rect 75852 34862 75854 34914
rect 75906 34862 76132 34914
rect 75852 34860 76132 34862
rect 75852 34850 75908 34860
rect 75964 34690 76020 34702
rect 75964 34638 75966 34690
rect 76018 34638 76020 34690
rect 75964 34356 76020 34638
rect 76076 34356 76132 34860
rect 76188 34822 76244 34860
rect 76188 34356 76244 34366
rect 76076 34354 76244 34356
rect 76076 34302 76190 34354
rect 76242 34302 76244 34354
rect 76076 34300 76244 34302
rect 75964 34290 76020 34300
rect 76188 34290 76244 34300
rect 76076 33124 76132 33134
rect 76412 33124 76468 36316
rect 76636 36306 76692 36316
rect 76748 35700 76804 36430
rect 76636 35698 76804 35700
rect 76636 35646 76750 35698
rect 76802 35646 76804 35698
rect 76636 35644 76804 35646
rect 76636 34692 76692 35644
rect 76748 35634 76804 35644
rect 76860 35810 76916 35822
rect 76860 35758 76862 35810
rect 76914 35758 76916 35810
rect 76636 34598 76692 34636
rect 76748 35476 76804 35486
rect 76076 33122 76468 33124
rect 76076 33070 76078 33122
rect 76130 33070 76468 33122
rect 76076 33068 76468 33070
rect 76748 34354 76804 35420
rect 76748 34302 76750 34354
rect 76802 34302 76804 34354
rect 76076 32676 76132 33068
rect 76076 32610 76132 32620
rect 76748 31780 76804 34302
rect 76860 34020 76916 35758
rect 77196 35588 77252 39200
rect 78092 36820 78148 39200
rect 78092 36754 78148 36764
rect 77196 35522 77252 35532
rect 77420 36482 77476 36494
rect 77420 36430 77422 36482
rect 77474 36430 77476 36482
rect 77308 34916 77364 34926
rect 77308 34822 77364 34860
rect 77420 34356 77476 36430
rect 78764 36372 78820 36382
rect 78764 36278 78820 36316
rect 77756 36258 77812 36270
rect 77756 36206 77758 36258
rect 77810 36206 77812 36258
rect 77532 36036 77588 36046
rect 77532 35698 77588 35980
rect 77532 35646 77534 35698
rect 77586 35646 77588 35698
rect 77532 35634 77588 35646
rect 77420 34290 77476 34300
rect 76860 33954 76916 33964
rect 77196 34020 77252 34030
rect 77196 33926 77252 33964
rect 76748 31714 76804 31724
rect 75740 11106 75796 11116
rect 74852 11004 75116 11014
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 74852 10938 75116 10948
rect 74852 9436 75116 9446
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 74852 9370 75116 9380
rect 74852 7868 75116 7878
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 74852 7802 75116 7812
rect 76300 7586 76356 7598
rect 76300 7534 76302 7586
rect 76354 7534 76356 7586
rect 75628 7364 75684 7374
rect 76300 7364 76356 7534
rect 75628 7362 76356 7364
rect 75628 7310 75630 7362
rect 75682 7310 76356 7362
rect 75628 7308 76356 7310
rect 76860 7586 76916 7598
rect 76860 7534 76862 7586
rect 76914 7534 76916 7586
rect 75628 7298 75684 7308
rect 75628 6804 75684 6814
rect 75628 6710 75684 6748
rect 75292 6468 75348 6478
rect 75180 6466 75348 6468
rect 75180 6414 75294 6466
rect 75346 6414 75348 6466
rect 75180 6412 75348 6414
rect 74852 6300 75116 6310
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 74852 6234 75116 6244
rect 75068 5908 75124 5918
rect 75180 5908 75236 6412
rect 75292 6402 75348 6412
rect 75068 5906 75236 5908
rect 75068 5854 75070 5906
rect 75122 5854 75236 5906
rect 75068 5852 75236 5854
rect 75292 6018 75348 6030
rect 75292 5966 75294 6018
rect 75346 5966 75348 6018
rect 75068 5842 75124 5852
rect 75292 5124 75348 5966
rect 75740 5684 75796 7308
rect 76412 7140 76468 7150
rect 76412 6690 76468 7084
rect 76860 7140 76916 7534
rect 77084 7476 77140 7486
rect 77084 7382 77140 7420
rect 76860 7074 76916 7084
rect 77420 7250 77476 7262
rect 77420 7198 77422 7250
rect 77474 7198 77476 7250
rect 76412 6638 76414 6690
rect 76466 6638 76468 6690
rect 76412 6626 76468 6638
rect 77420 6690 77476 7198
rect 77756 6804 77812 36206
rect 78428 36260 78484 36270
rect 78428 36166 78484 36204
rect 78540 35700 78596 35710
rect 78540 35606 78596 35644
rect 77868 35474 77924 35486
rect 77868 35422 77870 35474
rect 77922 35422 77924 35474
rect 77868 31948 77924 35422
rect 78092 35140 78148 35150
rect 78428 35140 78484 35150
rect 78148 35084 78428 35140
rect 78092 35074 78148 35084
rect 78428 35074 78484 35084
rect 77980 35028 78036 35038
rect 77980 34934 78036 34972
rect 78204 34356 78260 34366
rect 78204 34132 78260 34300
rect 78764 34356 78820 34366
rect 78764 34262 78820 34300
rect 78988 34356 79044 39200
rect 79436 36372 79492 36382
rect 79212 36260 79268 36270
rect 79100 36258 79268 36260
rect 79100 36206 79214 36258
rect 79266 36206 79268 36258
rect 79100 36204 79268 36206
rect 79100 35700 79156 36204
rect 79212 36194 79268 36204
rect 79100 35634 79156 35644
rect 79212 35588 79268 35598
rect 79212 35494 79268 35532
rect 79436 34692 79492 36316
rect 79884 35252 79940 39200
rect 80332 38836 80388 38846
rect 80332 36036 80388 38780
rect 80556 37604 80612 37614
rect 80332 35922 80388 35980
rect 80332 35870 80334 35922
rect 80386 35870 80388 35922
rect 80332 35858 80388 35870
rect 80444 36482 80500 36494
rect 80444 36430 80446 36482
rect 80498 36430 80500 36482
rect 79884 35186 79940 35196
rect 79548 34916 79604 34926
rect 79548 34914 80164 34916
rect 79548 34862 79550 34914
rect 79602 34862 80164 34914
rect 79548 34860 80164 34862
rect 79548 34850 79604 34860
rect 79436 34626 79492 34636
rect 79772 34690 79828 34702
rect 79772 34638 79774 34690
rect 79826 34638 79828 34690
rect 78988 34290 79044 34300
rect 79436 34356 79492 34366
rect 78204 34066 78260 34076
rect 79212 34242 79268 34254
rect 79212 34190 79214 34242
rect 79266 34190 79268 34242
rect 77868 31892 78484 31948
rect 78204 12740 78260 12750
rect 77980 7362 78036 7374
rect 77980 7310 77982 7362
rect 78034 7310 78036 7362
rect 77980 7140 78036 7310
rect 77980 6804 78036 7084
rect 78092 6804 78148 6814
rect 77980 6802 78148 6804
rect 77980 6750 78094 6802
rect 78146 6750 78148 6802
rect 77980 6748 78148 6750
rect 77756 6738 77812 6748
rect 78092 6738 78148 6748
rect 77420 6638 77422 6690
rect 77474 6638 77476 6690
rect 77420 6626 77476 6638
rect 75740 5590 75796 5628
rect 76300 6578 76356 6590
rect 76300 6526 76302 6578
rect 76354 6526 76356 6578
rect 76300 6468 76356 6526
rect 75516 5236 75572 5246
rect 75516 5142 75572 5180
rect 75292 5058 75348 5068
rect 74852 4732 75116 4742
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 74852 4666 75116 4676
rect 74844 4340 74900 4350
rect 74844 4246 74900 4284
rect 75628 3668 75684 3678
rect 75628 3574 75684 3612
rect 76300 3556 76356 6412
rect 77644 6466 77700 6478
rect 77644 6414 77646 6466
rect 77698 6414 77700 6466
rect 76524 6020 76580 6030
rect 76524 5926 76580 5964
rect 77644 5908 77700 6414
rect 77644 5842 77700 5852
rect 77420 5236 77476 5246
rect 77420 5122 77476 5180
rect 77420 5070 77422 5122
rect 77474 5070 77476 5122
rect 77420 5058 77476 5070
rect 77756 5124 77812 5134
rect 77756 5030 77812 5068
rect 76300 3490 76356 3500
rect 77532 3668 77588 3678
rect 77532 3554 77588 3612
rect 77532 3502 77534 3554
rect 77586 3502 77588 3554
rect 77532 3490 77588 3502
rect 74508 3444 74564 3454
rect 74508 3350 74564 3388
rect 74956 3444 75012 3454
rect 74956 3350 75012 3388
rect 75628 3444 75684 3454
rect 74172 3278 74174 3330
rect 74226 3278 74228 3330
rect 74172 2884 74228 3278
rect 74852 3164 75116 3174
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 74852 3098 75116 3108
rect 74172 2818 74228 2828
rect 75628 800 75684 3388
rect 76636 3444 76692 3454
rect 76636 3350 76692 3388
rect 76972 3444 77028 3454
rect 76972 800 77028 3388
rect 78092 3332 78148 3342
rect 78204 3332 78260 12684
rect 78428 7698 78484 31892
rect 79212 27636 79268 34190
rect 79436 34130 79492 34300
rect 79436 34078 79438 34130
rect 79490 34078 79492 34130
rect 79436 34066 79492 34078
rect 79772 32676 79828 34638
rect 79772 32610 79828 32620
rect 80108 34692 80164 34860
rect 80220 34692 80276 34702
rect 80108 34690 80276 34692
rect 80108 34638 80222 34690
rect 80274 34638 80276 34690
rect 80108 34636 80276 34638
rect 79212 27570 79268 27580
rect 80108 14308 80164 34636
rect 80220 34626 80276 34636
rect 80444 34244 80500 36430
rect 80556 35700 80612 37548
rect 80556 35634 80612 35644
rect 80780 35588 80836 39200
rect 80892 36820 80948 36830
rect 80892 36594 80948 36764
rect 80892 36542 80894 36594
rect 80946 36542 80948 36594
rect 80892 36530 80948 36542
rect 81340 35700 81396 35710
rect 80780 35522 80836 35532
rect 81228 35644 81340 35700
rect 80668 34692 80724 34702
rect 80668 34598 80724 34636
rect 81228 34356 81284 35644
rect 81340 35606 81396 35644
rect 81676 35028 81732 39200
rect 82012 38500 82068 38510
rect 82012 36484 82068 38444
rect 82012 36482 82180 36484
rect 82012 36430 82014 36482
rect 82066 36430 82180 36482
rect 82012 36428 82180 36430
rect 82012 36418 82068 36428
rect 82012 35588 82068 35598
rect 82012 35494 82068 35532
rect 81676 34962 81732 34972
rect 81900 34914 81956 34926
rect 81900 34862 81902 34914
rect 81954 34862 81956 34914
rect 81340 34692 81396 34702
rect 81900 34692 81956 34862
rect 82124 34692 82180 36428
rect 82572 35812 82628 39200
rect 83468 36820 83524 39200
rect 84364 39060 84420 39200
rect 84700 39060 84756 39228
rect 84364 39004 84756 39060
rect 83468 36754 83524 36764
rect 84812 36820 84868 36830
rect 81340 34690 81956 34692
rect 81340 34638 81342 34690
rect 81394 34638 81956 34690
rect 81340 34636 81956 34638
rect 82012 34636 82180 34692
rect 82348 35756 82628 35812
rect 82684 36594 82740 36606
rect 82684 36542 82686 36594
rect 82738 36542 82740 36594
rect 81340 34626 81396 34636
rect 81340 34356 81396 34366
rect 81228 34354 81396 34356
rect 81228 34302 81342 34354
rect 81394 34302 81396 34354
rect 81228 34300 81396 34302
rect 81340 34290 81396 34300
rect 80444 34178 80500 34188
rect 81452 30996 81508 34636
rect 81788 34356 81844 34366
rect 82012 34356 82068 34636
rect 81788 34354 82068 34356
rect 81788 34302 81790 34354
rect 81842 34302 82068 34354
rect 81788 34300 82068 34302
rect 82348 34354 82404 35756
rect 82684 35252 82740 36542
rect 84812 36594 84868 36764
rect 84812 36542 84814 36594
rect 84866 36542 84868 36594
rect 84812 36530 84868 36542
rect 84140 36484 84196 36494
rect 84028 36482 84196 36484
rect 84028 36430 84142 36482
rect 84194 36430 84196 36482
rect 84028 36428 84196 36430
rect 83468 35812 83524 35822
rect 83468 35718 83524 35756
rect 83244 35698 83300 35710
rect 83244 35646 83246 35698
rect 83298 35646 83300 35698
rect 83244 35588 83300 35646
rect 83916 35588 83972 35598
rect 83244 35586 83972 35588
rect 83244 35534 83918 35586
rect 83970 35534 83972 35586
rect 83244 35532 83972 35534
rect 82684 35186 82740 35196
rect 82572 35028 82628 35038
rect 82572 34934 82628 34972
rect 82348 34302 82350 34354
rect 82402 34302 82404 34354
rect 81788 34290 81844 34300
rect 82348 34244 82404 34302
rect 83692 34690 83748 34702
rect 83692 34638 83694 34690
rect 83746 34638 83748 34690
rect 82348 34178 82404 34188
rect 82796 34242 82852 34254
rect 82796 34190 82798 34242
rect 82850 34190 82852 34242
rect 81452 30930 81508 30940
rect 82796 25732 82852 34190
rect 83132 34244 83188 34254
rect 83132 34150 83188 34188
rect 83692 33572 83748 34638
rect 83692 33506 83748 33516
rect 83804 26516 83860 35532
rect 83916 35522 83972 35532
rect 84028 35308 84084 36428
rect 84140 36418 84196 36428
rect 84588 35700 84644 35710
rect 83916 35252 84084 35308
rect 84364 35698 84644 35700
rect 84364 35646 84590 35698
rect 84642 35646 84644 35698
rect 84364 35644 84644 35646
rect 83916 34354 83972 35252
rect 84028 34802 84084 34814
rect 84028 34750 84030 34802
rect 84082 34750 84084 34802
rect 84028 34468 84084 34750
rect 84028 34402 84084 34412
rect 83916 34302 83918 34354
rect 83970 34302 83972 34354
rect 83916 29316 83972 34302
rect 83916 29250 83972 29260
rect 84364 34354 84420 35644
rect 84588 35634 84644 35644
rect 85036 35588 85092 39228
rect 85232 39200 85344 40000
rect 86128 39200 86240 40000
rect 87024 39200 87136 40000
rect 87920 39200 88032 40000
rect 88816 39200 88928 40000
rect 89712 39200 89824 40000
rect 90608 39200 90720 40000
rect 91504 39200 91616 40000
rect 92400 39200 92512 40000
rect 93296 39200 93408 40000
rect 94192 39200 94304 40000
rect 95088 39200 95200 40000
rect 95984 39200 96096 40000
rect 96880 39200 96992 40000
rect 97776 39200 97888 40000
rect 98140 39228 98532 39284
rect 85260 36820 85316 39200
rect 86156 37044 86212 39200
rect 86940 37380 86996 37390
rect 86156 36988 86660 37044
rect 85260 36754 85316 36764
rect 86156 36820 86212 36830
rect 86156 36594 86212 36764
rect 86156 36542 86158 36594
rect 86210 36542 86212 36594
rect 86156 36530 86212 36542
rect 85260 35588 85316 35598
rect 85036 35586 85316 35588
rect 85036 35534 85262 35586
rect 85314 35534 85316 35586
rect 85036 35532 85316 35534
rect 85260 35522 85316 35532
rect 85260 34916 85316 34926
rect 85260 34802 85316 34860
rect 85260 34750 85262 34802
rect 85314 34750 85316 34802
rect 85260 34738 85316 34750
rect 85596 34802 85652 34814
rect 85596 34750 85598 34802
rect 85650 34750 85652 34802
rect 84364 34302 84366 34354
rect 84418 34302 84420 34354
rect 84364 29204 84420 34302
rect 84364 29138 84420 29148
rect 84588 34690 84644 34702
rect 84588 34638 84590 34690
rect 84642 34638 84644 34690
rect 84588 34468 84644 34638
rect 85596 34692 85652 34750
rect 86156 34692 86212 34702
rect 85596 34690 86212 34692
rect 85596 34638 86158 34690
rect 86210 34638 86212 34690
rect 85596 34636 86212 34638
rect 83804 26450 83860 26460
rect 82796 25666 82852 25676
rect 83132 26068 83188 26078
rect 80108 14242 80164 14252
rect 81452 24500 81508 24510
rect 81452 12740 81508 24444
rect 81452 8428 81508 12684
rect 81452 8372 82404 8428
rect 78428 7646 78430 7698
rect 78482 7646 78484 7698
rect 78428 7476 78484 7646
rect 78428 7410 78484 7420
rect 78540 6804 78596 6814
rect 78540 6690 78596 6748
rect 78540 6638 78542 6690
rect 78594 6638 78596 6690
rect 78540 6626 78596 6638
rect 79100 6468 79156 6478
rect 79100 6374 79156 6412
rect 80892 6468 80948 6478
rect 79884 6020 79940 6030
rect 79884 5926 79940 5964
rect 78764 5908 78820 5918
rect 78764 5814 78820 5852
rect 79436 5908 79492 5918
rect 79436 5814 79492 5852
rect 80444 5908 80500 5918
rect 79996 5796 80052 5806
rect 79884 5794 80052 5796
rect 79884 5742 79998 5794
rect 80050 5742 80052 5794
rect 79884 5740 80052 5742
rect 78988 5236 79044 5246
rect 78428 5124 78484 5134
rect 78428 4450 78484 5068
rect 78428 4398 78430 4450
rect 78482 4398 78484 4450
rect 78428 4386 78484 4398
rect 78988 3666 79044 5180
rect 79884 4452 79940 5740
rect 79996 5730 80052 5740
rect 80444 5794 80500 5852
rect 80444 5742 80446 5794
rect 80498 5742 80500 5794
rect 80444 5124 80500 5742
rect 80892 5346 80948 6412
rect 80892 5294 80894 5346
rect 80946 5294 80948 5346
rect 80892 5282 80948 5294
rect 81340 5794 81396 5806
rect 81340 5742 81342 5794
rect 81394 5742 81396 5794
rect 80444 5058 80500 5068
rect 81340 5012 81396 5742
rect 80108 4898 80164 4910
rect 80108 4846 80110 4898
rect 80162 4846 80164 4898
rect 79996 4564 80052 4574
rect 80108 4564 80164 4846
rect 79996 4562 80164 4564
rect 79996 4510 79998 4562
rect 80050 4510 80164 4562
rect 79996 4508 80164 4510
rect 79996 4498 80052 4508
rect 79884 4358 79940 4396
rect 80444 4452 80500 4462
rect 80444 4358 80500 4396
rect 81340 4452 81396 4956
rect 81340 4386 81396 4396
rect 79100 4340 79156 4350
rect 79100 4246 79156 4284
rect 78988 3614 78990 3666
rect 79042 3614 79044 3666
rect 78988 3602 79044 3614
rect 81788 4226 81844 4238
rect 81788 4174 81790 4226
rect 81842 4174 81844 4226
rect 81452 3556 81508 3566
rect 81452 3462 81508 3500
rect 78428 3444 78484 3454
rect 78428 3350 78484 3388
rect 79324 3444 79380 3454
rect 79324 3350 79380 3388
rect 79660 3444 79716 3454
rect 78092 3330 78260 3332
rect 78092 3278 78094 3330
rect 78146 3278 78260 3330
rect 78092 3276 78260 3278
rect 78092 3266 78148 3276
rect 78204 3220 78260 3276
rect 78204 3154 78260 3164
rect 79660 800 79716 3388
rect 80556 3444 80612 3454
rect 80556 3350 80612 3388
rect 81004 3444 81060 3454
rect 81004 800 81060 3388
rect 81788 3444 81844 4174
rect 81788 3378 81844 3388
rect 82012 3444 82068 3454
rect 82012 3350 82068 3388
rect 82348 3442 82404 8372
rect 82908 8148 82964 8158
rect 82908 3556 82964 8092
rect 82908 3462 82964 3500
rect 82348 3390 82350 3442
rect 82402 3390 82404 3442
rect 82348 3378 82404 3390
rect 83132 3220 83188 26012
rect 84588 6132 84644 34412
rect 86044 34244 86100 34636
rect 86156 34626 86212 34636
rect 86156 34356 86212 34366
rect 86268 34356 86324 36988
rect 86156 34354 86324 34356
rect 86156 34302 86158 34354
rect 86210 34302 86324 34354
rect 86156 34300 86324 34302
rect 86380 35810 86436 35822
rect 86380 35758 86382 35810
rect 86434 35758 86436 35810
rect 86156 34290 86212 34300
rect 86044 34178 86100 34188
rect 86380 26404 86436 35758
rect 86604 35698 86660 36988
rect 86940 36484 86996 37324
rect 86940 36352 86996 36428
rect 86604 35646 86606 35698
rect 86658 35646 86660 35698
rect 86604 35634 86660 35646
rect 87052 35588 87108 39200
rect 87052 35522 87108 35532
rect 87276 37156 87332 37166
rect 86940 34802 86996 34814
rect 86940 34750 86942 34802
rect 86994 34750 86996 34802
rect 86380 26338 86436 26348
rect 86604 34020 86660 34030
rect 86940 34020 86996 34750
rect 87276 34802 87332 37100
rect 87948 36820 88004 39200
rect 88172 38388 88228 38398
rect 87948 36764 88116 36820
rect 87948 36484 88004 36494
rect 87948 36390 88004 36428
rect 87388 35812 87444 35822
rect 87388 35698 87444 35756
rect 87388 35646 87390 35698
rect 87442 35646 87444 35698
rect 87388 35634 87444 35646
rect 87948 35588 88004 35598
rect 87948 35494 88004 35532
rect 88060 35140 88116 36764
rect 88060 35074 88116 35084
rect 88172 34916 88228 38332
rect 88844 37156 88900 39200
rect 88732 37100 88900 37156
rect 89068 37604 89124 37614
rect 87276 34750 87278 34802
rect 87330 34750 87332 34802
rect 87276 34738 87332 34750
rect 88060 34914 88228 34916
rect 88060 34862 88174 34914
rect 88226 34862 88228 34914
rect 88060 34860 88228 34862
rect 87388 34580 87444 34590
rect 87388 34354 87444 34524
rect 87388 34302 87390 34354
rect 87442 34302 87444 34354
rect 87388 34290 87444 34302
rect 87948 34580 88004 34590
rect 87948 34354 88004 34524
rect 87948 34302 87950 34354
rect 88002 34302 88004 34354
rect 87948 34290 88004 34302
rect 86604 34018 86996 34020
rect 86604 33966 86606 34018
rect 86658 33966 86996 34018
rect 86604 33964 86996 33966
rect 86604 21028 86660 33964
rect 87948 33460 88004 33470
rect 88060 33460 88116 34860
rect 88172 34850 88228 34860
rect 88620 36258 88676 36270
rect 88620 36206 88622 36258
rect 88674 36206 88676 36258
rect 88508 34018 88564 34030
rect 88508 33966 88510 34018
rect 88562 33966 88564 34018
rect 88508 33572 88564 33966
rect 88508 33506 88564 33516
rect 87948 33458 88116 33460
rect 87948 33406 87950 33458
rect 88002 33406 88116 33458
rect 87948 33404 88116 33406
rect 87948 33394 88004 33404
rect 88620 31948 88676 36206
rect 88732 35028 88788 37100
rect 89068 36932 89124 37548
rect 89740 37268 89796 39200
rect 89068 36866 89124 36876
rect 89628 37212 89796 37268
rect 88956 36484 89012 36494
rect 88956 36390 89012 36428
rect 89516 36370 89572 36382
rect 89516 36318 89518 36370
rect 89570 36318 89572 36370
rect 89516 36260 89572 36318
rect 89516 36194 89572 36204
rect 89404 35810 89460 35822
rect 89404 35758 89406 35810
rect 89458 35758 89460 35810
rect 88732 34962 88788 34972
rect 88844 35140 88900 35150
rect 88844 35026 88900 35084
rect 88844 34974 88846 35026
rect 88898 34974 88900 35026
rect 88844 34962 88900 34974
rect 89292 34580 89348 34590
rect 89292 34354 89348 34524
rect 89292 34302 89294 34354
rect 89346 34302 89348 34354
rect 89068 33460 89124 33470
rect 89292 33460 89348 34302
rect 89404 34020 89460 35758
rect 89628 35140 89684 37212
rect 89740 36484 89796 36494
rect 89740 36482 90020 36484
rect 89740 36430 89742 36482
rect 89794 36430 90020 36482
rect 89740 36428 90020 36430
rect 89740 36418 89796 36428
rect 89628 35074 89684 35084
rect 89740 36260 89796 36270
rect 89404 33964 89572 34020
rect 89068 33458 89348 33460
rect 89068 33406 89070 33458
rect 89122 33406 89348 33458
rect 89068 33404 89348 33406
rect 89404 33684 89460 33694
rect 89068 33394 89124 33404
rect 86604 20962 86660 20972
rect 87612 31892 88676 31948
rect 87612 20188 87668 31892
rect 87612 20132 87780 20188
rect 85820 17668 85876 17678
rect 85820 11732 85876 17612
rect 85484 8036 85540 8046
rect 85484 7698 85540 7980
rect 85484 7646 85486 7698
rect 85538 7646 85540 7698
rect 85484 7634 85540 7646
rect 84588 6066 84644 6076
rect 85260 5010 85316 5022
rect 85260 4958 85262 5010
rect 85314 4958 85316 5010
rect 84476 4898 84532 4910
rect 84476 4846 84478 4898
rect 84530 4846 84532 4898
rect 84476 4564 84532 4846
rect 84476 4498 84532 4508
rect 85260 4564 85316 4958
rect 85596 5012 85652 5022
rect 85596 4918 85652 4956
rect 85260 4498 85316 4508
rect 85372 3668 85428 3678
rect 85372 3554 85428 3612
rect 85372 3502 85374 3554
rect 85426 3502 85428 3554
rect 85372 3490 85428 3502
rect 83132 3154 83188 3164
rect 83692 3444 83748 3454
rect 83692 800 83748 3388
rect 84476 3444 84532 3454
rect 84476 3350 84532 3388
rect 85036 3444 85092 3454
rect 85036 800 85092 3388
rect 85820 3332 85876 11676
rect 86044 8036 86100 8046
rect 86604 8036 86660 8046
rect 87052 8036 87108 8046
rect 87612 8036 87668 8046
rect 86044 7698 86100 7980
rect 86044 7646 86046 7698
rect 86098 7646 86100 7698
rect 86044 7634 86100 7646
rect 86492 8034 87108 8036
rect 86492 7982 86606 8034
rect 86658 7982 87054 8034
rect 87106 7982 87108 8034
rect 86492 7980 87108 7982
rect 86268 7476 86324 7486
rect 85932 5124 85988 5134
rect 85932 4562 85988 5068
rect 85932 4510 85934 4562
rect 85986 4510 85988 4562
rect 85932 4498 85988 4510
rect 86268 4564 86324 7420
rect 86492 7362 86548 7980
rect 86604 7970 86660 7980
rect 87052 7588 87108 7980
rect 87052 7522 87108 7532
rect 87500 8034 87668 8036
rect 87500 7982 87614 8034
rect 87666 7982 87668 8034
rect 87500 7980 87668 7982
rect 86492 7310 86494 7362
rect 86546 7310 86548 7362
rect 86492 7140 86548 7310
rect 87276 7252 87332 7262
rect 86492 7074 86548 7084
rect 86716 7250 87332 7252
rect 86716 7198 87278 7250
rect 87330 7198 87332 7250
rect 86716 7196 87332 7198
rect 86380 6692 86436 6702
rect 86716 6692 86772 7196
rect 87276 7186 87332 7196
rect 86380 6690 86772 6692
rect 86380 6638 86382 6690
rect 86434 6638 86772 6690
rect 86380 6636 86772 6638
rect 87052 6692 87108 6702
rect 86380 6626 86436 6636
rect 86604 6468 86660 6478
rect 86604 6466 86772 6468
rect 86604 6414 86606 6466
rect 86658 6414 86772 6466
rect 86604 6412 86772 6414
rect 86604 6402 86660 6412
rect 86380 5124 86436 5134
rect 86380 5030 86436 5068
rect 86716 5122 86772 6412
rect 86828 5796 86884 5806
rect 87052 5796 87108 6636
rect 87500 6018 87556 7980
rect 87612 7970 87668 7980
rect 87724 7700 87780 20132
rect 89068 11284 89124 11294
rect 87948 8260 88004 8270
rect 87948 8166 88004 8204
rect 87612 7476 87668 7486
rect 87724 7476 87780 7644
rect 88284 8146 88340 8158
rect 88284 8094 88286 8146
rect 88338 8094 88340 8146
rect 87836 7588 87892 7598
rect 87836 7494 87892 7532
rect 88284 7588 88340 8094
rect 88508 8148 88564 8158
rect 88508 8054 88564 8092
rect 88284 7522 88340 7532
rect 88396 7586 88452 7598
rect 88396 7534 88398 7586
rect 88450 7534 88452 7586
rect 87612 7474 87780 7476
rect 87612 7422 87614 7474
rect 87666 7422 87780 7474
rect 87612 7420 87780 7422
rect 87612 7410 87668 7420
rect 88396 7364 88452 7534
rect 88396 7298 88452 7308
rect 87724 6690 87780 6702
rect 87724 6638 87726 6690
rect 87778 6638 87780 6690
rect 87724 6132 87780 6638
rect 87836 6132 87892 6142
rect 87724 6130 87892 6132
rect 87724 6078 87838 6130
rect 87890 6078 87892 6130
rect 87724 6076 87892 6078
rect 87836 6066 87892 6076
rect 87500 5966 87502 6018
rect 87554 5966 87556 6018
rect 87500 5954 87556 5966
rect 86828 5794 87108 5796
rect 86828 5742 86830 5794
rect 86882 5742 87108 5794
rect 86828 5740 87108 5742
rect 86828 5236 86884 5740
rect 86828 5170 86884 5180
rect 86716 5070 86718 5122
rect 86770 5070 86772 5122
rect 86716 5058 86772 5070
rect 86380 4564 86436 4574
rect 86268 4562 86436 4564
rect 86268 4510 86382 4562
rect 86434 4510 86436 4562
rect 86268 4508 86436 4510
rect 86268 3668 86324 4508
rect 86380 4498 86436 4508
rect 88508 4564 88564 4574
rect 88508 4470 88564 4508
rect 86268 3602 86324 3612
rect 86268 3444 86324 3454
rect 86268 3350 86324 3388
rect 86716 3444 86772 3454
rect 86716 3350 86772 3388
rect 87724 3444 87780 3454
rect 85932 3332 85988 3342
rect 85820 3330 85988 3332
rect 85820 3278 85934 3330
rect 85986 3278 85988 3330
rect 85820 3276 85988 3278
rect 85932 3266 85988 3276
rect 87724 800 87780 3388
rect 88396 3444 88452 3454
rect 88396 3350 88452 3388
rect 89068 3332 89124 11228
rect 89404 8260 89460 33628
rect 89516 33236 89572 33964
rect 89516 33142 89572 33180
rect 89740 31948 89796 36204
rect 89964 35812 90020 36428
rect 89852 34244 89908 34254
rect 89964 34244 90020 35756
rect 90412 36258 90468 36270
rect 90412 36206 90414 36258
rect 90466 36206 90468 36258
rect 90188 35700 90244 35710
rect 90188 35606 90244 35644
rect 90412 35476 90468 36206
rect 90636 36036 90692 39200
rect 90636 35970 90692 35980
rect 90748 36370 90804 36382
rect 90748 36318 90750 36370
rect 90802 36318 90804 36370
rect 90412 35410 90468 35420
rect 90524 35474 90580 35486
rect 90524 35422 90526 35474
rect 90578 35422 90580 35474
rect 90188 35028 90244 35038
rect 90188 34934 90244 34972
rect 89852 34242 90020 34244
rect 89852 34190 89854 34242
rect 89906 34190 90020 34242
rect 89852 34188 90020 34190
rect 89852 34178 89908 34188
rect 89628 31892 89796 31948
rect 90300 34020 90356 34030
rect 89628 26180 89684 31892
rect 89628 26114 89684 26124
rect 90300 25620 90356 33964
rect 90524 33684 90580 35422
rect 90748 35308 90804 36318
rect 91196 36372 91252 36382
rect 91196 36278 91252 36316
rect 91196 35698 91252 35710
rect 91196 35646 91198 35698
rect 91250 35646 91252 35698
rect 90636 35252 90804 35308
rect 90972 35476 91028 35486
rect 90636 34020 90692 35252
rect 90972 34914 91028 35420
rect 90972 34862 90974 34914
rect 91026 34862 91028 34914
rect 90972 34850 91028 34862
rect 90636 33954 90692 33964
rect 90860 34356 90916 34366
rect 91196 34356 91252 35646
rect 90860 34354 91252 34356
rect 90860 34302 90862 34354
rect 90914 34302 91252 34354
rect 90860 34300 91252 34302
rect 91532 34356 91588 39200
rect 92316 38276 92372 38286
rect 91980 36596 92036 36606
rect 91980 36370 92036 36540
rect 91980 36318 91982 36370
rect 92034 36318 92036 36370
rect 91980 36306 92036 36318
rect 92204 36482 92260 36494
rect 92204 36430 92206 36482
rect 92258 36430 92260 36482
rect 91868 36036 91924 36046
rect 91868 35586 91924 35980
rect 91868 35534 91870 35586
rect 91922 35534 91924 35586
rect 91868 35522 91924 35534
rect 90524 33618 90580 33628
rect 90860 27860 90916 34300
rect 91532 34290 91588 34300
rect 91868 35140 91924 35150
rect 91868 34916 91924 35084
rect 92204 34916 92260 36430
rect 92316 36036 92372 38220
rect 92316 35970 92372 35980
rect 92428 35028 92484 39200
rect 93324 37044 93380 39200
rect 93324 36988 93940 37044
rect 93262 36876 93526 36886
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93262 36810 93526 36820
rect 92988 36484 93044 36494
rect 92764 36260 92820 36270
rect 92764 36166 92820 36204
rect 92988 35922 93044 36428
rect 93660 36482 93716 36494
rect 93660 36430 93662 36482
rect 93714 36430 93716 36482
rect 92988 35870 92990 35922
rect 93042 35870 93044 35922
rect 92988 35700 93044 35870
rect 92988 35634 93044 35644
rect 93100 36148 93156 36158
rect 92428 34962 92484 34972
rect 91868 34860 92260 34916
rect 91756 34132 91812 34142
rect 91196 34130 91812 34132
rect 91196 34078 91758 34130
rect 91810 34078 91812 34130
rect 91196 34076 91812 34078
rect 91196 34018 91252 34076
rect 91756 34066 91812 34076
rect 91196 33966 91198 34018
rect 91250 33966 91252 34018
rect 91196 28868 91252 33966
rect 91756 33460 91812 33470
rect 91868 33460 91924 34860
rect 92428 34802 92484 34814
rect 92428 34750 92430 34802
rect 92482 34750 92484 34802
rect 91756 33458 91924 33460
rect 91756 33406 91758 33458
rect 91810 33406 91924 33458
rect 91756 33404 91924 33406
rect 92092 34690 92148 34702
rect 92092 34638 92094 34690
rect 92146 34638 92148 34690
rect 92092 33460 92148 34638
rect 92428 34580 92484 34750
rect 92428 34514 92484 34524
rect 92652 34356 92708 34366
rect 92652 34242 92708 34300
rect 92652 34190 92654 34242
rect 92706 34190 92708 34242
rect 92652 34178 92708 34190
rect 93100 33460 93156 36092
rect 93660 36036 93716 36430
rect 93772 36370 93828 36382
rect 93772 36318 93774 36370
rect 93826 36318 93828 36370
rect 93772 36148 93828 36318
rect 93772 36082 93828 36092
rect 93548 35980 93716 36036
rect 93548 35812 93604 35980
rect 93548 35698 93604 35756
rect 93548 35646 93550 35698
rect 93602 35646 93604 35698
rect 93548 35634 93604 35646
rect 93660 35810 93716 35822
rect 93660 35758 93662 35810
rect 93714 35758 93716 35810
rect 93262 35308 93526 35318
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93262 35242 93526 35252
rect 93660 35140 93716 35758
rect 93884 35252 93940 36988
rect 94220 36596 94276 39200
rect 94220 36530 94276 36540
rect 94332 36482 94388 36494
rect 94332 36430 94334 36482
rect 94386 36430 94388 36482
rect 94332 36372 94388 36430
rect 94332 36306 94388 36316
rect 94668 36260 94724 36270
rect 94668 36258 95060 36260
rect 94668 36206 94670 36258
rect 94722 36206 95060 36258
rect 94668 36204 95060 36206
rect 94668 36194 94724 36204
rect 94332 35700 94388 35710
rect 94332 35606 94388 35644
rect 93884 35186 93940 35196
rect 94668 35474 94724 35486
rect 94668 35422 94670 35474
rect 94722 35422 94724 35474
rect 93324 35084 93716 35140
rect 93324 34692 93380 35084
rect 93996 35028 94052 35038
rect 93996 34934 94052 34972
rect 93436 34916 93492 34926
rect 93436 34914 93940 34916
rect 93436 34862 93438 34914
rect 93490 34862 93940 34914
rect 93436 34860 93940 34862
rect 93436 34850 93492 34860
rect 93324 34626 93380 34636
rect 93436 34580 93492 34590
rect 93436 34354 93492 34524
rect 93436 34302 93438 34354
rect 93490 34302 93492 34354
rect 93436 34290 93492 34302
rect 93884 34018 93940 34860
rect 93884 33966 93886 34018
rect 93938 33966 93940 34018
rect 93262 33740 93526 33750
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93262 33674 93526 33684
rect 93212 33460 93268 33470
rect 93100 33458 93268 33460
rect 93100 33406 93214 33458
rect 93266 33406 93268 33458
rect 93100 33404 93268 33406
rect 91756 33394 91812 33404
rect 92092 33394 92148 33404
rect 93212 33394 93268 33404
rect 93262 32172 93526 32182
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93262 32106 93526 32116
rect 93262 30604 93526 30614
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93262 30538 93526 30548
rect 93262 29036 93526 29046
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93262 28970 93526 28980
rect 91196 28802 91252 28812
rect 90860 27794 90916 27804
rect 93262 27468 93526 27478
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93262 27402 93526 27412
rect 93884 27300 93940 33966
rect 94668 31948 94724 35422
rect 94668 31892 94836 31948
rect 93884 27234 93940 27244
rect 90300 25554 90356 25564
rect 91532 26180 91588 26190
rect 91532 11732 91588 26124
rect 93262 25900 93526 25910
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93262 25834 93526 25844
rect 93262 24332 93526 24342
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93262 24266 93526 24276
rect 93262 22764 93526 22774
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93262 22698 93526 22708
rect 93262 21196 93526 21206
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93262 21130 93526 21140
rect 93262 19628 93526 19638
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93262 19562 93526 19572
rect 93262 18060 93526 18070
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93262 17994 93526 18004
rect 93262 16492 93526 16502
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93262 16426 93526 16436
rect 93262 14924 93526 14934
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93262 14858 93526 14868
rect 93262 13356 93526 13366
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93262 13290 93526 13300
rect 93262 11788 93526 11798
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93262 11722 93526 11732
rect 91532 11666 91588 11676
rect 93262 10220 93526 10230
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93262 10154 93526 10164
rect 93262 8652 93526 8662
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93262 8586 93526 8596
rect 89404 8166 89460 8204
rect 90748 8260 90804 8270
rect 89852 8148 89908 8158
rect 89852 8054 89908 8092
rect 90076 8148 90132 8158
rect 89180 7700 89236 7710
rect 89180 7606 89236 7644
rect 89628 7364 89684 7374
rect 89684 7308 89796 7364
rect 89628 7232 89684 7308
rect 89404 5794 89460 5806
rect 89404 5742 89406 5794
rect 89458 5742 89460 5794
rect 89292 5682 89348 5694
rect 89292 5630 89294 5682
rect 89346 5630 89348 5682
rect 89292 4898 89348 5630
rect 89404 5012 89460 5742
rect 89404 4946 89460 4956
rect 89628 5684 89684 5694
rect 89292 4846 89294 4898
rect 89346 4846 89348 4898
rect 89292 4834 89348 4846
rect 89292 4564 89348 4574
rect 89292 4450 89348 4508
rect 89628 4562 89684 5628
rect 89740 5124 89796 7308
rect 89964 5794 90020 5806
rect 89964 5742 89966 5794
rect 90018 5742 90020 5794
rect 89852 5124 89908 5134
rect 89740 5122 89908 5124
rect 89740 5070 89854 5122
rect 89906 5070 89908 5122
rect 89740 5068 89908 5070
rect 89628 4510 89630 4562
rect 89682 4510 89684 4562
rect 89628 4498 89684 4510
rect 89292 4398 89294 4450
rect 89346 4398 89348 4450
rect 89292 4386 89348 4398
rect 89852 3780 89908 5068
rect 89964 5012 90020 5742
rect 89964 4946 90020 4956
rect 89852 3714 89908 3724
rect 90076 4562 90132 8092
rect 90748 6690 90804 8204
rect 94780 8260 94836 31892
rect 95004 20188 95060 36204
rect 95116 35140 95172 39200
rect 95900 36372 95956 36382
rect 95340 35812 95396 35822
rect 95340 35810 95508 35812
rect 95340 35758 95342 35810
rect 95394 35758 95508 35810
rect 95340 35756 95508 35758
rect 95340 35746 95396 35756
rect 95116 35074 95172 35084
rect 95340 34916 95396 34926
rect 95116 34914 95396 34916
rect 95116 34862 95342 34914
rect 95394 34862 95396 34914
rect 95116 34860 95396 34862
rect 95116 34018 95172 34860
rect 95340 34850 95396 34860
rect 95116 33966 95118 34018
rect 95170 33966 95172 34018
rect 95116 28420 95172 33966
rect 95452 33908 95508 35756
rect 95564 35698 95620 35710
rect 95564 35646 95566 35698
rect 95618 35646 95620 35698
rect 95564 35252 95620 35646
rect 95564 34354 95620 35196
rect 95564 34302 95566 34354
rect 95618 34302 95620 34354
rect 95564 34290 95620 34302
rect 95900 34020 95956 36316
rect 96012 35308 96068 39200
rect 96572 36596 96628 36606
rect 96572 36502 96628 36540
rect 96908 36596 96964 39200
rect 97804 39060 97860 39200
rect 98140 39060 98196 39228
rect 97804 39004 98196 39060
rect 96908 36530 96964 36540
rect 97244 36932 97300 36942
rect 96124 36484 96180 36494
rect 96124 36482 96404 36484
rect 96124 36430 96126 36482
rect 96178 36430 96404 36482
rect 96124 36428 96404 36430
rect 96124 36418 96180 36428
rect 96124 35588 96180 35598
rect 96124 35586 96292 35588
rect 96124 35534 96126 35586
rect 96178 35534 96292 35586
rect 96124 35532 96292 35534
rect 96124 35522 96180 35532
rect 96012 35252 96180 35308
rect 96012 35140 96068 35150
rect 96012 35026 96068 35084
rect 96012 34974 96014 35026
rect 96066 34974 96068 35026
rect 96012 34962 96068 34974
rect 96124 35028 96180 35252
rect 96124 34962 96180 34972
rect 96236 34692 96292 35532
rect 96236 34626 96292 34636
rect 96348 34354 96404 36428
rect 97244 35922 97300 36876
rect 98364 36596 98420 36606
rect 98364 36502 98420 36540
rect 97916 36484 97972 36494
rect 97916 36482 98308 36484
rect 97916 36430 97918 36482
rect 97970 36430 98308 36482
rect 97916 36428 98308 36430
rect 97916 36418 97972 36428
rect 97244 35870 97246 35922
rect 97298 35870 97300 35922
rect 97244 35700 97300 35870
rect 97244 35634 97300 35644
rect 98028 35698 98084 35710
rect 98028 35646 98030 35698
rect 98082 35646 98084 35698
rect 97356 35028 97412 35038
rect 97356 34914 97412 34972
rect 97356 34862 97358 34914
rect 97410 34862 97412 34914
rect 96348 34302 96350 34354
rect 96402 34302 96404 34354
rect 96012 34020 96068 34030
rect 95900 34018 96068 34020
rect 95900 33966 96014 34018
rect 96066 33966 96068 34018
rect 95900 33964 96068 33966
rect 95452 33842 95508 33852
rect 96012 33236 96068 33964
rect 96012 33170 96068 33180
rect 96348 31220 96404 34302
rect 96348 31154 96404 31164
rect 97132 34690 97188 34702
rect 97132 34638 97134 34690
rect 97186 34638 97188 34690
rect 95116 28354 95172 28364
rect 96572 27748 96628 27758
rect 95004 20132 95172 20188
rect 94780 8166 94836 8204
rect 93772 8148 93828 8158
rect 92540 8036 92596 8046
rect 92540 7698 92596 7980
rect 92540 7646 92542 7698
rect 92594 7646 92596 7698
rect 92540 7634 92596 7646
rect 93100 8036 93156 8046
rect 93100 7698 93156 7980
rect 93100 7646 93102 7698
rect 93154 7646 93156 7698
rect 93100 7634 93156 7646
rect 93660 7588 93716 7598
rect 93772 7588 93828 8092
rect 94892 8148 94948 8158
rect 94444 8036 94500 8046
rect 94444 8034 94612 8036
rect 94444 7982 94446 8034
rect 94498 7982 94612 8034
rect 94444 7980 94612 7982
rect 94444 7970 94500 7980
rect 93660 7586 94052 7588
rect 93660 7534 93662 7586
rect 93714 7534 94052 7586
rect 93660 7532 94052 7534
rect 93660 7522 93716 7532
rect 93262 7084 93526 7094
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93262 7018 93526 7028
rect 93996 6802 94052 7532
rect 94444 7586 94500 7598
rect 94444 7534 94446 7586
rect 94498 7534 94500 7586
rect 94444 7476 94500 7534
rect 94444 7410 94500 7420
rect 93996 6750 93998 6802
rect 94050 6750 94052 6802
rect 93996 6738 94052 6750
rect 90748 6638 90750 6690
rect 90802 6638 90804 6690
rect 90748 6626 90804 6638
rect 94556 6690 94612 7980
rect 94892 7586 94948 8092
rect 94892 7534 94894 7586
rect 94946 7534 94948 7586
rect 94892 7522 94948 7534
rect 95116 7700 95172 20132
rect 95564 8258 95620 8270
rect 95564 8206 95566 8258
rect 95618 8206 95620 8258
rect 95340 8146 95396 8158
rect 95340 8094 95342 8146
rect 95394 8094 95396 8146
rect 95340 8036 95396 8094
rect 95564 8148 95620 8206
rect 96124 8260 96180 8270
rect 96124 8166 96180 8204
rect 95564 8082 95620 8092
rect 95340 7970 95396 7980
rect 95116 7474 95172 7644
rect 96012 7700 96068 7710
rect 96012 7606 96068 7644
rect 95116 7422 95118 7474
rect 95170 7422 95172 7474
rect 95116 7410 95172 7422
rect 96460 7476 96516 7486
rect 96460 7382 96516 7420
rect 95452 7252 95508 7262
rect 94556 6638 94558 6690
rect 94610 6638 94612 6690
rect 94556 6626 94612 6638
rect 95228 7250 95508 7252
rect 95228 7198 95454 7250
rect 95506 7198 95508 7250
rect 95228 7196 95508 7198
rect 90188 6466 90244 6478
rect 90188 6414 90190 6466
rect 90242 6414 90244 6466
rect 90188 5348 90244 6414
rect 94780 6468 94836 6478
rect 94780 6466 94948 6468
rect 94780 6414 94782 6466
rect 94834 6414 94948 6466
rect 94780 6412 94948 6414
rect 94780 6402 94836 6412
rect 93262 5516 93526 5526
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93262 5450 93526 5460
rect 90300 5348 90356 5358
rect 90188 5346 90356 5348
rect 90188 5294 90302 5346
rect 90354 5294 90356 5346
rect 90188 5292 90356 5294
rect 90300 5282 90356 5292
rect 90412 5122 90468 5134
rect 90412 5070 90414 5122
rect 90466 5070 90468 5122
rect 90412 5012 90468 5070
rect 93884 5124 93940 5134
rect 93884 5030 93940 5068
rect 94556 5124 94612 5134
rect 94556 5030 94612 5068
rect 94892 5122 94948 6412
rect 95116 5908 95172 5918
rect 95228 5908 95284 7196
rect 95452 7186 95508 7196
rect 95452 6692 95508 6702
rect 95452 6598 95508 6636
rect 95676 6692 95732 6702
rect 95340 6468 95396 6478
rect 95340 6130 95396 6412
rect 95340 6078 95342 6130
rect 95394 6078 95396 6130
rect 95340 6066 95396 6078
rect 95564 6132 95620 6142
rect 95676 6132 95732 6636
rect 95788 6690 95844 6702
rect 95788 6638 95790 6690
rect 95842 6638 95844 6690
rect 95788 6468 95844 6638
rect 95788 6402 95844 6412
rect 95788 6132 95844 6142
rect 95676 6130 95844 6132
rect 95676 6078 95790 6130
rect 95842 6078 95844 6130
rect 95676 6076 95844 6078
rect 95116 5906 95284 5908
rect 95116 5854 95118 5906
rect 95170 5854 95284 5906
rect 95116 5852 95284 5854
rect 95116 5842 95172 5852
rect 94892 5070 94894 5122
rect 94946 5070 94948 5122
rect 94892 5058 94948 5070
rect 90412 4946 90468 4956
rect 90860 4900 90916 4910
rect 90860 4806 90916 4844
rect 90076 4510 90078 4562
rect 90130 4510 90132 4562
rect 89292 3556 89348 3566
rect 90076 3556 90132 4510
rect 93548 4228 93604 4238
rect 93548 4226 93716 4228
rect 93548 4174 93550 4226
rect 93602 4174 93716 4226
rect 93548 4172 93716 4174
rect 93548 4162 93604 4172
rect 93262 3948 93526 3958
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93262 3882 93526 3892
rect 89292 3554 90132 3556
rect 89292 3502 89294 3554
rect 89346 3502 90132 3554
rect 89292 3500 90132 3502
rect 93212 3668 93268 3678
rect 93212 3554 93268 3612
rect 93212 3502 93214 3554
rect 93266 3502 93268 3554
rect 89292 3490 89348 3500
rect 93212 3490 93268 3502
rect 89068 3266 89124 3276
rect 89180 3444 89236 3454
rect 89180 2548 89236 3388
rect 90188 3444 90244 3454
rect 90188 3350 90244 3388
rect 90636 3444 90692 3454
rect 90636 3350 90692 3388
rect 91756 3444 91812 3454
rect 89068 2492 89236 2548
rect 89852 3332 89908 3342
rect 89852 2548 89908 3276
rect 89068 800 89124 2492
rect 89852 2482 89908 2492
rect 91756 800 91812 3388
rect 92316 3444 92372 3454
rect 92316 3350 92372 3388
rect 93100 3444 93156 3454
rect 93660 3444 93716 4172
rect 94668 3668 94724 3678
rect 94668 3574 94724 3612
rect 93772 3444 93828 3454
rect 93660 3388 93772 3444
rect 93100 800 93156 3388
rect 93772 3350 93828 3388
rect 94108 3330 94164 3342
rect 94108 3278 94110 3330
rect 94162 3278 94164 3330
rect 94108 3220 94164 3278
rect 95564 3332 95620 6076
rect 95788 6066 95844 6076
rect 96572 6020 96628 27692
rect 97132 27188 97188 34638
rect 97244 34356 97300 34366
rect 97356 34356 97412 34862
rect 97244 34354 97412 34356
rect 97244 34302 97246 34354
rect 97298 34302 97412 34354
rect 97244 34300 97412 34302
rect 98028 34690 98084 35646
rect 98028 34638 98030 34690
rect 98082 34638 98084 34690
rect 97244 34290 97300 34300
rect 97132 27122 97188 27132
rect 98028 26292 98084 34638
rect 98252 34692 98308 36428
rect 98476 35588 98532 39228
rect 98672 39200 98784 40000
rect 99568 39200 99680 40000
rect 100464 39200 100576 40000
rect 101360 39200 101472 40000
rect 102256 39200 102368 40000
rect 103152 39200 103264 40000
rect 104048 39200 104160 40000
rect 104944 39200 105056 40000
rect 105840 39200 105952 40000
rect 106736 39200 106848 40000
rect 107100 39228 107492 39284
rect 98700 35812 98756 39200
rect 99596 37828 99652 39200
rect 99596 37772 100100 37828
rect 100044 36594 100100 37772
rect 100044 36542 100046 36594
rect 100098 36542 100100 36594
rect 100044 36530 100100 36542
rect 100492 36596 100548 39200
rect 100492 36530 100548 36540
rect 101052 36708 101108 36718
rect 100828 36484 100884 36494
rect 100604 36482 100884 36484
rect 100604 36430 100830 36482
rect 100882 36430 100884 36482
rect 100604 36428 100884 36430
rect 100604 36036 100660 36428
rect 100828 36418 100884 36428
rect 99820 35924 99876 35934
rect 99820 35830 99876 35868
rect 100604 35922 100660 35980
rect 100604 35870 100606 35922
rect 100658 35870 100660 35922
rect 100604 35858 100660 35870
rect 101052 35812 101108 36652
rect 101388 36708 101444 39200
rect 102172 37044 102228 37054
rect 101388 36652 101892 36708
rect 101164 35924 101220 35934
rect 101388 35924 101444 36652
rect 101612 36484 101668 36494
rect 101164 35922 101444 35924
rect 101164 35870 101166 35922
rect 101218 35870 101444 35922
rect 101164 35868 101444 35870
rect 101500 36482 101668 36484
rect 101500 36430 101614 36482
rect 101666 36430 101668 36482
rect 101500 36428 101668 36430
rect 101164 35858 101220 35868
rect 98700 35756 98868 35812
rect 98700 35588 98756 35598
rect 98476 35586 98756 35588
rect 98476 35534 98702 35586
rect 98754 35534 98756 35586
rect 98476 35532 98756 35534
rect 98700 35522 98756 35532
rect 98812 35252 98868 35756
rect 101052 35746 101108 35756
rect 100044 35698 100100 35710
rect 100044 35646 100046 35698
rect 100098 35646 100100 35698
rect 98812 35186 98868 35196
rect 99596 35252 99652 35262
rect 99596 35026 99652 35196
rect 100044 35252 100100 35646
rect 100044 35186 100100 35196
rect 99596 34974 99598 35026
rect 99650 34974 99652 35026
rect 99596 34962 99652 34974
rect 98364 34692 98420 34702
rect 98252 34690 98420 34692
rect 98252 34638 98366 34690
rect 98418 34638 98420 34690
rect 98252 34636 98420 34638
rect 98364 29652 98420 34636
rect 98364 29586 98420 29596
rect 99932 34692 99988 34702
rect 98028 26226 98084 26236
rect 98140 19348 98196 19358
rect 98140 11844 98196 19292
rect 96684 8036 96740 8046
rect 96684 7942 96740 7980
rect 98028 8036 98084 8046
rect 96460 5964 96628 6020
rect 95564 3266 95620 3276
rect 95788 3444 95844 3454
rect 94108 2660 94164 3164
rect 94108 2594 94164 2604
rect 95788 800 95844 3388
rect 96348 3444 96404 3454
rect 96348 3350 96404 3388
rect 96460 3220 96516 5964
rect 96572 5794 96628 5806
rect 96572 5742 96574 5794
rect 96626 5742 96628 5794
rect 96572 5684 96628 5742
rect 96572 5618 96628 5628
rect 97244 5794 97300 5806
rect 97244 5742 97246 5794
rect 97298 5742 97300 5794
rect 97244 5684 97300 5742
rect 97244 5618 97300 5628
rect 97356 5682 97412 5694
rect 97356 5630 97358 5682
rect 97410 5630 97412 5682
rect 97356 4898 97412 5630
rect 98028 5346 98084 7980
rect 98028 5294 98030 5346
rect 98082 5294 98084 5346
rect 98028 5282 98084 5294
rect 97356 4846 97358 4898
rect 97410 4846 97412 4898
rect 97356 4834 97412 4846
rect 97580 4226 97636 4238
rect 97580 4174 97582 4226
rect 97634 4174 97636 4226
rect 97244 3556 97300 3566
rect 97244 3462 97300 3500
rect 96460 3154 96516 3164
rect 97132 3444 97188 3454
rect 97132 800 97188 3388
rect 97580 3444 97636 4174
rect 97580 3378 97636 3388
rect 97804 3444 97860 3454
rect 97804 3350 97860 3388
rect 98140 3330 98196 11788
rect 98924 7476 98980 7486
rect 98924 6690 98980 7420
rect 98924 6638 98926 6690
rect 98978 6638 98980 6690
rect 98924 6626 98980 6638
rect 98252 6466 98308 6478
rect 98252 6414 98254 6466
rect 98306 6414 98308 6466
rect 98252 6130 98308 6414
rect 98252 6078 98254 6130
rect 98306 6078 98308 6130
rect 98252 6066 98308 6078
rect 98364 5794 98420 5806
rect 98364 5742 98366 5794
rect 98418 5742 98420 5794
rect 98364 5684 98420 5742
rect 98364 5618 98420 5628
rect 98924 5794 98980 5806
rect 98924 5742 98926 5794
rect 98978 5742 98980 5794
rect 98924 5684 98980 5742
rect 98924 5618 98980 5628
rect 98700 3556 98756 3566
rect 98700 3462 98756 3500
rect 98140 3278 98142 3330
rect 98194 3278 98196 3330
rect 98140 3266 98196 3278
rect 99820 3444 99876 3454
rect 99820 800 99876 3388
rect 99932 2772 99988 34636
rect 101164 34692 101220 34702
rect 101500 34692 101556 36428
rect 101612 36418 101668 36428
rect 101612 35812 101668 35822
rect 101612 35718 101668 35756
rect 101836 35698 101892 36652
rect 101836 35646 101838 35698
rect 101890 35646 101892 35698
rect 101836 35634 101892 35646
rect 101164 34690 101556 34692
rect 101164 34638 101166 34690
rect 101218 34638 101556 34690
rect 101164 34636 101556 34638
rect 101612 34692 101668 34702
rect 100716 33796 100772 33806
rect 100716 32788 100772 33740
rect 100716 32722 100772 32732
rect 101164 28084 101220 34636
rect 101612 34598 101668 34636
rect 102060 34690 102116 34702
rect 102060 34638 102062 34690
rect 102114 34638 102116 34690
rect 101164 28018 101220 28028
rect 101612 32788 101668 32798
rect 101612 8428 101668 32732
rect 102060 29540 102116 34638
rect 102172 34244 102228 36988
rect 102284 35812 102340 39200
rect 102396 36596 102452 36606
rect 102396 36502 102452 36540
rect 103180 36596 103236 39200
rect 103740 38052 103796 38062
rect 103180 36530 103236 36540
rect 103516 37156 103572 37166
rect 102284 35746 102340 35756
rect 102844 35812 102900 35822
rect 102844 35718 102900 35756
rect 103516 35698 103572 37100
rect 103740 36484 103796 37996
rect 103516 35646 103518 35698
rect 103570 35646 103572 35698
rect 103516 35634 103572 35646
rect 103628 36482 103796 36484
rect 103628 36430 103742 36482
rect 103794 36430 103796 36482
rect 103628 36428 103796 36430
rect 102172 34178 102228 34188
rect 102396 34802 102452 34814
rect 102396 34750 102398 34802
rect 102450 34750 102452 34802
rect 102396 34020 102452 34750
rect 102956 34802 103012 34814
rect 102956 34750 102958 34802
rect 103010 34750 103012 34802
rect 102956 34692 103012 34750
rect 103292 34804 103348 34814
rect 103292 34710 103348 34748
rect 102956 34626 103012 34636
rect 103516 34356 103572 34366
rect 103628 34356 103684 36428
rect 103740 36418 103796 36428
rect 103516 34354 103684 34356
rect 103516 34302 103518 34354
rect 103570 34302 103684 34354
rect 103516 34300 103684 34302
rect 103740 35812 103796 35822
rect 103516 34290 103572 34300
rect 102620 34020 102676 34030
rect 102396 34018 102676 34020
rect 102396 33966 102622 34018
rect 102674 33966 102676 34018
rect 102396 33964 102676 33966
rect 102508 33684 102564 33694
rect 102508 33348 102564 33628
rect 102508 33282 102564 33292
rect 102620 33124 102676 33964
rect 102620 33058 102676 33068
rect 103740 31108 103796 35756
rect 103852 35028 103908 35038
rect 104076 35028 104132 39200
rect 104188 37156 104244 37166
rect 104188 35922 104244 37100
rect 104412 36596 104468 36606
rect 104412 36502 104468 36540
rect 104188 35870 104190 35922
rect 104242 35870 104244 35922
rect 104188 35858 104244 35870
rect 104972 35028 105028 39200
rect 105644 36372 105700 36382
rect 105420 36370 105700 36372
rect 105420 36318 105646 36370
rect 105698 36318 105700 36370
rect 105420 36316 105700 36318
rect 105196 35700 105252 35710
rect 103852 35026 104580 35028
rect 103852 34974 103854 35026
rect 103906 34974 104580 35026
rect 103852 34972 104580 34974
rect 103852 34962 103908 34972
rect 104524 34914 104580 34972
rect 104972 34962 105028 34972
rect 105084 35698 105252 35700
rect 105084 35646 105198 35698
rect 105250 35646 105252 35698
rect 105084 35644 105252 35646
rect 104524 34862 104526 34914
rect 104578 34862 104580 34914
rect 104524 34850 104580 34862
rect 104300 34690 104356 34702
rect 104300 34638 104302 34690
rect 104354 34638 104356 34690
rect 104300 33796 104356 34638
rect 104300 33730 104356 33740
rect 104412 34020 104468 34030
rect 105084 34020 105140 35644
rect 105196 35634 105252 35644
rect 104412 34018 105140 34020
rect 104412 33966 104414 34018
rect 104466 33966 105140 34018
rect 104412 33964 105140 33966
rect 105196 34914 105252 34926
rect 105196 34862 105198 34914
rect 105250 34862 105252 34914
rect 105196 34018 105252 34862
rect 105196 33966 105198 34018
rect 105250 33966 105252 34018
rect 103740 31042 103796 31052
rect 102060 29474 102116 29484
rect 103292 24724 103348 24734
rect 103292 8932 103348 24668
rect 104412 17780 104468 33964
rect 105084 33122 105140 33134
rect 105084 33070 105086 33122
rect 105138 33070 105140 33122
rect 105084 32452 105140 33070
rect 105196 32676 105252 33966
rect 105196 32610 105252 32620
rect 105420 32452 105476 36316
rect 105644 36306 105700 36316
rect 105532 35810 105588 35822
rect 105532 35758 105534 35810
rect 105586 35758 105588 35810
rect 105532 35476 105588 35758
rect 105532 35410 105588 35420
rect 105868 35252 105924 39200
rect 106764 39060 106820 39200
rect 107100 39060 107156 39228
rect 106764 39004 107156 39060
rect 105644 35196 105924 35252
rect 106204 36484 106260 36494
rect 106204 36370 106260 36428
rect 106204 36318 106206 36370
rect 106258 36318 106260 36370
rect 106204 35698 106260 36318
rect 106428 36482 106484 36494
rect 106428 36430 106430 36482
rect 106482 36430 106484 36482
rect 106428 36372 106484 36430
rect 106428 36306 106484 36316
rect 107212 36372 107268 36382
rect 106764 36258 106820 36270
rect 106764 36206 106766 36258
rect 106818 36206 106820 36258
rect 106316 35812 106372 35822
rect 106316 35718 106372 35756
rect 106204 35646 106206 35698
rect 106258 35646 106260 35698
rect 105084 32396 105476 32452
rect 105532 34468 105588 34478
rect 105084 30884 105140 32396
rect 105084 30818 105140 30828
rect 105532 29988 105588 34412
rect 105644 34354 105700 35196
rect 105868 35028 105924 35038
rect 105868 34934 105924 34972
rect 105644 34302 105646 34354
rect 105698 34302 105700 34354
rect 105644 34244 105700 34302
rect 105644 34178 105700 34188
rect 106092 34242 106148 34254
rect 106092 34190 106094 34242
rect 106146 34190 106148 34242
rect 106092 33684 106148 34190
rect 106092 33618 106148 33628
rect 105756 33572 105812 33582
rect 105756 33458 105812 33516
rect 105756 33406 105758 33458
rect 105810 33406 105812 33458
rect 105756 33394 105812 33406
rect 106204 33572 106260 35646
rect 106540 35588 106596 35598
rect 106428 34244 106484 34254
rect 106428 34150 106484 34188
rect 106204 33458 106260 33516
rect 106204 33406 106206 33458
rect 106258 33406 106260 33458
rect 106204 33394 106260 33406
rect 105532 29922 105588 29932
rect 106540 20188 106596 35532
rect 106652 33570 106708 33582
rect 106652 33518 106654 33570
rect 106706 33518 106708 33570
rect 106652 33122 106708 33518
rect 106652 33070 106654 33122
rect 106706 33070 106708 33122
rect 106652 24612 106708 33070
rect 106652 24546 106708 24556
rect 106540 20132 106708 20188
rect 104412 17714 104468 17724
rect 104188 17668 104244 17678
rect 104188 11844 104244 17612
rect 104188 11778 104244 11788
rect 103292 8866 103348 8876
rect 105196 8930 105252 8942
rect 105196 8878 105198 8930
rect 105250 8878 105252 8930
rect 101500 8372 101668 8428
rect 105196 8428 105252 8878
rect 105196 8372 105588 8428
rect 101276 3780 101332 3790
rect 101276 3554 101332 3724
rect 101276 3502 101278 3554
rect 101330 3502 101332 3554
rect 101276 3490 101332 3502
rect 100380 3444 100436 3454
rect 100380 3350 100436 3388
rect 101164 3444 101220 3454
rect 99932 2706 99988 2716
rect 101164 800 101220 3388
rect 101500 2884 101556 8372
rect 104524 8260 104580 8270
rect 104524 8258 105364 8260
rect 104524 8206 104526 8258
rect 104578 8206 105364 8258
rect 104524 8204 105364 8206
rect 104524 8194 104580 8204
rect 102956 8036 103012 8046
rect 102508 6692 102564 6702
rect 102508 6466 102564 6636
rect 102508 6414 102510 6466
rect 102562 6414 102564 6466
rect 102508 5908 102564 6414
rect 102508 5842 102564 5852
rect 102956 6466 103012 7980
rect 103964 8036 104020 8046
rect 103964 7942 104020 7980
rect 104748 8034 104804 8046
rect 104748 7982 104750 8034
rect 104802 7982 104804 8034
rect 104076 7588 104132 7598
rect 104076 7494 104132 7532
rect 104412 7586 104468 7598
rect 104412 7534 104414 7586
rect 104466 7534 104468 7586
rect 102956 6414 102958 6466
rect 103010 6414 103012 6466
rect 102732 5794 102788 5806
rect 102732 5742 102734 5794
rect 102786 5742 102788 5794
rect 102732 5684 102788 5742
rect 102732 5618 102788 5628
rect 102620 5124 102676 5134
rect 102620 5030 102676 5068
rect 101612 4226 101668 4238
rect 101612 4174 101614 4226
rect 101666 4174 101668 4226
rect 101612 3444 101668 4174
rect 102732 3780 102788 3790
rect 102732 3666 102788 3724
rect 102732 3614 102734 3666
rect 102786 3614 102788 3666
rect 102732 3602 102788 3614
rect 102956 3556 103012 6414
rect 103068 7364 103124 7374
rect 103068 5346 103124 7308
rect 103516 7364 103572 7374
rect 103516 7270 103572 7308
rect 104412 6692 104468 7534
rect 104412 6626 104468 6636
rect 104748 6580 104804 7982
rect 105308 7364 105364 8204
rect 105532 8148 105588 8372
rect 105756 8260 105812 8270
rect 105756 8166 105812 8204
rect 106652 8260 106708 20132
rect 106652 8194 106708 8204
rect 105532 8082 105588 8092
rect 105980 8148 106036 8158
rect 105420 8034 105476 8046
rect 105420 7982 105422 8034
rect 105474 7982 105476 8034
rect 105420 7588 105476 7982
rect 105420 7522 105476 7532
rect 105980 7700 106036 8092
rect 106316 8146 106372 8158
rect 106316 8094 106318 8146
rect 106370 8094 106372 8146
rect 106316 8036 106372 8094
rect 106316 7970 106372 7980
rect 105980 7586 106036 7644
rect 105980 7534 105982 7586
rect 106034 7534 106036 7586
rect 105980 7522 106036 7534
rect 106316 7586 106372 7598
rect 106316 7534 106318 7586
rect 106370 7534 106372 7586
rect 105756 7476 105812 7486
rect 105756 7382 105812 7420
rect 105420 7364 105476 7374
rect 105308 7362 105476 7364
rect 105308 7310 105422 7362
rect 105474 7310 105476 7362
rect 105308 7308 105476 7310
rect 105420 7298 105476 7308
rect 106316 7364 106372 7534
rect 106764 7476 106820 36206
rect 106988 35474 107044 35486
rect 106988 35422 106990 35474
rect 107042 35422 107044 35474
rect 106988 35140 107044 35422
rect 106988 35074 107044 35084
rect 106988 34914 107044 34926
rect 106988 34862 106990 34914
rect 107042 34862 107044 34914
rect 106988 34804 107044 34862
rect 106988 34738 107044 34748
rect 106988 34130 107044 34142
rect 106988 34078 106990 34130
rect 107042 34078 107044 34130
rect 106988 33570 107044 34078
rect 106988 33518 106990 33570
rect 107042 33518 107044 33570
rect 106988 33506 107044 33518
rect 107212 33458 107268 36316
rect 107324 35588 107380 35598
rect 107324 35494 107380 35532
rect 107324 35252 107380 35262
rect 107436 35252 107492 39228
rect 107632 39200 107744 40000
rect 108528 39200 108640 40000
rect 109424 39200 109536 40000
rect 110320 39200 110432 40000
rect 111216 39200 111328 40000
rect 112112 39200 112224 40000
rect 113008 39200 113120 40000
rect 113904 39200 114016 40000
rect 114800 39200 114912 40000
rect 115696 39200 115808 40000
rect 116592 39200 116704 40000
rect 117488 39200 117600 40000
rect 118384 39200 118496 40000
rect 119280 39200 119392 40000
rect 119644 39228 120036 39284
rect 107548 36258 107604 36270
rect 107548 36206 107550 36258
rect 107602 36206 107604 36258
rect 107548 35812 107604 36206
rect 107548 35746 107604 35756
rect 107660 35476 107716 39200
rect 108556 37268 108612 39200
rect 108556 37212 109060 37268
rect 108668 36484 108724 36494
rect 108556 36370 108612 36382
rect 108556 36318 108558 36370
rect 108610 36318 108612 36370
rect 108332 35810 108388 35822
rect 108332 35758 108334 35810
rect 108386 35758 108388 35810
rect 107996 35700 108052 35710
rect 107996 35698 108276 35700
rect 107996 35646 107998 35698
rect 108050 35646 108276 35698
rect 107996 35644 108276 35646
rect 107996 35634 108052 35644
rect 107660 35420 108164 35476
rect 107436 35196 107716 35252
rect 107324 34354 107380 35196
rect 107660 35026 107716 35196
rect 107660 34974 107662 35026
rect 107714 34974 107716 35026
rect 107660 34962 107716 34974
rect 107324 34302 107326 34354
rect 107378 34302 107380 34354
rect 107324 34290 107380 34302
rect 107884 34244 107940 34254
rect 107212 33406 107214 33458
rect 107266 33406 107268 33458
rect 107212 33394 107268 33406
rect 107548 34242 107940 34244
rect 107548 34190 107886 34242
rect 107938 34190 107940 34242
rect 107548 34188 107940 34190
rect 106764 7410 106820 7420
rect 106876 33124 106932 33134
rect 106316 7298 106372 7308
rect 105980 6692 106036 6702
rect 105980 6598 106036 6636
rect 106652 6690 106708 6702
rect 106652 6638 106654 6690
rect 106706 6638 106708 6690
rect 104748 6514 104804 6524
rect 106092 6580 106148 6590
rect 103740 6466 103796 6478
rect 103740 6414 103742 6466
rect 103794 6414 103796 6466
rect 103740 6132 103796 6414
rect 105756 6468 105812 6478
rect 103740 6066 103796 6076
rect 104412 6132 104468 6142
rect 104412 6038 104468 6076
rect 104524 5908 104580 5918
rect 103180 5794 103236 5806
rect 103180 5742 103182 5794
rect 103234 5742 103236 5794
rect 103180 5684 103236 5742
rect 103180 5618 103236 5628
rect 103628 5794 103684 5806
rect 103628 5742 103630 5794
rect 103682 5742 103684 5794
rect 103628 5684 103684 5742
rect 104300 5794 104356 5806
rect 104300 5742 104302 5794
rect 104354 5742 104356 5794
rect 103628 5618 103684 5628
rect 103740 5682 103796 5694
rect 103740 5630 103742 5682
rect 103794 5630 103796 5682
rect 103068 5294 103070 5346
rect 103122 5294 103124 5346
rect 103068 3668 103124 5294
rect 103740 4898 103796 5630
rect 104300 5684 104356 5742
rect 104300 5618 104356 5628
rect 103740 4846 103742 4898
rect 103794 4846 103796 4898
rect 103740 4834 103796 4846
rect 103964 5124 104020 5134
rect 103964 4562 104020 5068
rect 103964 4510 103966 4562
rect 104018 4510 104020 4562
rect 103964 4498 104020 4510
rect 104412 4564 104468 4574
rect 104524 4564 104580 5852
rect 105308 5908 105364 5918
rect 105308 5814 105364 5852
rect 105756 5906 105812 6412
rect 105756 5854 105758 5906
rect 105810 5854 105812 5906
rect 105756 5842 105812 5854
rect 104412 4562 104580 4564
rect 104412 4510 104414 4562
rect 104466 4510 104580 4562
rect 104412 4508 104580 4510
rect 105308 5124 105364 5134
rect 104412 4498 104468 4508
rect 105308 4338 105364 5068
rect 106092 5122 106148 6524
rect 106652 5908 106708 6638
rect 106652 5842 106708 5852
rect 106092 5070 106094 5122
rect 106146 5070 106148 5122
rect 106092 5058 106148 5070
rect 106764 5124 106820 5134
rect 106764 5030 106820 5068
rect 105308 4286 105310 4338
rect 105362 4286 105364 4338
rect 105308 4274 105364 4286
rect 105756 4340 105812 4350
rect 105756 4246 105812 4284
rect 103068 3602 103124 3612
rect 102956 3490 103012 3500
rect 105308 3556 105364 3566
rect 105308 3462 105364 3500
rect 101612 3378 101668 3388
rect 101836 3444 101892 3454
rect 101836 3350 101892 3388
rect 103852 3444 103908 3454
rect 102172 3332 102228 3342
rect 102172 3238 102228 3276
rect 101500 2818 101556 2828
rect 103852 800 103908 3388
rect 104412 3444 104468 3454
rect 104412 3350 104468 3388
rect 105196 3444 105252 3454
rect 105196 800 105252 3388
rect 106204 3444 106260 3454
rect 106204 3350 106260 3388
rect 106652 3444 106708 3454
rect 106652 3350 106708 3388
rect 105868 3330 105924 3342
rect 105868 3278 105870 3330
rect 105922 3278 105924 3330
rect 105868 2994 105924 3278
rect 105868 2942 105870 2994
rect 105922 2942 105924 2994
rect 105868 2930 105924 2942
rect 106876 2994 106932 33068
rect 107548 32564 107604 34188
rect 107884 34178 107940 34188
rect 108108 34132 108164 35420
rect 107996 34130 108164 34132
rect 107996 34078 108110 34130
rect 108162 34078 108164 34130
rect 107996 34076 108164 34078
rect 107660 33460 107716 33470
rect 107996 33460 108052 34076
rect 108108 34066 108164 34076
rect 107660 33458 108052 33460
rect 107660 33406 107662 33458
rect 107714 33406 108052 33458
rect 107660 33404 108052 33406
rect 107660 33394 107716 33404
rect 107996 33124 108052 33134
rect 108220 33124 108276 35644
rect 108332 35364 108388 35758
rect 108332 35298 108388 35308
rect 108556 34692 108612 36318
rect 108668 36148 108724 36428
rect 108668 36082 108724 36092
rect 108556 34626 108612 34636
rect 108780 35140 108836 35150
rect 108780 34354 108836 35084
rect 109004 35140 109060 37212
rect 109340 36484 109396 36494
rect 109340 36390 109396 36428
rect 109228 36148 109284 36158
rect 109228 35698 109284 36092
rect 109228 35646 109230 35698
rect 109282 35646 109284 35698
rect 109228 35634 109284 35646
rect 109340 35810 109396 35822
rect 109340 35758 109342 35810
rect 109394 35758 109396 35810
rect 109004 35074 109060 35084
rect 109228 35476 109284 35486
rect 109228 34914 109284 35420
rect 109228 34862 109230 34914
rect 109282 34862 109284 34914
rect 109228 34850 109284 34862
rect 108780 34302 108782 34354
rect 108834 34302 108836 34354
rect 108780 33908 108836 34302
rect 109228 34468 109284 34478
rect 109228 34354 109284 34412
rect 109228 34302 109230 34354
rect 109282 34302 109284 34354
rect 109228 34290 109284 34302
rect 108780 33842 108836 33852
rect 109340 33684 109396 35758
rect 109452 34468 109508 39200
rect 110236 37940 110292 37950
rect 110124 36484 110180 36494
rect 109676 36260 109732 36270
rect 109452 34402 109508 34412
rect 109564 36258 109732 36260
rect 109564 36206 109678 36258
rect 109730 36206 109732 36258
rect 109564 36204 109732 36206
rect 109228 33628 109396 33684
rect 108052 33068 108276 33124
rect 108332 33572 108388 33582
rect 107996 33030 108052 33068
rect 108220 32788 108276 32798
rect 108332 32788 108388 33516
rect 109228 33460 109284 33628
rect 108220 32786 108388 32788
rect 108220 32734 108222 32786
rect 108274 32734 108388 32786
rect 108220 32732 108388 32734
rect 109116 33404 109284 33460
rect 109452 33572 109508 33582
rect 109452 33458 109508 33516
rect 109452 33406 109454 33458
rect 109506 33406 109508 33458
rect 109116 33122 109172 33404
rect 109452 33394 109508 33406
rect 109116 33070 109118 33122
rect 109170 33070 109172 33122
rect 108220 32722 108276 32732
rect 107548 32498 107604 32508
rect 109116 31556 109172 33070
rect 109116 31490 109172 31500
rect 107100 8260 107156 8270
rect 107100 8166 107156 8204
rect 107100 7700 107156 7710
rect 107100 7606 107156 7644
rect 107548 7476 107604 7486
rect 107548 7382 107604 7420
rect 107436 6578 107492 6590
rect 107436 6526 107438 6578
rect 107490 6526 107492 6578
rect 107100 6468 107156 6478
rect 107100 6374 107156 6412
rect 107212 4898 107268 4910
rect 107212 4846 107214 4898
rect 107266 4846 107268 4898
rect 107212 4340 107268 4846
rect 107212 4274 107268 4284
rect 107436 3780 107492 6526
rect 109116 6468 109172 6478
rect 109116 6466 109396 6468
rect 109116 6414 109118 6466
rect 109170 6414 109396 6466
rect 109116 6412 109396 6414
rect 109116 6402 109172 6412
rect 108220 6132 108276 6142
rect 108220 6038 108276 6076
rect 109228 6132 109284 6142
rect 109228 6038 109284 6076
rect 108332 6020 108388 6030
rect 107548 5236 107604 5246
rect 107548 5010 107604 5180
rect 108220 5236 108276 5246
rect 108332 5236 108388 5964
rect 109340 6020 109396 6412
rect 109340 5926 109396 5964
rect 108780 5684 108836 5694
rect 108780 5682 108948 5684
rect 108780 5630 108782 5682
rect 108834 5630 108948 5682
rect 108780 5628 108948 5630
rect 108780 5618 108836 5628
rect 108220 5234 108388 5236
rect 108220 5182 108222 5234
rect 108274 5182 108388 5234
rect 108220 5180 108388 5182
rect 108220 5170 108276 5180
rect 107548 4958 107550 5010
rect 107602 4958 107604 5010
rect 107548 4946 107604 4958
rect 108108 4898 108164 4910
rect 108108 4846 108110 4898
rect 108162 4846 108164 4898
rect 108108 4562 108164 4846
rect 108108 4510 108110 4562
rect 108162 4510 108164 4562
rect 108108 4498 108164 4510
rect 108444 4564 108500 4574
rect 107436 3714 107492 3724
rect 107884 4228 107940 4238
rect 106876 2942 106878 2994
rect 106930 2942 106932 2994
rect 106876 2930 106932 2942
rect 107884 800 107940 4172
rect 108108 3780 108164 3790
rect 108108 3686 108164 3724
rect 108444 3778 108500 4508
rect 108780 4114 108836 4126
rect 108780 4062 108782 4114
rect 108834 4062 108836 4114
rect 108780 3892 108836 4062
rect 108780 3826 108836 3836
rect 108444 3726 108446 3778
rect 108498 3726 108500 3778
rect 108444 3714 108500 3726
rect 108892 3556 108948 5628
rect 109564 5346 109620 36204
rect 109676 36194 109732 36204
rect 110012 35474 110068 35486
rect 110012 35422 110014 35474
rect 110066 35422 110068 35474
rect 109788 35140 109844 35150
rect 109788 35026 109844 35084
rect 109788 34974 109790 35026
rect 109842 34974 109844 35026
rect 109788 34962 109844 34974
rect 109900 34468 109956 34478
rect 109676 34242 109732 34254
rect 109676 34190 109678 34242
rect 109730 34190 109732 34242
rect 109676 25508 109732 34190
rect 109900 34130 109956 34412
rect 109900 34078 109902 34130
rect 109954 34078 109956 34130
rect 109900 34066 109956 34078
rect 110012 33460 110068 35422
rect 110012 33394 110068 33404
rect 110124 33458 110180 36428
rect 110236 36372 110292 37884
rect 110348 36708 110404 39200
rect 110348 36642 110404 36652
rect 111132 38836 111188 38846
rect 110348 36372 110404 36382
rect 110236 36370 110404 36372
rect 110236 36318 110350 36370
rect 110402 36318 110404 36370
rect 110236 36316 110404 36318
rect 110348 36306 110404 36316
rect 110684 36370 110740 36382
rect 110684 36318 110686 36370
rect 110738 36318 110740 36370
rect 110348 35476 110404 35486
rect 110348 35382 110404 35420
rect 110124 33406 110126 33458
rect 110178 33406 110180 33458
rect 110124 33348 110180 33406
rect 110124 33282 110180 33292
rect 110684 33236 110740 36318
rect 111020 35698 111076 35710
rect 111020 35646 111022 35698
rect 111074 35646 111076 35698
rect 110796 34692 110852 34702
rect 110796 34598 110852 34636
rect 110796 34018 110852 34030
rect 110796 33966 110798 34018
rect 110850 33966 110852 34018
rect 110796 33460 110852 33966
rect 110796 33394 110852 33404
rect 111020 33572 111076 35646
rect 111132 34804 111188 38780
rect 111244 35028 111300 39200
rect 112140 36596 112196 39200
rect 112140 36530 112196 36540
rect 112252 36708 112308 36718
rect 112252 36594 112308 36652
rect 112252 36542 112254 36594
rect 112306 36542 112308 36594
rect 112252 36530 112308 36542
rect 111580 36484 111636 36494
rect 111468 36482 111636 36484
rect 111468 36430 111582 36482
rect 111634 36430 111636 36482
rect 111468 36428 111636 36430
rect 111356 35924 111412 35934
rect 111356 35830 111412 35868
rect 111468 35252 111524 36428
rect 111580 36418 111636 36428
rect 111672 36092 111936 36102
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111672 36026 111936 36036
rect 112252 35812 112308 35822
rect 112252 35718 112308 35756
rect 111468 35186 111524 35196
rect 112028 35698 112084 35710
rect 112028 35646 112030 35698
rect 112082 35646 112084 35698
rect 111244 34972 111748 35028
rect 111468 34804 111524 34814
rect 111132 34802 111524 34804
rect 111132 34750 111470 34802
rect 111522 34750 111524 34802
rect 111132 34748 111524 34750
rect 111468 34738 111524 34748
rect 111580 34692 111636 34972
rect 111692 34914 111748 34972
rect 111692 34862 111694 34914
rect 111746 34862 111748 34914
rect 111692 34850 111748 34862
rect 111580 34626 111636 34636
rect 111244 34580 111300 34590
rect 111244 34354 111300 34524
rect 111672 34524 111936 34534
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111672 34458 111936 34468
rect 111244 34302 111246 34354
rect 111298 34302 111300 34354
rect 111244 34290 111300 34302
rect 111580 34020 111636 34030
rect 112028 34020 112084 35646
rect 112812 35476 112868 35486
rect 110908 33236 110964 33246
rect 110684 33234 110964 33236
rect 110684 33182 110910 33234
rect 110962 33182 110964 33234
rect 110684 33180 110964 33182
rect 110684 31948 110740 33180
rect 110908 33124 110964 33180
rect 110908 33058 110964 33068
rect 111020 32788 111076 33516
rect 111020 32722 111076 32732
rect 111468 34018 112084 34020
rect 111468 33966 111582 34018
rect 111634 33966 112084 34018
rect 111468 33964 112084 33966
rect 112252 34690 112308 34702
rect 112252 34638 112254 34690
rect 112306 34638 112308 34690
rect 109676 25442 109732 25452
rect 110348 31892 110740 31948
rect 110236 6020 110292 6030
rect 110236 5926 110292 5964
rect 109564 5294 109566 5346
rect 109618 5294 109620 5346
rect 109228 5236 109284 5246
rect 109228 5142 109284 5180
rect 109564 5236 109620 5294
rect 109564 5170 109620 5180
rect 109900 5794 109956 5806
rect 109900 5742 109902 5794
rect 109954 5742 109956 5794
rect 109900 5012 109956 5742
rect 110236 5684 110292 5694
rect 110236 5122 110292 5628
rect 110236 5070 110238 5122
rect 110290 5070 110292 5122
rect 110236 5058 110292 5070
rect 110124 5012 110180 5022
rect 109900 5010 110180 5012
rect 109900 4958 110126 5010
rect 110178 4958 110180 5010
rect 109900 4956 110180 4958
rect 109452 4228 109508 4238
rect 109452 4134 109508 4172
rect 110124 3892 110180 4956
rect 110124 3826 110180 3836
rect 109004 3556 109060 3566
rect 108892 3500 109004 3556
rect 109004 3442 109060 3500
rect 109228 3556 109284 3566
rect 109228 3462 109284 3500
rect 109004 3390 109006 3442
rect 109058 3390 109060 3442
rect 109004 3378 109060 3390
rect 109900 3444 109956 3454
rect 109228 924 109508 980
rect 109228 800 109284 924
rect 69132 700 69524 756
rect 70224 0 70336 800
rect 71568 0 71680 800
rect 72912 0 73024 800
rect 74256 0 74368 800
rect 75600 0 75712 800
rect 76944 0 77056 800
rect 78288 0 78400 800
rect 79632 0 79744 800
rect 80976 0 81088 800
rect 82320 0 82432 800
rect 83664 0 83776 800
rect 85008 0 85120 800
rect 86352 0 86464 800
rect 87696 0 87808 800
rect 89040 0 89152 800
rect 90384 0 90496 800
rect 91728 0 91840 800
rect 93072 0 93184 800
rect 94416 0 94528 800
rect 95760 0 95872 800
rect 97104 0 97216 800
rect 98448 0 98560 800
rect 99792 0 99904 800
rect 101136 0 101248 800
rect 102480 0 102592 800
rect 103824 0 103936 800
rect 105168 0 105280 800
rect 106512 0 106624 800
rect 107856 0 107968 800
rect 109200 0 109312 800
rect 109452 756 109508 924
rect 109900 756 109956 3388
rect 110236 3332 110292 3342
rect 110348 3332 110404 31892
rect 111468 26068 111524 33964
rect 111580 33954 111636 33964
rect 112252 33572 112308 34638
rect 112252 33506 112308 33516
rect 111672 32956 111936 32966
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111672 32890 111936 32900
rect 111672 31388 111936 31398
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111672 31322 111936 31332
rect 111672 29820 111936 29830
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111672 29754 111936 29764
rect 111672 28252 111936 28262
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111672 28186 111936 28196
rect 111672 26684 111936 26694
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111672 26618 111936 26628
rect 111468 26002 111524 26012
rect 111672 25116 111936 25126
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111672 25050 111936 25060
rect 111672 23548 111936 23558
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111672 23482 111936 23492
rect 111672 21980 111936 21990
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111672 21914 111936 21924
rect 111672 20412 111936 20422
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111672 20346 111936 20356
rect 111672 18844 111936 18854
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111672 18778 111936 18788
rect 111672 17276 111936 17286
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111672 17210 111936 17220
rect 111672 15708 111936 15718
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111672 15642 111936 15652
rect 111672 14140 111936 14150
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111672 14074 111936 14084
rect 111672 12572 111936 12582
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111672 12506 111936 12516
rect 111672 11004 111936 11014
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111672 10938 111936 10948
rect 111672 9436 111936 9446
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111672 9370 111936 9380
rect 111672 7868 111936 7878
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111672 7802 111936 7812
rect 110796 6466 110852 6478
rect 110796 6414 110798 6466
rect 110850 6414 110852 6466
rect 110796 6132 110852 6414
rect 111672 6300 111936 6310
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111672 6234 111936 6244
rect 110796 5908 110852 6076
rect 111020 5908 111076 5918
rect 110796 5906 111076 5908
rect 110796 5854 111022 5906
rect 111074 5854 111076 5906
rect 110796 5852 111076 5854
rect 110908 5684 110964 5694
rect 110908 5236 110964 5628
rect 111020 5348 111076 5852
rect 112364 5908 112420 5918
rect 112364 5814 112420 5852
rect 111580 5796 111636 5806
rect 111580 5702 111636 5740
rect 111020 5282 111076 5292
rect 110684 5234 110964 5236
rect 110684 5182 110910 5234
rect 110962 5182 110964 5234
rect 110684 5180 110964 5182
rect 110460 4452 110516 4462
rect 110460 4338 110516 4396
rect 110460 4286 110462 4338
rect 110514 4286 110516 4338
rect 110460 4274 110516 4286
rect 110684 3666 110740 5180
rect 110908 5170 110964 5180
rect 111356 5236 111412 5246
rect 111356 5142 111412 5180
rect 111672 4732 111936 4742
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111672 4666 111936 4676
rect 110908 4564 110964 4574
rect 110908 4470 110964 4508
rect 112812 4564 112868 35420
rect 113036 35140 113092 39200
rect 113148 37716 113204 37726
rect 113148 35922 113204 37660
rect 113148 35870 113150 35922
rect 113202 35870 113204 35922
rect 113148 35858 113204 35870
rect 113372 36482 113428 36494
rect 113372 36430 113374 36482
rect 113426 36430 113428 36482
rect 113372 35924 113428 36430
rect 113372 35858 113428 35868
rect 113484 35700 113540 35710
rect 113484 35606 113540 35644
rect 113932 35588 113988 39200
rect 114044 36596 114100 36606
rect 114044 36502 114100 36540
rect 114828 36148 114884 39200
rect 115724 36596 115780 39200
rect 116620 36820 116676 39200
rect 116620 36764 117124 36820
rect 115724 36530 115780 36540
rect 116620 36596 116676 36606
rect 116620 36502 116676 36540
rect 115948 36482 116004 36494
rect 115948 36430 115950 36482
rect 116002 36430 116004 36482
rect 115500 36258 115556 36270
rect 115500 36206 115502 36258
rect 115554 36206 115556 36258
rect 114828 36092 115332 36148
rect 114268 35812 114324 35822
rect 114268 35698 114324 35756
rect 114268 35646 114270 35698
rect 114322 35646 114324 35698
rect 114268 35634 114324 35646
rect 113932 35522 113988 35532
rect 114828 35588 114884 35598
rect 114828 35494 114884 35532
rect 115052 35476 115108 35486
rect 113036 35074 113092 35084
rect 114380 35140 114436 35150
rect 113148 34802 113204 34814
rect 113148 34750 113150 34802
rect 113202 34750 113204 34802
rect 113036 34020 113092 34030
rect 113148 34020 113204 34750
rect 114380 34804 114436 35084
rect 114380 34710 114436 34748
rect 113484 34692 113540 34702
rect 113484 34598 113540 34636
rect 114044 34690 114100 34702
rect 114044 34638 114046 34690
rect 114098 34638 114100 34690
rect 113036 34018 113204 34020
rect 113036 33966 113038 34018
rect 113090 33966 113204 34018
rect 113036 33964 113204 33966
rect 113036 33954 113092 33964
rect 113148 12740 113204 33964
rect 113596 34242 113652 34254
rect 113596 34190 113598 34242
rect 113650 34190 113652 34242
rect 113596 27972 113652 34190
rect 114044 34244 114100 34638
rect 115052 34690 115108 35420
rect 115276 34916 115332 36092
rect 115500 35700 115556 36206
rect 115500 35140 115556 35644
rect 115500 35074 115556 35084
rect 115052 34638 115054 34690
rect 115106 34638 115108 34690
rect 115052 34626 115108 34638
rect 115164 34914 115332 34916
rect 115164 34862 115278 34914
rect 115330 34862 115332 34914
rect 115164 34860 115332 34862
rect 115164 34468 115220 34860
rect 115276 34850 115332 34860
rect 115836 34804 115892 34814
rect 115836 34710 115892 34748
rect 115948 34692 116004 36430
rect 116844 36260 116900 36270
rect 116844 35922 116900 36204
rect 116844 35870 116846 35922
rect 116898 35870 116900 35922
rect 116844 35858 116900 35870
rect 116284 35812 116340 35822
rect 116284 35718 116340 35756
rect 116060 35698 116116 35710
rect 116060 35646 116062 35698
rect 116114 35646 116116 35698
rect 116060 34692 116116 35646
rect 117068 35698 117124 36764
rect 117068 35646 117070 35698
rect 117122 35646 117124 35698
rect 117068 35026 117124 35646
rect 117516 35588 117572 39200
rect 117852 36482 117908 36494
rect 117852 36430 117854 36482
rect 117906 36430 117908 36482
rect 117516 35522 117572 35532
rect 117628 36260 117684 36270
rect 117068 34974 117070 35026
rect 117122 34974 117124 35026
rect 117068 34962 117124 34974
rect 117516 35140 117572 35150
rect 116284 34692 116340 34702
rect 116060 34690 116340 34692
rect 116060 34638 116286 34690
rect 116338 34638 116340 34690
rect 116060 34636 116340 34638
rect 115948 34626 116004 34636
rect 114940 34412 115220 34468
rect 114940 34354 114996 34412
rect 114940 34302 114942 34354
rect 114994 34302 114996 34354
rect 114940 34290 114996 34302
rect 114044 34178 114100 34188
rect 113932 34130 113988 34142
rect 113932 34078 113934 34130
rect 113986 34078 113988 34130
rect 113932 33796 113988 34078
rect 113932 33730 113988 33740
rect 114380 34018 114436 34030
rect 114380 33966 114382 34018
rect 114434 33966 114436 34018
rect 114380 33796 114436 33966
rect 114380 33730 114436 33740
rect 113596 27906 113652 27916
rect 116284 26180 116340 34636
rect 116284 26114 116340 26124
rect 117516 34354 117572 35084
rect 117516 34302 117518 34354
rect 117570 34302 117572 34354
rect 113148 12674 113204 12684
rect 113372 12628 113428 12638
rect 113260 5908 113316 5918
rect 113260 5814 113316 5852
rect 112812 4498 112868 4508
rect 111356 4452 111412 4462
rect 111356 4358 111412 4396
rect 113372 4340 113428 12572
rect 115388 7588 115444 7598
rect 115388 7362 115444 7532
rect 116620 7588 116676 7598
rect 116620 7494 116676 7532
rect 116956 7586 117012 7598
rect 116956 7534 116958 7586
rect 117010 7534 117012 7586
rect 116396 7476 116452 7486
rect 116396 7382 116452 7420
rect 115388 7310 115390 7362
rect 115442 7310 115444 7362
rect 115052 7252 115108 7262
rect 114268 6804 114324 6814
rect 113708 6468 113764 6478
rect 113708 5906 113764 6412
rect 113708 5854 113710 5906
rect 113762 5854 113764 5906
rect 113708 5842 113764 5854
rect 113260 4284 113428 4340
rect 112364 3668 112420 3678
rect 110684 3614 110686 3666
rect 110738 3614 110740 3666
rect 110684 3556 110740 3614
rect 110684 3490 110740 3500
rect 112028 3666 112420 3668
rect 112028 3614 112366 3666
rect 112418 3614 112420 3666
rect 112028 3612 112420 3614
rect 111468 3444 111524 3454
rect 111468 3350 111524 3388
rect 110236 3330 110404 3332
rect 110236 3278 110238 3330
rect 110290 3278 110404 3330
rect 110236 3276 110404 3278
rect 110236 3266 110292 3276
rect 111672 3164 111936 3174
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111672 3098 111936 3108
rect 112028 980 112084 3612
rect 112364 3602 112420 3612
rect 113260 2548 113316 4284
rect 113708 4226 113764 4238
rect 113708 4174 113710 4226
rect 113762 4174 113764 4226
rect 113372 4116 113428 4126
rect 113372 3554 113428 4060
rect 113372 3502 113374 3554
rect 113426 3502 113428 3554
rect 113372 3490 113428 3502
rect 113708 3444 113764 4174
rect 113932 3444 113988 3454
rect 113708 3442 113988 3444
rect 113708 3390 113934 3442
rect 113986 3390 113988 3442
rect 113708 3388 113988 3390
rect 113260 2482 113316 2492
rect 111916 924 112084 980
rect 113260 924 113652 980
rect 111916 800 111972 924
rect 113260 800 113316 924
rect 109452 700 109956 756
rect 110544 0 110656 800
rect 111888 0 112000 800
rect 113232 0 113344 800
rect 113596 756 113652 924
rect 113932 756 113988 3388
rect 114268 3330 114324 6748
rect 115052 6690 115108 7196
rect 115052 6638 115054 6690
rect 115106 6638 115108 6690
rect 115052 6626 115108 6638
rect 114716 6468 114772 6478
rect 114716 6374 114772 6412
rect 114940 6020 114996 6030
rect 114940 5236 114996 5964
rect 115388 5796 115444 7310
rect 116956 7364 117012 7534
rect 116060 7252 116116 7262
rect 116060 7158 116116 7196
rect 115948 6020 116004 6030
rect 115388 5730 115444 5740
rect 115612 6018 116004 6020
rect 115612 5966 115950 6018
rect 116002 5966 116004 6018
rect 115612 5964 116004 5966
rect 115612 5346 115668 5964
rect 115948 5954 116004 5964
rect 115612 5294 115614 5346
rect 115666 5294 115668 5346
rect 115612 5282 115668 5294
rect 116732 5684 116788 5694
rect 116956 5684 117012 7308
rect 117516 6804 117572 34302
rect 117628 20188 117684 36204
rect 117852 36148 117908 36430
rect 118076 36484 118132 36494
rect 118412 36484 118468 39200
rect 119308 39060 119364 39200
rect 119644 39060 119700 39228
rect 119308 39004 119700 39060
rect 118748 37828 118804 37838
rect 119980 37828 120036 39228
rect 120176 39200 120288 40000
rect 120540 39228 120932 39284
rect 120204 39060 120260 39200
rect 120540 39060 120596 39228
rect 120204 39004 120596 39060
rect 119980 37772 120260 37828
rect 118412 36428 118692 36484
rect 118076 36370 118132 36428
rect 118076 36318 118078 36370
rect 118130 36318 118132 36370
rect 118076 36306 118132 36318
rect 118524 36258 118580 36270
rect 118524 36206 118526 36258
rect 118578 36206 118580 36258
rect 118524 36148 118580 36206
rect 117852 36092 118580 36148
rect 117740 35812 117796 35822
rect 117740 35698 117796 35756
rect 117740 35646 117742 35698
rect 117794 35646 117796 35698
rect 117740 35634 117796 35646
rect 118412 35588 118468 35598
rect 118412 35494 118468 35532
rect 117852 35140 117908 35150
rect 117852 34914 117908 35084
rect 117852 34862 117854 34914
rect 117906 34862 117908 34914
rect 117852 34850 117908 34862
rect 118188 34690 118244 34702
rect 118188 34638 118190 34690
rect 118242 34638 118244 34690
rect 118076 34468 118132 34478
rect 118076 33796 118132 34412
rect 117628 20132 117796 20188
rect 117740 7476 117796 20132
rect 118076 8428 118132 33740
rect 118188 33012 118244 34638
rect 118188 32946 118244 32956
rect 118524 12628 118580 36092
rect 118636 35140 118692 36428
rect 118636 35074 118692 35084
rect 118748 34802 118804 37772
rect 120204 36594 120260 37772
rect 120204 36542 120206 36594
rect 120258 36542 120260 36594
rect 120204 36530 120260 36542
rect 119532 36484 119588 36494
rect 119532 36390 119588 36428
rect 119868 35924 119924 35934
rect 119868 35830 119924 35868
rect 119644 35698 119700 35710
rect 119644 35646 119646 35698
rect 119698 35646 119700 35698
rect 119644 35588 119700 35646
rect 120316 35588 120372 35598
rect 119644 35586 120372 35588
rect 119644 35534 120318 35586
rect 120370 35534 120372 35586
rect 119644 35532 120372 35534
rect 120876 35588 120932 39228
rect 121072 39200 121184 40000
rect 121436 39228 121828 39284
rect 121100 39060 121156 39200
rect 121436 39060 121492 39228
rect 121100 39004 121492 39060
rect 121772 37828 121828 39228
rect 121968 39200 122080 40000
rect 122864 39200 122976 40000
rect 123760 39200 123872 40000
rect 124656 39200 124768 40000
rect 125552 39200 125664 40000
rect 126448 39200 126560 40000
rect 127344 39200 127456 40000
rect 128240 39200 128352 40000
rect 129136 39200 129248 40000
rect 130032 39200 130144 40000
rect 130928 39200 131040 40000
rect 131824 39200 131936 40000
rect 132720 39200 132832 40000
rect 133616 39200 133728 40000
rect 134512 39200 134624 40000
rect 135408 39200 135520 40000
rect 136304 39200 136416 40000
rect 137200 39200 137312 40000
rect 138096 39200 138208 40000
rect 138992 39200 139104 40000
rect 139888 39200 140000 40000
rect 140784 39200 140896 40000
rect 141680 39200 141792 40000
rect 142576 39200 142688 40000
rect 143472 39200 143584 40000
rect 144368 39200 144480 40000
rect 145264 39200 145376 40000
rect 121996 37940 122052 39200
rect 121996 37884 122164 37940
rect 121772 37772 122052 37828
rect 121548 37492 121604 37502
rect 121100 36820 121156 36830
rect 121100 35922 121156 36764
rect 121100 35870 121102 35922
rect 121154 35870 121156 35922
rect 121100 35858 121156 35870
rect 121324 36482 121380 36494
rect 121324 36430 121326 36482
rect 121378 36430 121380 36482
rect 121324 35924 121380 36430
rect 121324 35858 121380 35868
rect 121324 35698 121380 35710
rect 121324 35646 121326 35698
rect 121378 35646 121380 35698
rect 121324 35588 121380 35646
rect 120876 35532 121380 35588
rect 119532 35476 119588 35486
rect 118748 34750 118750 34802
rect 118802 34750 118804 34802
rect 118748 34738 118804 34750
rect 119084 34802 119140 34814
rect 119084 34750 119086 34802
rect 119138 34750 119140 34802
rect 119084 34020 119140 34750
rect 119308 34020 119364 34030
rect 119084 34018 119364 34020
rect 119084 33966 119310 34018
rect 119362 33966 119364 34018
rect 119084 33964 119364 33966
rect 119308 33796 119364 33964
rect 119308 33730 119364 33740
rect 118524 12562 118580 12572
rect 117740 7382 117796 7420
rect 117852 8372 118132 8428
rect 117516 6738 117572 6748
rect 117292 6466 117348 6478
rect 117292 6414 117294 6466
rect 117346 6414 117348 6466
rect 116732 5682 117012 5684
rect 116732 5630 116734 5682
rect 116786 5630 117012 5682
rect 116732 5628 117012 5630
rect 117180 6356 117236 6366
rect 114380 5124 114436 5134
rect 114940 5104 114996 5180
rect 115500 5236 115556 5246
rect 115500 5142 115556 5180
rect 116284 5236 116340 5246
rect 116284 5142 116340 5180
rect 115612 5124 115668 5134
rect 114380 4340 114436 5068
rect 114380 4246 114436 4284
rect 114828 5012 114884 5022
rect 114828 4562 114884 4956
rect 114828 4510 114830 4562
rect 114882 4510 114884 4562
rect 114828 4116 114884 4510
rect 115612 4562 115668 5068
rect 116172 5124 116228 5134
rect 116172 5030 116228 5068
rect 115612 4510 115614 4562
rect 115666 4510 115668 4562
rect 115612 4498 115668 4510
rect 116732 4452 116788 5628
rect 116956 5236 117012 5246
rect 116956 5142 117012 5180
rect 116732 4386 116788 4396
rect 114828 4050 114884 4060
rect 117068 4004 117124 4014
rect 115724 3668 115780 3678
rect 115724 3574 115780 3612
rect 114268 3278 114270 3330
rect 114322 3278 114324 3330
rect 114268 3266 114324 3278
rect 115948 3444 116004 3454
rect 115948 800 116004 3388
rect 116508 3444 116564 3454
rect 116508 3350 116564 3388
rect 117068 2996 117124 3948
rect 117180 3668 117236 6300
rect 117292 5908 117348 6414
rect 117852 6130 117908 8372
rect 118300 7588 118356 7598
rect 118188 7364 118244 7374
rect 118188 7270 118244 7308
rect 117852 6078 117854 6130
rect 117906 6078 117908 6130
rect 117852 6066 117908 6078
rect 118300 6130 118356 7532
rect 118300 6078 118302 6130
rect 118354 6078 118356 6130
rect 117516 5908 117572 5918
rect 117292 5906 117572 5908
rect 117292 5854 117518 5906
rect 117570 5854 117572 5906
rect 117292 5852 117572 5854
rect 117516 4116 117572 5852
rect 117852 5236 117908 5246
rect 117740 5012 117796 5022
rect 117740 4918 117796 4956
rect 117180 3554 117236 3612
rect 117180 3502 117182 3554
rect 117234 3502 117236 3554
rect 117180 3490 117236 3502
rect 117292 4060 117572 4116
rect 117068 2930 117124 2940
rect 117292 800 117348 4060
rect 117852 3332 117908 5180
rect 118300 5010 118356 6078
rect 118524 5348 118580 5358
rect 118524 5254 118580 5292
rect 119532 5348 119588 35420
rect 119868 35140 119924 35150
rect 119868 34914 119924 35084
rect 119868 34862 119870 34914
rect 119922 34862 119924 34914
rect 119868 34850 119924 34862
rect 119644 34690 119700 34702
rect 119644 34638 119646 34690
rect 119698 34638 119700 34690
rect 119644 33236 119700 34638
rect 119644 33170 119700 33180
rect 120316 27748 120372 35532
rect 120428 35140 120484 35150
rect 120428 35026 120484 35084
rect 120428 34974 120430 35026
rect 120482 34974 120484 35026
rect 120428 34962 120484 34974
rect 120988 35026 121044 35532
rect 120988 34974 120990 35026
rect 121042 34974 121044 35026
rect 120988 34962 121044 34974
rect 121548 34802 121604 37436
rect 121996 36594 122052 37772
rect 121996 36542 121998 36594
rect 122050 36542 122052 36594
rect 121996 36530 122052 36542
rect 121996 35698 122052 35710
rect 121996 35646 121998 35698
rect 122050 35646 122052 35698
rect 121996 35588 122052 35646
rect 121548 34750 121550 34802
rect 121602 34750 121604 34802
rect 121548 34738 121604 34750
rect 121884 34802 121940 34814
rect 121884 34750 121886 34802
rect 121938 34750 121940 34802
rect 121884 34692 121940 34750
rect 121884 34626 121940 34636
rect 120316 27682 120372 27692
rect 121996 17668 122052 35532
rect 122108 34916 122164 37884
rect 122892 36596 122948 39200
rect 122892 36530 122948 36540
rect 123116 38612 123172 38622
rect 122444 36372 122500 36382
rect 122332 35924 122388 35934
rect 122332 35830 122388 35868
rect 122108 34850 122164 34860
rect 122444 34802 122500 36316
rect 123116 35812 123172 38556
rect 123788 36708 123844 39200
rect 123788 36652 124068 36708
rect 123788 36482 123844 36494
rect 123788 36430 123790 36482
rect 123842 36430 123844 36482
rect 123452 36260 123508 36270
rect 123452 36166 123508 36204
rect 123116 35746 123172 35756
rect 123676 35700 123732 35710
rect 122780 35588 122836 35598
rect 122780 35494 122836 35532
rect 123564 35476 123620 35486
rect 123564 35382 123620 35420
rect 122444 34750 122446 34802
rect 122498 34750 122500 34802
rect 122444 34738 122500 34750
rect 122668 34916 122724 34926
rect 122108 34692 122164 34702
rect 122108 34018 122164 34636
rect 122668 34354 122724 34860
rect 123340 34802 123396 34814
rect 123340 34750 123342 34802
rect 123394 34750 123396 34802
rect 122668 34302 122670 34354
rect 122722 34302 122724 34354
rect 122668 34290 122724 34302
rect 123004 34356 123060 34366
rect 123004 34262 123060 34300
rect 123340 34356 123396 34750
rect 123676 34802 123732 35644
rect 123676 34750 123678 34802
rect 123730 34750 123732 34802
rect 123676 34738 123732 34750
rect 123340 34290 123396 34300
rect 123788 34132 123844 36430
rect 123900 35476 123956 35486
rect 123900 35382 123956 35420
rect 124012 34916 124068 36652
rect 124572 36482 124628 36494
rect 124572 36430 124574 36482
rect 124626 36430 124628 36482
rect 124348 36370 124404 36382
rect 124348 36318 124350 36370
rect 124402 36318 124404 36370
rect 124012 34850 124068 34860
rect 124124 35812 124180 35822
rect 124124 34692 124180 35756
rect 124236 34692 124292 34702
rect 124124 34690 124292 34692
rect 124124 34638 124238 34690
rect 124290 34638 124292 34690
rect 124124 34636 124292 34638
rect 124236 34626 124292 34636
rect 123788 34066 123844 34076
rect 122108 33966 122110 34018
rect 122162 33966 122164 34018
rect 122108 26908 122164 33966
rect 123564 34020 123620 34030
rect 123564 30100 123620 33964
rect 124348 34020 124404 36318
rect 124460 35812 124516 35822
rect 124460 35718 124516 35756
rect 124572 35698 124628 36430
rect 124684 35812 124740 39200
rect 125244 36482 125300 36494
rect 125244 36430 125246 36482
rect 125298 36430 125300 36482
rect 125244 35924 125300 36430
rect 125244 35858 125300 35868
rect 124684 35746 124740 35756
rect 124572 35646 124574 35698
rect 124626 35646 124628 35698
rect 124572 35588 124628 35646
rect 125356 35700 125412 35710
rect 125356 35606 125412 35644
rect 124572 35522 124628 35532
rect 125132 35476 125188 35486
rect 124796 34916 124852 34926
rect 124796 34354 124852 34860
rect 124796 34302 124798 34354
rect 124850 34302 124852 34354
rect 124796 34290 124852 34302
rect 125020 34690 125076 34702
rect 125020 34638 125022 34690
rect 125074 34638 125076 34690
rect 124348 33954 124404 33964
rect 125020 33908 125076 34638
rect 125132 34354 125188 35420
rect 125244 34916 125300 34926
rect 125244 34822 125300 34860
rect 125580 34916 125636 39200
rect 126028 36596 126084 36606
rect 126028 36502 126084 36540
rect 126476 36596 126532 39200
rect 126476 36530 126532 36540
rect 127260 36482 127316 36494
rect 127260 36430 127262 36482
rect 127314 36430 127316 36482
rect 126252 35812 126308 35822
rect 126252 35718 126308 35756
rect 127260 35364 127316 36430
rect 127372 35812 127428 39200
rect 127932 36596 127988 36606
rect 127932 36502 127988 36540
rect 128268 36596 128324 39200
rect 128268 36530 128324 36540
rect 128156 36260 128212 36270
rect 127372 35756 127540 35812
rect 127372 35588 127428 35598
rect 127372 35494 127428 35532
rect 127148 35308 127260 35364
rect 125580 34850 125636 34860
rect 126588 34916 126644 34926
rect 126252 34802 126308 34814
rect 126252 34750 126254 34802
rect 126306 34750 126308 34802
rect 125132 34302 125134 34354
rect 125186 34302 125188 34354
rect 125132 34290 125188 34302
rect 125916 34690 125972 34702
rect 125916 34638 125918 34690
rect 125970 34638 125972 34690
rect 125580 34132 125636 34142
rect 125580 34038 125636 34076
rect 125020 33842 125076 33852
rect 125916 31668 125972 34638
rect 125916 31602 125972 31612
rect 126140 34242 126196 34254
rect 126140 34190 126142 34242
rect 126194 34190 126196 34242
rect 123564 30034 123620 30044
rect 126140 28532 126196 34190
rect 126252 33572 126308 34750
rect 126476 34130 126532 34142
rect 126476 34078 126478 34130
rect 126530 34078 126532 34130
rect 126476 34020 126532 34078
rect 126476 33954 126532 33964
rect 126476 33572 126532 33582
rect 126252 33516 126476 33572
rect 126140 28466 126196 28476
rect 122108 26852 122388 26908
rect 122332 20188 122388 26852
rect 122332 20132 122612 20188
rect 121996 17602 122052 17612
rect 120764 11172 120820 11182
rect 120764 8372 120820 11116
rect 120764 8306 120820 8316
rect 121884 8372 121940 8382
rect 121884 8278 121940 8316
rect 122444 8034 122500 8046
rect 122444 7982 122446 8034
rect 122498 7982 122500 8034
rect 122444 7812 122500 7982
rect 122108 7756 122500 7812
rect 121772 7588 121828 7598
rect 121324 7586 121828 7588
rect 121324 7534 121774 7586
rect 121826 7534 121828 7586
rect 121324 7532 121828 7534
rect 121212 7364 121268 7374
rect 121100 7362 121268 7364
rect 121100 7310 121214 7362
rect 121266 7310 121268 7362
rect 121100 7308 121268 7310
rect 120652 6692 120708 6702
rect 121100 6692 121156 7308
rect 121212 7298 121268 7308
rect 120652 6690 121156 6692
rect 120652 6638 120654 6690
rect 120706 6638 121156 6690
rect 120652 6636 121156 6638
rect 121324 6690 121380 7532
rect 121772 7522 121828 7532
rect 122108 7586 122164 7756
rect 122108 7534 122110 7586
rect 122162 7534 122164 7586
rect 122108 7522 122164 7534
rect 121324 6638 121326 6690
rect 121378 6638 121380 6690
rect 120204 6468 120260 6478
rect 120652 6468 120708 6636
rect 121324 6626 121380 6638
rect 120204 6466 120708 6468
rect 120204 6414 120206 6466
rect 120258 6414 120708 6466
rect 120204 6412 120708 6414
rect 120204 5908 120260 6412
rect 122556 6132 122612 20132
rect 124684 9154 124740 9166
rect 124684 9102 124686 9154
rect 124738 9102 124740 9154
rect 123116 8932 123172 8942
rect 123116 8838 123172 8876
rect 124124 8932 124180 8942
rect 124124 8838 124180 8876
rect 124348 8932 124404 8942
rect 123788 8818 123844 8830
rect 123788 8766 123790 8818
rect 123842 8766 123844 8818
rect 123564 8484 123620 8494
rect 122780 8372 122836 8382
rect 122780 8278 122836 8316
rect 123564 8258 123620 8428
rect 123564 8206 123566 8258
rect 123618 8206 123620 8258
rect 123564 8194 123620 8206
rect 123788 8260 123844 8766
rect 124124 8484 124180 8494
rect 124348 8428 124404 8876
rect 124124 8372 124404 8428
rect 124684 8428 124740 9102
rect 124908 9042 124964 9054
rect 124908 8990 124910 9042
rect 124962 8990 124964 9042
rect 124908 8932 124964 8990
rect 124908 8866 124964 8876
rect 125468 8932 125524 8942
rect 125468 8838 125524 8876
rect 125916 8930 125972 8942
rect 125916 8878 125918 8930
rect 125970 8878 125972 8930
rect 124684 8372 124852 8428
rect 124124 8370 124180 8372
rect 124124 8318 124126 8370
rect 124178 8318 124180 8370
rect 124124 8306 124180 8318
rect 124796 8306 124852 8316
rect 125916 8372 125972 8878
rect 123788 8194 123844 8204
rect 125244 8260 125300 8270
rect 125916 8260 125972 8316
rect 125916 8204 126196 8260
rect 125244 8166 125300 8204
rect 123452 8148 123508 8158
rect 123452 8054 123508 8092
rect 124348 8148 124404 8158
rect 123116 8036 123172 8046
rect 122332 6076 122612 6132
rect 122668 7474 122724 7486
rect 122668 7422 122670 7474
rect 122722 7422 122724 7474
rect 122668 6692 122724 7422
rect 120204 5842 120260 5852
rect 121996 5908 122052 5918
rect 121996 5814 122052 5852
rect 121548 5794 121604 5806
rect 121548 5742 121550 5794
rect 121602 5742 121604 5794
rect 119532 5234 119588 5292
rect 119532 5182 119534 5234
rect 119586 5182 119588 5234
rect 119532 5170 119588 5182
rect 121212 5348 121268 5358
rect 118300 4958 118302 5010
rect 118354 4958 118356 5010
rect 118300 4946 118356 4958
rect 120204 5122 120260 5134
rect 120204 5070 120206 5122
rect 120258 5070 120260 5122
rect 120204 5012 120260 5070
rect 120204 4946 120260 4956
rect 120876 5122 120932 5134
rect 120876 5070 120878 5122
rect 120930 5070 120932 5122
rect 120876 5012 120932 5070
rect 121212 5122 121268 5292
rect 121212 5070 121214 5122
rect 121266 5070 121268 5122
rect 121212 5058 121268 5070
rect 121324 5124 121380 5134
rect 118860 4900 118916 4910
rect 118860 4898 119364 4900
rect 118860 4846 118862 4898
rect 118914 4846 119364 4898
rect 118860 4844 119364 4846
rect 118860 4834 118916 4844
rect 118972 4564 119028 4574
rect 117964 4562 119028 4564
rect 117964 4510 118974 4562
rect 119026 4510 119028 4562
rect 117964 4508 119028 4510
rect 117964 4338 118020 4508
rect 118972 4498 119028 4508
rect 119308 4450 119364 4844
rect 119308 4398 119310 4450
rect 119362 4398 119364 4450
rect 119308 4386 119364 4398
rect 117964 4286 117966 4338
rect 118018 4286 118020 4338
rect 117964 4274 118020 4286
rect 118524 4340 118580 4350
rect 118524 4246 118580 4284
rect 120876 4340 120932 4956
rect 121324 4562 121380 5068
rect 121324 4510 121326 4562
rect 121378 4510 121380 4562
rect 121324 4498 121380 4510
rect 120876 4274 120932 4284
rect 121548 4340 121604 5742
rect 121548 4274 121604 4284
rect 122220 4340 122276 4350
rect 122220 4246 122276 4284
rect 121772 4226 121828 4238
rect 121772 4174 121774 4226
rect 121826 4174 121828 4226
rect 118300 4004 118356 4014
rect 118300 3554 118356 3948
rect 119308 4004 119364 4014
rect 119308 3666 119364 3948
rect 119308 3614 119310 3666
rect 119362 3614 119364 3666
rect 119308 3602 119364 3614
rect 121436 3668 121492 3678
rect 118300 3502 118302 3554
rect 118354 3502 118356 3554
rect 118300 3490 118356 3502
rect 121436 3554 121492 3612
rect 121436 3502 121438 3554
rect 121490 3502 121492 3554
rect 121436 3490 121492 3502
rect 119980 3444 120036 3454
rect 117964 3332 118020 3342
rect 117852 3330 118020 3332
rect 117852 3278 117966 3330
rect 118018 3278 118020 3330
rect 117852 3276 118020 3278
rect 117964 3266 118020 3276
rect 119980 800 120036 3388
rect 120540 3444 120596 3454
rect 120540 3350 120596 3388
rect 121324 3444 121380 3454
rect 121324 800 121380 3388
rect 121772 3444 121828 4174
rect 121772 3378 121828 3388
rect 121996 3444 122052 3454
rect 121996 3350 122052 3388
rect 122332 3330 122388 6076
rect 122444 5908 122500 5918
rect 122668 5908 122724 6636
rect 122500 5852 122724 5908
rect 123116 5906 123172 7980
rect 123340 7924 123396 7934
rect 123340 7474 123396 7868
rect 123340 7422 123342 7474
rect 123394 7422 123396 7474
rect 123340 7410 123396 7422
rect 123116 5854 123118 5906
rect 123170 5854 123172 5906
rect 122444 5814 122500 5852
rect 123116 5842 123172 5854
rect 123340 7140 123396 7150
rect 122892 4340 122948 4350
rect 122892 4246 122948 4284
rect 123340 4338 123396 7084
rect 124348 6914 124404 8092
rect 125020 8036 125076 8046
rect 125020 7942 125076 7980
rect 125916 8036 125972 8046
rect 125916 7812 125972 7980
rect 125916 7746 125972 7756
rect 125804 7700 125860 7710
rect 125804 7606 125860 7644
rect 124348 6862 124350 6914
rect 124402 6862 124404 6914
rect 124348 6850 124404 6862
rect 126140 6916 126196 8204
rect 124908 6692 124964 6702
rect 124908 6598 124964 6636
rect 125468 6690 125524 6702
rect 125468 6638 125470 6690
rect 125522 6638 125524 6690
rect 123788 6468 123844 6478
rect 123788 6374 123844 6412
rect 125244 5908 125300 5918
rect 123900 5348 123956 5358
rect 123788 4898 123844 4910
rect 123788 4846 123790 4898
rect 123842 4846 123844 4898
rect 123788 4564 123844 4846
rect 123788 4498 123844 4508
rect 123340 4286 123342 4338
rect 123394 4286 123396 4338
rect 123340 4274 123396 4286
rect 123340 3668 123396 3678
rect 123340 3574 123396 3612
rect 123788 3668 123844 3678
rect 123900 3668 123956 5292
rect 124348 5236 124404 5246
rect 124348 5142 124404 5180
rect 124908 5124 124964 5134
rect 124908 5030 124964 5068
rect 125244 5124 125300 5852
rect 123788 3666 123956 3668
rect 123788 3614 123790 3666
rect 123842 3614 123956 3666
rect 123788 3612 123956 3614
rect 123788 3602 123844 3612
rect 125244 3554 125300 5068
rect 125468 4788 125524 6638
rect 125580 6132 125636 6142
rect 125580 6038 125636 6076
rect 126140 6130 126196 6860
rect 126252 8034 126308 8046
rect 126252 7982 126254 8034
rect 126306 7982 126308 8034
rect 126252 6692 126308 7982
rect 126364 7252 126420 7262
rect 126364 7158 126420 7196
rect 126252 6626 126308 6636
rect 126140 6078 126142 6130
rect 126194 6078 126196 6130
rect 126140 6066 126196 6078
rect 125804 5684 125860 5694
rect 125468 4722 125524 4732
rect 125692 4898 125748 4910
rect 125692 4846 125694 4898
rect 125746 4846 125748 4898
rect 125692 3780 125748 4846
rect 125804 4562 125860 5628
rect 125804 4510 125806 4562
rect 125858 4510 125860 4562
rect 125804 4498 125860 4510
rect 126364 4228 126420 4238
rect 126364 4134 126420 4172
rect 125692 3714 125748 3724
rect 125244 3502 125246 3554
rect 125298 3502 125300 3554
rect 125244 3490 125300 3502
rect 125356 3556 125412 3566
rect 122332 3278 122334 3330
rect 122386 3278 122388 3330
rect 122332 3266 122388 3278
rect 124012 3444 124068 3454
rect 124012 800 124068 3388
rect 124572 3444 124628 3454
rect 124572 3350 124628 3388
rect 125356 800 125412 3500
rect 126140 3556 126196 3566
rect 126140 3462 126196 3500
rect 126364 3332 126420 3342
rect 126476 3332 126532 33516
rect 126588 33458 126644 34860
rect 127036 34916 127092 34926
rect 127036 34822 127092 34860
rect 126588 33406 126590 33458
rect 126642 33406 126644 33458
rect 126588 33394 126644 33406
rect 126812 34690 126868 34702
rect 126812 34638 126814 34690
rect 126866 34638 126868 34690
rect 126812 33348 126868 34638
rect 126924 34020 126980 34030
rect 126924 33926 126980 33964
rect 127036 33460 127092 33470
rect 127148 33460 127204 35308
rect 127260 35298 127316 35308
rect 127484 34916 127540 35756
rect 127484 34850 127540 34860
rect 127932 35700 127988 35710
rect 127708 34802 127764 34814
rect 127708 34750 127710 34802
rect 127762 34750 127764 34802
rect 127708 34692 127764 34750
rect 127708 34356 127764 34636
rect 127820 34356 127876 34366
rect 127708 34354 127876 34356
rect 127708 34302 127822 34354
rect 127874 34302 127876 34354
rect 127708 34300 127876 34302
rect 127820 34290 127876 34300
rect 127372 34018 127428 34030
rect 127372 33966 127374 34018
rect 127426 33966 127428 34018
rect 127372 33572 127428 33966
rect 127372 33506 127428 33516
rect 127036 33458 127204 33460
rect 127036 33406 127038 33458
rect 127090 33406 127204 33458
rect 127036 33404 127204 33406
rect 127036 33394 127092 33404
rect 126812 33282 126868 33292
rect 127932 26908 127988 35644
rect 128044 35140 128100 35150
rect 128044 34802 128100 35084
rect 128044 34750 128046 34802
rect 128098 34750 128100 34802
rect 128044 34738 128100 34750
rect 128156 32004 128212 36204
rect 129052 35700 129108 35710
rect 129052 35606 129108 35644
rect 128828 34916 128884 34926
rect 128828 34822 128884 34860
rect 128604 34690 128660 34702
rect 128604 34638 128606 34690
rect 128658 34638 128660 34690
rect 128268 34018 128324 34030
rect 128268 33966 128270 34018
rect 128322 33966 128324 34018
rect 128268 33124 128324 33966
rect 128604 33460 128660 34638
rect 129164 34244 129220 39200
rect 130060 37044 130116 39200
rect 129948 36988 130116 37044
rect 130844 37268 130900 37278
rect 129724 36596 129780 36606
rect 129724 36502 129780 36540
rect 129276 36484 129332 36494
rect 129276 36482 129556 36484
rect 129276 36430 129278 36482
rect 129330 36430 129556 36482
rect 129276 36428 129556 36430
rect 129276 36418 129332 36428
rect 129388 34916 129444 34926
rect 129388 34822 129444 34860
rect 129388 34356 129444 34366
rect 129500 34356 129556 36428
rect 129612 36372 129668 36382
rect 129612 35810 129668 36316
rect 129612 35758 129614 35810
rect 129666 35758 129668 35810
rect 129612 35746 129668 35758
rect 129948 34916 130004 36988
rect 130082 36876 130346 36886
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130082 36810 130346 36820
rect 130844 35812 130900 37212
rect 130956 36036 131012 39200
rect 131852 36932 131908 39200
rect 131852 36866 131908 36876
rect 132412 36708 132468 36718
rect 131852 36706 132468 36708
rect 131852 36654 132414 36706
rect 132466 36654 132468 36706
rect 131852 36652 132468 36654
rect 131404 36482 131460 36494
rect 131404 36430 131406 36482
rect 131458 36430 131460 36482
rect 131292 36370 131348 36382
rect 131292 36318 131294 36370
rect 131346 36318 131348 36370
rect 131292 36260 131348 36318
rect 131292 36194 131348 36204
rect 130956 35980 131124 36036
rect 130060 35700 130116 35710
rect 130844 35680 130900 35756
rect 130060 35606 130116 35644
rect 130082 35308 130346 35318
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130082 35242 130346 35252
rect 131068 35252 131124 35980
rect 131404 35810 131460 36430
rect 131404 35758 131406 35810
rect 131458 35758 131460 35810
rect 131068 35186 131124 35196
rect 131292 35700 131348 35710
rect 131068 35026 131124 35038
rect 131068 34974 131070 35026
rect 131122 34974 131124 35026
rect 129948 34850 130004 34860
rect 130508 34916 130564 34926
rect 131068 34916 131124 34974
rect 130508 34914 130676 34916
rect 130508 34862 130510 34914
rect 130562 34862 130676 34914
rect 130508 34860 130676 34862
rect 130508 34850 130564 34860
rect 129388 34354 129556 34356
rect 129388 34302 129390 34354
rect 129442 34302 129556 34354
rect 129388 34300 129556 34302
rect 130284 34356 130340 34366
rect 129388 34290 129444 34300
rect 130284 34262 130340 34300
rect 129164 34178 129220 34188
rect 129052 34130 129108 34142
rect 129052 34078 129054 34130
rect 129106 34078 129108 34130
rect 128604 33394 128660 33404
rect 128716 33572 128772 33582
rect 128716 33458 128772 33516
rect 128716 33406 128718 33458
rect 128770 33406 128772 33458
rect 128716 33394 128772 33406
rect 128268 33058 128324 33068
rect 129052 33124 129108 34078
rect 130060 34130 130116 34142
rect 130060 34078 130062 34130
rect 130114 34078 130116 34130
rect 130060 34020 130116 34078
rect 130060 33908 130116 33964
rect 130060 33852 130564 33908
rect 130082 33740 130346 33750
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130082 33674 130346 33684
rect 129276 33572 129332 33582
rect 129276 33346 129332 33516
rect 129276 33294 129278 33346
rect 129330 33294 129332 33346
rect 129276 33282 129332 33294
rect 129612 33236 129668 33246
rect 129612 33142 129668 33180
rect 129052 33058 129108 33068
rect 130172 33122 130228 33134
rect 130172 33070 130174 33122
rect 130226 33070 130228 33122
rect 130172 33012 130228 33070
rect 130172 32946 130228 32956
rect 130508 33122 130564 33852
rect 130508 33070 130510 33122
rect 130562 33070 130564 33122
rect 130082 32172 130346 32182
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130082 32106 130346 32116
rect 128156 31938 128212 31948
rect 130082 30604 130346 30614
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130082 30538 130346 30548
rect 130082 29036 130346 29046
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130082 28970 130346 28980
rect 130082 27468 130346 27478
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130082 27402 130346 27412
rect 127932 26852 128212 26908
rect 128156 26786 128212 26796
rect 130082 25900 130346 25910
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130082 25834 130346 25844
rect 130082 24332 130346 24342
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130082 24266 130346 24276
rect 130082 22764 130346 22774
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130082 22698 130346 22708
rect 130082 21196 130346 21206
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130082 21130 130346 21140
rect 130082 19628 130346 19638
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130082 19562 130346 19572
rect 130082 18060 130346 18070
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130082 17994 130346 18004
rect 130082 16492 130346 16502
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130082 16426 130346 16436
rect 130082 14924 130346 14934
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130082 14858 130346 14868
rect 130082 13356 130346 13366
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130082 13290 130346 13300
rect 130082 11788 130346 11798
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130082 11722 130346 11732
rect 130082 10220 130346 10230
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130082 10154 130346 10164
rect 130082 8652 130346 8662
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130082 8586 130346 8596
rect 126812 8036 126868 8046
rect 126812 7942 126868 7980
rect 127260 8034 127316 8046
rect 127260 7982 127262 8034
rect 127314 7982 127316 8034
rect 127260 7924 127316 7982
rect 126812 7700 126868 7710
rect 126812 7606 126868 7644
rect 126924 7362 126980 7374
rect 126924 7310 126926 7362
rect 126978 7310 126980 7362
rect 126588 6468 126644 6478
rect 126588 6130 126644 6412
rect 126588 6078 126590 6130
rect 126642 6078 126644 6130
rect 126588 6066 126644 6078
rect 126700 5796 126756 5806
rect 126924 5796 126980 7310
rect 127260 7140 127316 7868
rect 127260 7074 127316 7084
rect 127484 7362 127540 7374
rect 127484 7310 127486 7362
rect 127538 7310 127540 7362
rect 127260 6132 127316 6142
rect 127260 6038 127316 6076
rect 127484 6132 127540 7310
rect 126700 5794 126980 5796
rect 126700 5742 126702 5794
rect 126754 5742 126980 5794
rect 126700 5740 126980 5742
rect 127372 5794 127428 5806
rect 127372 5742 127374 5794
rect 127426 5742 127428 5794
rect 126700 5572 126756 5740
rect 126700 5506 126756 5516
rect 127372 5572 127428 5742
rect 127372 5506 127428 5516
rect 127260 5236 127316 5246
rect 127260 4338 127316 5180
rect 127484 4676 127540 6076
rect 127596 7250 127652 7262
rect 127596 7198 127598 7250
rect 127650 7198 127652 7250
rect 127596 5796 127652 7198
rect 130082 7084 130346 7094
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130082 7018 130346 7028
rect 128044 6466 128100 6478
rect 128044 6414 128046 6466
rect 128098 6414 128100 6466
rect 128044 6020 128100 6414
rect 128044 5954 128100 5964
rect 128380 6468 128436 6478
rect 127596 5730 127652 5740
rect 128044 5794 128100 5806
rect 128044 5742 128046 5794
rect 128098 5742 128100 5794
rect 127932 5684 127988 5694
rect 127932 5590 127988 5628
rect 128044 5572 128100 5742
rect 128044 5506 128100 5516
rect 128044 5122 128100 5134
rect 128044 5070 128046 5122
rect 128098 5070 128100 5122
rect 128044 5012 128100 5070
rect 128044 4946 128100 4956
rect 128380 5122 128436 6412
rect 128604 6466 128660 6478
rect 128604 6414 128606 6466
rect 128658 6414 128660 6466
rect 128604 6356 128660 6414
rect 129052 6468 129108 6478
rect 129388 6468 129444 6478
rect 129052 6466 129220 6468
rect 129052 6414 129054 6466
rect 129106 6414 129220 6466
rect 129052 6412 129220 6414
rect 129052 6402 129108 6412
rect 128604 6290 128660 6300
rect 129164 5908 129220 6412
rect 129388 6374 129444 6412
rect 129388 6132 129444 6142
rect 129388 6038 129444 6076
rect 129164 5906 129332 5908
rect 129164 5854 129166 5906
rect 129218 5854 129332 5906
rect 129164 5852 129332 5854
rect 129164 5842 129220 5852
rect 129276 5796 129332 5852
rect 129836 5796 129892 5806
rect 130284 5796 130340 5806
rect 129276 5794 129892 5796
rect 129276 5742 129838 5794
rect 129890 5742 129892 5794
rect 129276 5740 129892 5742
rect 128380 5070 128382 5122
rect 128434 5070 128436 5122
rect 127260 4286 127262 4338
rect 127314 4286 127316 4338
rect 127260 4274 127316 4286
rect 127372 4620 127484 4676
rect 127260 3780 127316 3790
rect 127260 3686 127316 3724
rect 127372 3666 127428 4620
rect 127484 4610 127540 4620
rect 128156 4676 128212 4686
rect 128044 4564 128100 4574
rect 128044 4470 128100 4508
rect 127484 4452 127540 4462
rect 127484 4358 127540 4396
rect 128156 4450 128212 4620
rect 128156 4398 128158 4450
rect 128210 4398 128212 4450
rect 128156 4386 128212 4398
rect 128380 4340 128436 5070
rect 129052 5572 129108 5582
rect 129052 5010 129108 5516
rect 129052 4958 129054 5010
rect 129106 4958 129108 5010
rect 129052 4946 129108 4958
rect 129276 5122 129332 5740
rect 129836 5730 129892 5740
rect 129948 5794 130340 5796
rect 129948 5742 130286 5794
rect 130338 5742 130340 5794
rect 129948 5740 130340 5742
rect 129948 5572 130004 5740
rect 130284 5730 130340 5740
rect 129836 5516 130004 5572
rect 130082 5516 130346 5526
rect 129276 5070 129278 5122
rect 129330 5070 129332 5122
rect 128380 4274 128436 4284
rect 128940 4340 128996 4350
rect 128940 4246 128996 4284
rect 129276 4004 129332 5070
rect 129276 3938 129332 3948
rect 129388 5124 129444 5134
rect 129388 3780 129444 5068
rect 129500 4452 129556 4462
rect 129500 4338 129556 4396
rect 129500 4286 129502 4338
rect 129554 4286 129556 4338
rect 129500 4274 129556 4286
rect 129500 3780 129556 3790
rect 129388 3724 129500 3780
rect 127372 3614 127374 3666
rect 127426 3614 127428 3666
rect 127372 3602 127428 3614
rect 129500 3554 129556 3724
rect 129500 3502 129502 3554
rect 129554 3502 129556 3554
rect 129500 3490 129556 3502
rect 126364 3330 126532 3332
rect 126364 3278 126366 3330
rect 126418 3278 126532 3330
rect 126364 3276 126532 3278
rect 128044 3444 128100 3454
rect 126364 3266 126420 3276
rect 128044 800 128100 3388
rect 128604 3444 128660 3454
rect 129836 3444 129892 5516
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130082 5450 130346 5460
rect 130284 5124 130340 5134
rect 130284 5010 130340 5068
rect 130284 4958 130286 5010
rect 130338 4958 130340 5010
rect 130284 4946 130340 4958
rect 129948 4898 130004 4910
rect 129948 4846 129950 4898
rect 130002 4846 130004 4898
rect 129948 4788 130004 4846
rect 129948 4722 130004 4732
rect 130082 3948 130346 3958
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130082 3882 130346 3892
rect 130060 3444 130116 3454
rect 129836 3442 130116 3444
rect 129836 3390 130062 3442
rect 130114 3390 130116 3442
rect 129836 3388 130116 3390
rect 128604 3350 128660 3388
rect 129388 924 129668 980
rect 129388 800 129444 924
rect 113596 700 113988 756
rect 114576 0 114688 800
rect 115920 0 116032 800
rect 117264 0 117376 800
rect 118608 0 118720 800
rect 119952 0 120064 800
rect 121296 0 121408 800
rect 122640 0 122752 800
rect 123984 0 124096 800
rect 125328 0 125440 800
rect 126672 0 126784 800
rect 128016 0 128128 800
rect 129360 0 129472 800
rect 129612 756 129668 924
rect 130060 756 130116 3388
rect 130396 3332 130452 3342
rect 130508 3332 130564 33070
rect 130620 33012 130676 34860
rect 131068 34850 131124 34860
rect 131292 34916 131348 35644
rect 131404 35588 131460 35758
rect 131404 35522 131460 35532
rect 131628 35588 131684 35598
rect 131628 35494 131684 35532
rect 131740 35476 131796 35486
rect 131292 34850 131348 34860
rect 131516 35252 131572 35262
rect 130844 34242 130900 34254
rect 130844 34190 130846 34242
rect 130898 34190 130900 34242
rect 130844 34132 130900 34190
rect 130844 34066 130900 34076
rect 131180 34244 131236 34254
rect 131068 33460 131124 33470
rect 131180 33460 131236 34188
rect 131068 33458 131236 33460
rect 131068 33406 131070 33458
rect 131122 33406 131236 33458
rect 131068 33404 131236 33406
rect 131516 33458 131572 35196
rect 131740 34354 131796 35420
rect 131740 34302 131742 34354
rect 131794 34302 131796 34354
rect 131740 34290 131796 34302
rect 131516 33406 131518 33458
rect 131570 33406 131572 33458
rect 131068 33394 131124 33404
rect 131516 33394 131572 33406
rect 130620 32946 130676 32956
rect 130844 6020 130900 6030
rect 130844 5346 130900 5964
rect 130844 5294 130846 5346
rect 130898 5294 130900 5346
rect 130844 5282 130900 5294
rect 131852 5348 131908 36652
rect 132412 36642 132468 36652
rect 132076 36482 132132 36494
rect 132076 36430 132078 36482
rect 132130 36430 132132 36482
rect 132076 35700 132132 36430
rect 132076 35634 132132 35644
rect 132524 35812 132580 35822
rect 131964 35476 132020 35486
rect 131964 35474 132468 35476
rect 131964 35422 131966 35474
rect 132018 35422 132468 35474
rect 131964 35420 132468 35422
rect 131964 35410 132020 35420
rect 132076 35252 132132 35262
rect 131964 34916 132020 34926
rect 131964 34822 132020 34860
rect 132076 34242 132132 35196
rect 132076 34190 132078 34242
rect 132130 34190 132132 34242
rect 132076 34178 132132 34190
rect 132188 6356 132244 6366
rect 131852 5234 131908 5292
rect 131852 5182 131854 5234
rect 131906 5182 131908 5234
rect 131852 5170 131908 5182
rect 131964 5796 132020 5806
rect 130956 5122 131012 5134
rect 130956 5070 130958 5122
rect 131010 5070 131012 5122
rect 130956 4676 131012 5070
rect 130956 4610 131012 4620
rect 131964 4562 132020 5740
rect 132076 5682 132132 5694
rect 132076 5630 132078 5682
rect 132130 5630 132132 5682
rect 132076 5236 132132 5630
rect 132076 5170 132132 5180
rect 132188 5572 132244 6300
rect 132412 6132 132468 35420
rect 132524 34354 132580 35756
rect 132636 35698 132692 35710
rect 132636 35646 132638 35698
rect 132690 35646 132692 35698
rect 132636 34692 132692 35646
rect 132748 34916 132804 39200
rect 133084 36482 133140 36494
rect 133084 36430 133086 36482
rect 133138 36430 133140 36482
rect 132972 35924 133028 35934
rect 133084 35924 133140 36430
rect 132972 35922 133140 35924
rect 132972 35870 132974 35922
rect 133026 35870 133140 35922
rect 132972 35868 133140 35870
rect 132972 35858 133028 35868
rect 133644 35812 133700 39200
rect 133756 36932 133812 36942
rect 133756 36594 133812 36876
rect 133756 36542 133758 36594
rect 133810 36542 133812 36594
rect 133756 36530 133812 36542
rect 133644 35746 133700 35756
rect 132972 35700 133028 35710
rect 132804 34860 132916 34916
rect 132748 34850 132804 34860
rect 132636 34626 132692 34636
rect 132524 34302 132526 34354
rect 132578 34302 132580 34354
rect 132524 34290 132580 34302
rect 132860 34356 132916 34860
rect 132972 34802 133028 35644
rect 133868 35698 133924 35710
rect 133868 35646 133870 35698
rect 133922 35646 133924 35698
rect 133868 35140 133924 35646
rect 134540 35700 134596 39200
rect 135212 38164 135268 38174
rect 134988 36260 135044 36270
rect 134988 36166 135044 36204
rect 134764 35812 134820 35822
rect 134764 35718 134820 35756
rect 134540 35634 134596 35644
rect 133868 35074 133924 35084
rect 133196 34916 133252 34926
rect 133196 34822 133252 34860
rect 132972 34750 132974 34802
rect 133026 34750 133028 34802
rect 132972 34738 133028 34750
rect 134428 34802 134484 34814
rect 134428 34750 134430 34802
rect 134482 34750 134484 34802
rect 133756 34692 133812 34702
rect 133756 34598 133812 34636
rect 132972 34356 133028 34366
rect 132860 34354 133028 34356
rect 132860 34302 132974 34354
rect 133026 34302 133028 34354
rect 132860 34300 133028 34302
rect 132972 34290 133028 34300
rect 134092 34018 134148 34030
rect 134092 33966 134094 34018
rect 134146 33966 134148 34018
rect 132412 5906 132468 6076
rect 133532 33908 133588 33918
rect 132412 5854 132414 5906
rect 132466 5854 132468 5906
rect 132412 5842 132468 5854
rect 132972 6018 133028 6030
rect 132972 5966 132974 6018
rect 133026 5966 133028 6018
rect 132188 5234 132244 5516
rect 132972 5684 133028 5966
rect 133196 5908 133252 5918
rect 133196 5814 133252 5852
rect 132188 5182 132190 5234
rect 132242 5182 132244 5234
rect 132188 5170 132244 5182
rect 132300 5236 132356 5246
rect 131964 4510 131966 4562
rect 132018 4510 132020 4562
rect 131964 4498 132020 4510
rect 131628 3780 131684 3790
rect 131628 3666 131684 3724
rect 132300 3780 132356 5180
rect 132972 5124 133028 5628
rect 133420 5348 133476 5358
rect 133420 5254 133476 5292
rect 132300 3714 132356 3724
rect 132636 5068 133028 5124
rect 133084 5124 133140 5134
rect 132636 4114 132692 5068
rect 133084 5030 133140 5068
rect 133308 4900 133364 4910
rect 132972 4228 133028 4238
rect 132972 4134 133028 4172
rect 133308 4228 133364 4844
rect 133532 4564 133588 33852
rect 134092 33908 134148 33966
rect 134092 33842 134148 33852
rect 134428 33908 134484 34750
rect 134764 34690 134820 34702
rect 134764 34638 134766 34690
rect 134818 34638 134820 34690
rect 134764 34580 134820 34638
rect 134764 34514 134820 34524
rect 135212 34354 135268 38108
rect 135436 35140 135492 39200
rect 135772 38164 135828 38174
rect 135436 35074 135492 35084
rect 135548 36372 135604 36382
rect 135212 34302 135214 34354
rect 135266 34302 135268 34354
rect 135212 34290 135268 34302
rect 135548 34356 135604 36316
rect 135772 36370 135828 38108
rect 136332 36484 136388 39200
rect 137228 36596 137284 39200
rect 137228 36540 137508 36596
rect 136332 36418 136388 36428
rect 136556 36482 136612 36494
rect 136556 36430 136558 36482
rect 136610 36430 136612 36482
rect 135772 36318 135774 36370
rect 135826 36318 135828 36370
rect 135772 36306 135828 36318
rect 136220 36372 136276 36382
rect 136220 36036 136276 36316
rect 136556 36148 136612 36430
rect 136892 36260 136948 36270
rect 137340 36260 137396 36270
rect 136892 36258 137284 36260
rect 136892 36206 136894 36258
rect 136946 36206 137284 36258
rect 136892 36204 137284 36206
rect 136892 36194 136948 36204
rect 136556 36082 136612 36092
rect 136220 35970 136276 35980
rect 137116 36036 137172 36046
rect 135660 35810 135716 35822
rect 135660 35758 135662 35810
rect 135714 35758 135716 35810
rect 135660 35588 135716 35758
rect 135884 35700 135940 35710
rect 135884 35606 135940 35644
rect 136892 35700 136948 35710
rect 136892 35606 136948 35644
rect 135660 35522 135716 35532
rect 136332 35140 136388 35150
rect 136332 35026 136388 35084
rect 136332 34974 136334 35026
rect 136386 34974 136388 35026
rect 136332 34962 136388 34974
rect 135772 34914 135828 34926
rect 135772 34862 135774 34914
rect 135826 34862 135828 34914
rect 135660 34356 135716 34366
rect 135548 34354 135716 34356
rect 135548 34302 135662 34354
rect 135714 34302 135716 34354
rect 135548 34300 135716 34302
rect 135660 34290 135716 34300
rect 134428 33842 134484 33852
rect 135772 33236 135828 34862
rect 137116 34692 137172 35980
rect 137116 34626 137172 34636
rect 135772 33170 135828 33180
rect 135996 34020 136052 34030
rect 135996 30212 136052 33964
rect 135996 30146 136052 30156
rect 136780 8932 136836 8942
rect 135660 7924 135716 7934
rect 135660 6578 135716 7868
rect 135660 6526 135662 6578
rect 135714 6526 135716 6578
rect 135660 6514 135716 6526
rect 135772 7252 135828 7262
rect 135772 6244 135828 7196
rect 136780 6692 136836 8876
rect 137116 8036 137172 8046
rect 137116 7698 137172 7980
rect 137116 7646 137118 7698
rect 137170 7646 137172 7698
rect 137116 7634 137172 7646
rect 135996 6580 136052 6590
rect 135996 6486 136052 6524
rect 136668 6578 136724 6590
rect 136668 6526 136670 6578
rect 136722 6526 136724 6578
rect 136780 6560 136836 6636
rect 134204 6132 134260 6142
rect 134204 6038 134260 6076
rect 135772 6132 135828 6188
rect 135772 6130 135940 6132
rect 135772 6078 135774 6130
rect 135826 6078 135940 6130
rect 135772 6076 135940 6078
rect 135772 6066 135828 6076
rect 133756 5908 133812 5918
rect 133756 5794 133812 5852
rect 133756 5742 133758 5794
rect 133810 5742 133812 5794
rect 133756 5236 133812 5742
rect 134652 5794 134708 5806
rect 134652 5742 134654 5794
rect 134706 5742 134708 5794
rect 134652 5684 134708 5742
rect 134652 5618 134708 5628
rect 135212 5796 135268 5806
rect 133756 5170 133812 5180
rect 133980 5572 134036 5582
rect 133980 5010 134036 5516
rect 134204 5236 134260 5246
rect 134204 5122 134260 5180
rect 134764 5236 134820 5246
rect 134764 5142 134820 5180
rect 135212 5234 135268 5740
rect 135212 5182 135214 5234
rect 135266 5182 135268 5234
rect 135212 5170 135268 5182
rect 134204 5070 134206 5122
rect 134258 5070 134260 5122
rect 134204 5058 134260 5070
rect 133980 4958 133982 5010
rect 134034 4958 134036 5010
rect 133980 4946 134036 4958
rect 135772 5012 135828 5022
rect 135772 4918 135828 4956
rect 133644 4564 133700 4574
rect 133532 4562 133700 4564
rect 133532 4510 133646 4562
rect 133698 4510 133700 4562
rect 133532 4508 133700 4510
rect 133644 4498 133700 4508
rect 132636 4062 132638 4114
rect 132690 4062 132692 4114
rect 131628 3614 131630 3666
rect 131682 3614 131684 3666
rect 131628 3602 131684 3614
rect 132636 3668 132692 4062
rect 132636 3602 132692 3612
rect 131068 3556 131124 3566
rect 131068 3462 131124 3500
rect 133308 3554 133364 4172
rect 133308 3502 133310 3554
rect 133362 3502 133364 3554
rect 133308 3490 133364 3502
rect 133868 4338 133924 4350
rect 133868 4286 133870 4338
rect 133922 4286 133924 4338
rect 133868 4228 133924 4286
rect 130396 3330 130564 3332
rect 130396 3278 130398 3330
rect 130450 3278 130564 3330
rect 130396 3276 130564 3278
rect 132076 3444 132132 3454
rect 130396 3266 130452 3276
rect 132076 800 132132 3388
rect 132636 3444 132692 3454
rect 132636 3350 132692 3388
rect 133868 2884 133924 4172
rect 134428 4228 134484 4238
rect 134428 4134 134484 4172
rect 135884 3666 135940 6076
rect 136220 5796 136276 5806
rect 136668 5796 136724 6526
rect 136220 5794 136724 5796
rect 136220 5742 136222 5794
rect 136274 5742 136724 5794
rect 136220 5740 136724 5742
rect 136220 5236 136276 5740
rect 135996 5180 136276 5236
rect 137004 5460 137060 5470
rect 135996 4900 136052 5180
rect 136108 5012 136164 5022
rect 136780 5012 136836 5022
rect 136108 5010 136836 5012
rect 136108 4958 136110 5010
rect 136162 4958 136782 5010
rect 136834 4958 136836 5010
rect 136108 4956 136836 4958
rect 136108 4946 136164 4956
rect 136780 4946 136836 4956
rect 135996 4834 136052 4844
rect 137004 4564 137060 5404
rect 137116 5348 137172 5358
rect 137228 5348 137284 36204
rect 137340 34354 137396 36204
rect 137452 35252 137508 36540
rect 137788 36484 137844 36494
rect 137788 36390 137844 36428
rect 137564 36258 137620 36270
rect 137564 36206 137566 36258
rect 137618 36206 137620 36258
rect 137564 36148 137620 36206
rect 137564 36082 137620 36092
rect 137900 35924 137956 35934
rect 137900 35830 137956 35868
rect 137676 35700 137732 35710
rect 138124 35700 138180 39200
rect 139020 36708 139076 39200
rect 139916 36708 139972 39200
rect 140588 38724 140644 38734
rect 139916 36652 140084 36708
rect 139020 36642 139076 36652
rect 139244 36482 139300 36494
rect 139244 36430 139246 36482
rect 139298 36430 139300 36482
rect 139132 36372 139188 36382
rect 138908 36370 139188 36372
rect 138908 36318 139134 36370
rect 139186 36318 139188 36370
rect 138908 36316 139188 36318
rect 138572 36036 138628 36046
rect 137676 35698 138404 35700
rect 137676 35646 137678 35698
rect 137730 35646 138404 35698
rect 137676 35644 138404 35646
rect 137676 35634 137732 35644
rect 137452 35186 137508 35196
rect 138124 35252 138180 35262
rect 138124 35026 138180 35196
rect 138124 34974 138126 35026
rect 138178 34974 138180 35026
rect 138124 34962 138180 34974
rect 137340 34302 137342 34354
rect 137394 34302 137396 34354
rect 137340 34290 137396 34302
rect 137452 34914 137508 34926
rect 137452 34862 137454 34914
rect 137506 34862 137508 34914
rect 137452 34356 137508 34862
rect 137452 34290 137508 34300
rect 138348 34242 138404 35644
rect 138572 35698 138628 35980
rect 138572 35646 138574 35698
rect 138626 35646 138628 35698
rect 138572 35634 138628 35646
rect 138684 35810 138740 35822
rect 138684 35758 138686 35810
rect 138738 35758 138740 35810
rect 138348 34190 138350 34242
rect 138402 34190 138404 34242
rect 138348 34178 138404 34190
rect 138012 34018 138068 34030
rect 138012 33966 138014 34018
rect 138066 33966 138068 34018
rect 138012 33906 138068 33966
rect 138012 33854 138014 33906
rect 138066 33854 138068 33906
rect 138012 31892 138068 33854
rect 138684 33906 138740 35758
rect 138908 34354 138964 36316
rect 139132 36306 139188 36316
rect 139132 35028 139188 35038
rect 139244 35028 139300 36430
rect 139916 36482 139972 36494
rect 139916 36430 139918 36482
rect 139970 36430 139972 36482
rect 139916 35924 139972 36430
rect 139916 35858 139972 35868
rect 139356 35476 139412 35486
rect 139356 35382 139412 35420
rect 139692 35474 139748 35486
rect 139692 35422 139694 35474
rect 139746 35422 139748 35474
rect 139132 35026 139412 35028
rect 139132 34974 139134 35026
rect 139186 34974 139412 35026
rect 139132 34972 139412 34974
rect 139132 34692 139188 34972
rect 139132 34626 139188 34636
rect 138908 34302 138910 34354
rect 138962 34302 138964 34354
rect 138908 34020 138964 34302
rect 139356 34354 139412 34972
rect 139356 34302 139358 34354
rect 139410 34302 139412 34354
rect 139356 34290 139412 34302
rect 138908 33954 138964 33964
rect 138684 33854 138686 33906
rect 138738 33854 138740 33906
rect 138684 33842 138740 33854
rect 138012 31826 138068 31836
rect 137564 7700 137620 7710
rect 137340 7474 137396 7486
rect 137340 7422 137342 7474
rect 137394 7422 137396 7474
rect 137340 6132 137396 7422
rect 137452 6916 137508 6926
rect 137564 6916 137620 7644
rect 139132 7700 139188 7710
rect 139132 7606 139188 7644
rect 139692 7700 139748 35422
rect 139804 35476 139860 35486
rect 139804 34802 139860 35420
rect 139804 34750 139806 34802
rect 139858 34750 139860 34802
rect 139804 34738 139860 34750
rect 140028 34914 140084 36652
rect 140028 34862 140030 34914
rect 140082 34862 140084 34914
rect 140028 34356 140084 34862
rect 140028 34290 140084 34300
rect 140252 36258 140308 36270
rect 140252 36206 140254 36258
rect 140306 36206 140308 36258
rect 139916 34018 139972 34030
rect 139916 33966 139918 34018
rect 139970 33966 139972 34018
rect 139916 33906 139972 33966
rect 139916 33854 139918 33906
rect 139970 33854 139972 33906
rect 139916 33842 139972 33854
rect 139692 7634 139748 7644
rect 139916 7812 139972 7822
rect 137452 6914 137620 6916
rect 137452 6862 137454 6914
rect 137506 6862 137620 6914
rect 137452 6860 137620 6862
rect 138124 7362 138180 7374
rect 138124 7310 138126 7362
rect 138178 7310 138180 7362
rect 137452 6850 137508 6860
rect 138124 6692 138180 7310
rect 137788 6580 137844 6590
rect 137788 6486 137844 6524
rect 137340 6066 137396 6076
rect 137452 6244 137508 6254
rect 137452 6020 137508 6188
rect 138012 6020 138068 6030
rect 138124 6020 138180 6636
rect 138684 7362 138740 7374
rect 138684 7310 138686 7362
rect 138738 7310 138740 7362
rect 137452 6018 137620 6020
rect 137452 5966 137454 6018
rect 137506 5966 137620 6018
rect 137452 5964 137620 5966
rect 137452 5954 137508 5964
rect 137116 5346 137228 5348
rect 137116 5294 137118 5346
rect 137170 5294 137228 5346
rect 137116 5292 137228 5294
rect 137116 5282 137172 5292
rect 137228 5216 137284 5292
rect 137452 5124 137508 5134
rect 137116 4564 137172 4574
rect 137004 4562 137172 4564
rect 137004 4510 137118 4562
rect 137170 4510 137172 4562
rect 137004 4508 137172 4510
rect 137116 4498 137172 4508
rect 137452 4450 137508 5068
rect 137452 4398 137454 4450
rect 137506 4398 137508 4450
rect 137452 4386 137508 4398
rect 135884 3614 135886 3666
rect 135938 3614 135940 3666
rect 135884 3602 135940 3614
rect 137564 3554 137620 5964
rect 138012 6018 138180 6020
rect 138012 5966 138014 6018
rect 138066 5966 138180 6018
rect 138012 5964 138180 5966
rect 138012 5954 138068 5964
rect 137900 5908 137956 5918
rect 137788 5460 137844 5470
rect 137788 5236 137844 5404
rect 137788 5122 137844 5180
rect 137788 5070 137790 5122
rect 137842 5070 137844 5122
rect 137788 5058 137844 5070
rect 137900 5010 137956 5852
rect 138124 5908 138180 5964
rect 138124 5842 138180 5852
rect 138460 6580 138516 6590
rect 138236 5682 138292 5694
rect 138236 5630 138238 5682
rect 138290 5630 138292 5682
rect 138236 5236 138292 5630
rect 138236 5170 138292 5180
rect 138460 5460 138516 6524
rect 138684 6578 138740 7310
rect 139356 6804 139412 6814
rect 139356 6710 139412 6748
rect 138684 6526 138686 6578
rect 138738 6526 138740 6578
rect 138572 6132 138628 6142
rect 138572 6038 138628 6076
rect 138684 5572 138740 6526
rect 139132 6580 139188 6590
rect 139132 6486 139188 6524
rect 139692 6466 139748 6478
rect 139692 6414 139694 6466
rect 139746 6414 139748 6466
rect 138684 5506 138740 5516
rect 139020 5908 139076 5918
rect 138460 5234 138516 5404
rect 138460 5182 138462 5234
rect 138514 5182 138516 5234
rect 138460 5170 138516 5182
rect 138796 5348 138852 5358
rect 137900 4958 137902 5010
rect 137954 4958 137956 5010
rect 137900 4946 137956 4958
rect 138348 4564 138404 4574
rect 138348 4470 138404 4508
rect 138796 4562 138852 5292
rect 139020 5234 139076 5852
rect 139580 5908 139636 5918
rect 139580 5814 139636 5852
rect 139020 5182 139022 5234
rect 139074 5182 139076 5234
rect 139020 5170 139076 5182
rect 139468 5236 139524 5246
rect 139468 5142 139524 5180
rect 139692 5124 139748 6414
rect 139804 6020 139860 6030
rect 139804 5234 139860 5964
rect 139804 5182 139806 5234
rect 139858 5182 139860 5234
rect 139804 5170 139860 5182
rect 139692 5058 139748 5068
rect 138796 4510 138798 4562
rect 138850 4510 138852 4562
rect 138796 4498 138852 4510
rect 137564 3502 137566 3554
rect 137618 3502 137620 3554
rect 137564 3490 137620 3502
rect 138012 4338 138068 4350
rect 138012 4286 138014 4338
rect 138066 4286 138068 4338
rect 138012 3666 138068 4286
rect 138012 3614 138014 3666
rect 138066 3614 138068 3666
rect 133420 2828 133924 2884
rect 136108 3444 136164 3454
rect 133420 800 133476 2828
rect 136108 800 136164 3388
rect 136668 3444 136724 3454
rect 136668 3350 136724 3388
rect 137452 3444 137508 3454
rect 137452 800 137508 3388
rect 138012 3444 138068 3614
rect 139916 3668 139972 7756
rect 140252 6804 140308 36206
rect 140476 36036 140532 36046
rect 140476 35698 140532 35980
rect 140476 35646 140478 35698
rect 140530 35646 140532 35698
rect 140476 35634 140532 35646
rect 140588 35810 140644 38668
rect 140812 36596 140868 39200
rect 140812 36530 140868 36540
rect 140924 37044 140980 37054
rect 140588 35758 140590 35810
rect 140642 35758 140644 35810
rect 140364 34356 140420 34366
rect 140364 34262 140420 34300
rect 140588 33906 140644 35758
rect 140924 34914 140980 36988
rect 141596 36708 141652 36718
rect 141596 36594 141652 36652
rect 141596 36542 141598 36594
rect 141650 36542 141652 36594
rect 141596 36530 141652 36542
rect 140924 34862 140926 34914
rect 140978 34862 140980 34914
rect 140812 34356 140868 34366
rect 140924 34356 140980 34862
rect 141036 36482 141092 36494
rect 141036 36430 141038 36482
rect 141090 36430 141092 36482
rect 141036 34580 141092 36430
rect 141708 35812 141764 39200
rect 142156 36036 142212 36046
rect 142156 35922 142212 35980
rect 142156 35870 142158 35922
rect 142210 35870 142212 35922
rect 142156 35858 142212 35870
rect 142604 35924 142660 39200
rect 142604 35858 142660 35868
rect 142940 36482 142996 36494
rect 142940 36430 142942 36482
rect 142994 36430 142996 36482
rect 141484 35756 141764 35812
rect 141260 35588 141316 35626
rect 141260 35522 141316 35532
rect 141260 35364 141316 35374
rect 141260 34802 141316 35308
rect 141260 34750 141262 34802
rect 141314 34750 141316 34802
rect 141260 34738 141316 34750
rect 141036 34514 141092 34524
rect 140812 34354 140980 34356
rect 140812 34302 140814 34354
rect 140866 34302 140980 34354
rect 140812 34300 140980 34302
rect 140812 34290 140868 34300
rect 140588 33854 140590 33906
rect 140642 33854 140644 33906
rect 140588 33842 140644 33854
rect 140252 6738 140308 6748
rect 140812 6804 140868 6814
rect 140812 6690 140868 6748
rect 140812 6638 140814 6690
rect 140866 6638 140868 6690
rect 140812 6626 140868 6638
rect 140140 6020 140196 6030
rect 140140 5926 140196 5964
rect 140700 6020 140756 6030
rect 140700 5236 140756 5964
rect 140812 5236 140868 5246
rect 140700 5234 140868 5236
rect 140700 5182 140814 5234
rect 140866 5182 140868 5234
rect 140700 5180 140868 5182
rect 140812 5170 140868 5180
rect 140924 4564 140980 34300
rect 141484 34354 141540 35756
rect 142828 35700 142884 35710
rect 142492 35698 142884 35700
rect 142492 35646 142830 35698
rect 142882 35646 142884 35698
rect 142492 35644 142884 35646
rect 141932 35588 141988 35598
rect 141484 34302 141486 34354
rect 141538 34302 141540 34354
rect 141484 34244 141540 34302
rect 141484 34178 141540 34188
rect 141596 35474 141652 35486
rect 141596 35422 141598 35474
rect 141650 35422 141652 35474
rect 141260 6580 141316 6590
rect 141260 6466 141316 6524
rect 141260 6414 141262 6466
rect 141314 6414 141316 6466
rect 141260 6018 141316 6414
rect 141260 5966 141262 6018
rect 141314 5966 141316 6018
rect 141260 5954 141316 5966
rect 141596 5236 141652 35422
rect 141932 34354 141988 35532
rect 141932 34302 141934 34354
rect 141986 34302 141988 34354
rect 141932 34290 141988 34302
rect 142156 34804 142212 34814
rect 142156 31948 142212 34748
rect 142492 34802 142548 35644
rect 142828 35634 142884 35644
rect 142940 35364 142996 36430
rect 142940 35298 142996 35308
rect 143500 34916 143556 39200
rect 143612 36596 143668 36606
rect 143612 36502 143668 36540
rect 144396 36596 144452 39200
rect 144396 36530 144452 36540
rect 144956 36482 145012 36494
rect 144956 36430 144958 36482
rect 145010 36430 145012 36482
rect 143724 35924 143780 35934
rect 143724 35810 143780 35868
rect 144956 35922 145012 36430
rect 144956 35870 144958 35922
rect 145010 35870 145012 35922
rect 144956 35858 145012 35870
rect 145292 35924 145348 39200
rect 145852 37604 145908 37614
rect 145404 36596 145460 36606
rect 145404 36502 145460 36540
rect 145292 35858 145348 35868
rect 145852 35922 145908 37548
rect 148492 36092 148756 36102
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148492 36026 148756 36036
rect 145852 35870 145854 35922
rect 145906 35870 145908 35922
rect 145852 35858 145908 35870
rect 146188 35924 146244 35934
rect 143724 35758 143726 35810
rect 143778 35758 143780 35810
rect 143724 35746 143780 35758
rect 146188 35810 146244 35868
rect 146636 35924 146692 35934
rect 146636 35830 146692 35868
rect 146188 35758 146190 35810
rect 146242 35758 146244 35810
rect 146188 35746 146244 35758
rect 145180 35698 145236 35710
rect 145180 35646 145182 35698
rect 145234 35646 145236 35698
rect 145180 35028 145236 35646
rect 145180 34962 145236 34972
rect 145516 35028 145572 35038
rect 142492 34750 142494 34802
rect 142546 34750 142548 34802
rect 142492 34738 142548 34750
rect 142940 34804 142996 34814
rect 142940 34710 142996 34748
rect 143500 34354 143556 34860
rect 143948 34916 144004 34926
rect 143948 34822 144004 34860
rect 143500 34302 143502 34354
rect 143554 34302 143556 34354
rect 143500 34290 143556 34302
rect 143724 34690 143780 34702
rect 143724 34638 143726 34690
rect 143778 34638 143780 34690
rect 142268 34244 142324 34254
rect 142268 34150 142324 34188
rect 141596 5170 141652 5180
rect 142044 31892 142212 31948
rect 140924 4498 140980 4508
rect 142044 4562 142100 31892
rect 143724 31780 143780 34638
rect 145516 31948 145572 34972
rect 148492 34524 148756 34534
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148492 34458 148756 34468
rect 148492 32956 148756 32966
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148492 32890 148756 32900
rect 145516 31892 145796 31948
rect 143724 31714 143780 31724
rect 142044 4510 142046 4562
rect 142098 4510 142100 4562
rect 142044 4498 142100 4510
rect 143948 6916 144004 6926
rect 141708 4338 141764 4350
rect 141708 4286 141710 4338
rect 141762 4286 141764 4338
rect 141260 4228 141316 4238
rect 141708 4228 141764 4286
rect 141260 4226 141764 4228
rect 141260 4174 141262 4226
rect 141314 4174 141764 4226
rect 141260 4172 141764 4174
rect 141260 4162 141316 4172
rect 139916 3666 140420 3668
rect 139916 3614 139918 3666
rect 139970 3614 140420 3666
rect 139916 3612 140420 3614
rect 139916 3602 139972 3612
rect 140364 3554 140420 3612
rect 140364 3502 140366 3554
rect 140418 3502 140420 3554
rect 140364 3490 140420 3502
rect 138012 3378 138068 3388
rect 140140 3444 140196 3454
rect 140140 800 140196 3388
rect 141260 3444 141316 3454
rect 141260 3350 141316 3388
rect 141484 800 141540 4172
rect 143948 3668 144004 6860
rect 145740 4562 145796 31892
rect 148492 31388 148756 31398
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148492 31322 148756 31332
rect 148492 29820 148756 29830
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148492 29754 148756 29764
rect 148492 28252 148756 28262
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148492 28186 148756 28196
rect 148492 26684 148756 26694
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148492 26618 148756 26628
rect 148492 25116 148756 25126
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148492 25050 148756 25060
rect 148492 23548 148756 23558
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148492 23482 148756 23492
rect 148492 21980 148756 21990
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148492 21914 148756 21924
rect 148492 20412 148756 20422
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148492 20346 148756 20356
rect 148492 18844 148756 18854
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148492 18778 148756 18788
rect 148492 17276 148756 17286
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148492 17210 148756 17220
rect 148492 15708 148756 15718
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148492 15642 148756 15652
rect 148492 14140 148756 14150
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148492 14074 148756 14084
rect 148492 12572 148756 12582
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148492 12506 148756 12516
rect 148492 11004 148756 11014
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148492 10938 148756 10948
rect 148492 9436 148756 9446
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148492 9370 148756 9380
rect 148492 7868 148756 7878
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148492 7802 148756 7812
rect 148492 6300 148756 6310
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148492 6234 148756 6244
rect 148492 4732 148756 4742
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148492 4666 148756 4676
rect 145740 4510 145742 4562
rect 145794 4510 145796 4562
rect 145740 4498 145796 4510
rect 145964 4338 146020 4350
rect 145964 4286 145966 4338
rect 146018 4286 146020 4338
rect 145292 4228 145348 4238
rect 145964 4228 146020 4286
rect 145292 4226 146020 4228
rect 145292 4174 145294 4226
rect 145346 4174 146020 4226
rect 145292 4172 146020 4174
rect 145292 4162 145348 4172
rect 143948 3666 144452 3668
rect 143948 3614 143950 3666
rect 144002 3614 144452 3666
rect 143948 3612 144452 3614
rect 143948 3602 144004 3612
rect 144396 3554 144452 3612
rect 144396 3502 144398 3554
rect 144450 3502 144452 3554
rect 144396 3490 144452 3502
rect 144172 3444 144228 3454
rect 144172 800 144228 3388
rect 145292 3444 145348 3454
rect 145292 3350 145348 3388
rect 145516 800 145572 4172
rect 148492 3164 148756 3174
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148492 3098 148756 3108
rect 129612 700 130116 756
rect 130704 0 130816 800
rect 132048 0 132160 800
rect 133392 0 133504 800
rect 134736 0 134848 800
rect 136080 0 136192 800
rect 137424 0 137536 800
rect 138768 0 138880 800
rect 140112 0 140224 800
rect 141456 0 141568 800
rect 142800 0 142912 800
rect 144144 0 144256 800
rect 145488 0 145600 800
<< via2 >>
rect 6076 35922 6132 35924
rect 6076 35870 6078 35922
rect 6078 35870 6130 35922
rect 6130 35870 6132 35922
rect 6076 35868 6132 35870
rect 8876 37100 8932 37156
rect 6972 35868 7028 35924
rect 6412 35756 6468 35812
rect 7532 35810 7588 35812
rect 7532 35758 7534 35810
rect 7534 35758 7586 35810
rect 7586 35758 7588 35810
rect 7532 35756 7588 35758
rect 6188 34914 6244 34916
rect 6188 34862 6190 34914
rect 6190 34862 6242 34914
rect 6242 34862 6244 34914
rect 6188 34860 6244 34862
rect 6972 34914 7028 34916
rect 6972 34862 6974 34914
rect 6974 34862 7026 34914
rect 7026 34862 7028 34914
rect 6972 34860 7028 34862
rect 7868 35084 7924 35140
rect 8764 35532 8820 35588
rect 8988 36428 9044 36484
rect 8876 35084 8932 35140
rect 9772 36482 9828 36484
rect 9772 36430 9774 36482
rect 9774 36430 9826 36482
rect 9826 36430 9828 36482
rect 9772 36428 9828 36430
rect 10892 35980 10948 36036
rect 11788 35980 11844 36036
rect 9660 35586 9716 35588
rect 9660 35534 9662 35586
rect 9662 35534 9714 35586
rect 9714 35534 9716 35586
rect 9660 35532 9716 35534
rect 9100 35084 9156 35140
rect 10108 35084 10164 35140
rect 10332 34972 10388 35028
rect 11004 35026 11060 35028
rect 11004 34974 11006 35026
rect 11006 34974 11058 35026
rect 11058 34974 11060 35026
rect 11004 34972 11060 34974
rect 8540 34412 8596 34468
rect 8876 34412 8932 34468
rect 8764 34242 8820 34244
rect 8764 34190 8766 34242
rect 8766 34190 8818 34242
rect 8818 34190 8820 34242
rect 8764 34188 8820 34190
rect 7868 7532 7924 7588
rect 9660 34412 9716 34468
rect 11004 34300 11060 34356
rect 11116 34748 11172 34804
rect 12012 35644 12068 35700
rect 13244 35810 13300 35812
rect 13244 35758 13246 35810
rect 13246 35758 13298 35810
rect 13298 35758 13300 35810
rect 13244 35756 13300 35758
rect 13804 35756 13860 35812
rect 12908 34914 12964 34916
rect 12908 34862 12910 34914
rect 12910 34862 12962 34914
rect 12962 34862 12964 34914
rect 12908 34860 12964 34862
rect 13580 34914 13636 34916
rect 13580 34862 13582 34914
rect 13582 34862 13634 34914
rect 13634 34862 13636 34914
rect 13580 34860 13636 34862
rect 14588 34914 14644 34916
rect 14588 34862 14590 34914
rect 14590 34862 14642 34914
rect 14642 34862 14644 34914
rect 14588 34860 14644 34862
rect 13020 33964 13076 34020
rect 13468 34018 13524 34020
rect 13468 33966 13470 34018
rect 13470 33966 13522 34018
rect 13522 33966 13524 34018
rect 13468 33964 13524 33966
rect 14252 31052 14308 31108
rect 8876 5180 8932 5236
rect 7756 5122 7812 5124
rect 7756 5070 7758 5122
rect 7758 5070 7810 5122
rect 7810 5070 7812 5122
rect 7756 5068 7812 5070
rect 5852 4732 5908 4788
rect 6188 4732 6244 4788
rect 7756 4450 7812 4452
rect 7756 4398 7758 4450
rect 7758 4398 7810 4450
rect 7810 4398 7812 4450
rect 7756 4396 7812 4398
rect 6972 4338 7028 4340
rect 6972 4286 6974 4338
rect 6974 4286 7026 4338
rect 7026 4286 7028 4338
rect 6972 4284 7028 4286
rect 5852 3554 5908 3556
rect 5852 3502 5854 3554
rect 5854 3502 5906 3554
rect 5906 3502 5908 3554
rect 5852 3500 5908 3502
rect 6300 3442 6356 3444
rect 6300 3390 6302 3442
rect 6302 3390 6354 3442
rect 6354 3390 6356 3442
rect 6300 3388 6356 3390
rect 8316 3612 8372 3668
rect 8540 3836 8596 3892
rect 7308 3554 7364 3556
rect 7308 3502 7310 3554
rect 7310 3502 7362 3554
rect 7362 3502 7364 3554
rect 7308 3500 7364 3502
rect 8428 3500 8484 3556
rect 6524 3388 6580 3444
rect 7084 3388 7140 3444
rect 6636 3330 6692 3332
rect 6636 3278 6638 3330
rect 6638 3278 6690 3330
rect 6690 3278 6692 3330
rect 6636 3276 6692 3278
rect 7532 2940 7588 2996
rect 8764 3612 8820 3668
rect 8652 3276 8708 3332
rect 8988 4338 9044 4340
rect 8988 4286 8990 4338
rect 8990 4286 9042 4338
rect 9042 4286 9044 4338
rect 8988 4284 9044 4286
rect 8988 3836 9044 3892
rect 9884 5068 9940 5124
rect 9772 3836 9828 3892
rect 9996 3612 10052 3668
rect 8876 3276 8932 3332
rect 9772 3388 9828 3444
rect 10220 4396 10276 4452
rect 10444 3724 10500 3780
rect 10108 3388 10164 3444
rect 10332 3442 10388 3444
rect 10332 3390 10334 3442
rect 10334 3390 10386 3442
rect 10386 3390 10388 3442
rect 10332 3388 10388 3390
rect 11116 3388 11172 3444
rect 11676 5068 11732 5124
rect 12124 5010 12180 5012
rect 12124 4958 12126 5010
rect 12126 4958 12178 5010
rect 12178 4958 12180 5010
rect 12124 4956 12180 4958
rect 12684 4956 12740 5012
rect 11340 4898 11396 4900
rect 11340 4846 11342 4898
rect 11342 4846 11394 4898
rect 11394 4846 11396 4898
rect 11340 4844 11396 4846
rect 12348 4396 12404 4452
rect 12236 3778 12292 3780
rect 12236 3726 12238 3778
rect 12238 3726 12290 3778
rect 12290 3726 12292 3778
rect 12236 3724 12292 3726
rect 13692 4956 13748 5012
rect 13356 4732 13412 4788
rect 14812 34860 14868 34916
rect 15820 37324 15876 37380
rect 16044 36594 16100 36596
rect 16044 36542 16046 36594
rect 16046 36542 16098 36594
rect 16098 36542 16100 36594
rect 16044 36540 16100 36542
rect 15484 34690 15540 34692
rect 15484 34638 15486 34690
rect 15486 34638 15538 34690
rect 15538 34638 15540 34690
rect 15484 34636 15540 34638
rect 15820 34860 15876 34916
rect 17164 36540 17220 36596
rect 17500 36370 17556 36372
rect 17500 36318 17502 36370
rect 17502 36318 17554 36370
rect 17554 36318 17556 36370
rect 17500 36316 17556 36318
rect 17500 34188 17556 34244
rect 18172 36316 18228 36372
rect 18284 35420 18340 35476
rect 17836 34188 17892 34244
rect 17052 33180 17108 33236
rect 18956 35644 19012 35700
rect 18620 33516 18676 33572
rect 18396 33404 18452 33460
rect 18284 32732 18340 32788
rect 16492 29372 16548 29428
rect 18172 9324 18228 9380
rect 14588 9212 14644 9268
rect 15708 7532 15764 7588
rect 14588 6466 14644 6468
rect 14588 6414 14590 6466
rect 14590 6414 14642 6466
rect 14642 6414 14644 6466
rect 14588 6412 14644 6414
rect 14252 4844 14308 4900
rect 15036 5180 15092 5236
rect 12684 4396 12740 4452
rect 12908 4396 12964 4452
rect 14476 4226 14532 4228
rect 14476 4174 14478 4226
rect 14478 4174 14530 4226
rect 14530 4174 14532 4226
rect 14476 4172 14532 4174
rect 14924 4060 14980 4116
rect 11676 3442 11732 3444
rect 11676 3390 11678 3442
rect 11678 3390 11730 3442
rect 11730 3390 11732 3442
rect 11676 3388 11732 3390
rect 13804 3388 13860 3444
rect 11340 3330 11396 3332
rect 11340 3278 11342 3330
rect 11342 3278 11394 3330
rect 11394 3278 11396 3330
rect 11340 3276 11396 3278
rect 11228 3164 11284 3220
rect 14364 3442 14420 3444
rect 14364 3390 14366 3442
rect 14366 3390 14418 3442
rect 14418 3390 14420 3442
rect 14364 3388 14420 3390
rect 15372 4508 15428 4564
rect 15484 6412 15540 6468
rect 15036 3276 15092 3332
rect 15148 4172 15204 4228
rect 16156 6130 16212 6132
rect 16156 6078 16158 6130
rect 16158 6078 16210 6130
rect 16210 6078 16212 6130
rect 16156 6076 16212 6078
rect 18284 6690 18340 6692
rect 18284 6638 18286 6690
rect 18286 6638 18338 6690
rect 18338 6638 18340 6690
rect 18284 6636 18340 6638
rect 17612 6076 17668 6132
rect 18732 6412 18788 6468
rect 17724 5964 17780 6020
rect 15932 5906 15988 5908
rect 15932 5854 15934 5906
rect 15934 5854 15986 5906
rect 15986 5854 15988 5906
rect 15932 5852 15988 5854
rect 16716 5740 16772 5796
rect 17500 5740 17556 5796
rect 17276 5122 17332 5124
rect 17276 5070 17278 5122
rect 17278 5070 17330 5122
rect 17330 5070 17332 5122
rect 17276 5068 17332 5070
rect 16940 4732 16996 4788
rect 16156 4396 16212 4452
rect 16268 4620 16324 4676
rect 16828 4450 16884 4452
rect 16828 4398 16830 4450
rect 16830 4398 16882 4450
rect 16882 4398 16884 4450
rect 16828 4396 16884 4398
rect 16268 4284 16324 4340
rect 16940 4226 16996 4228
rect 16940 4174 16942 4226
rect 16942 4174 16994 4226
rect 16994 4174 16996 4226
rect 16940 4172 16996 4174
rect 16492 4060 16548 4116
rect 15932 3442 15988 3444
rect 15932 3390 15934 3442
rect 15934 3390 15986 3442
rect 15986 3390 15988 3442
rect 15932 3388 15988 3390
rect 17836 5906 17892 5908
rect 17836 5854 17838 5906
rect 17838 5854 17890 5906
rect 17890 5854 17892 5906
rect 17836 5852 17892 5854
rect 18172 5906 18228 5908
rect 18172 5854 18174 5906
rect 18174 5854 18226 5906
rect 18226 5854 18228 5906
rect 18172 5852 18228 5854
rect 19622 36874 19678 36876
rect 19622 36822 19624 36874
rect 19624 36822 19676 36874
rect 19676 36822 19678 36874
rect 19622 36820 19678 36822
rect 19726 36874 19782 36876
rect 19726 36822 19728 36874
rect 19728 36822 19780 36874
rect 19780 36822 19782 36874
rect 19726 36820 19782 36822
rect 19830 36874 19886 36876
rect 19830 36822 19832 36874
rect 19832 36822 19884 36874
rect 19884 36822 19886 36874
rect 19830 36820 19886 36822
rect 19516 36370 19572 36372
rect 19516 36318 19518 36370
rect 19518 36318 19570 36370
rect 19570 36318 19572 36370
rect 19516 36316 19572 36318
rect 20188 36316 20244 36372
rect 19740 36092 19796 36148
rect 19404 35420 19460 35476
rect 19622 35306 19678 35308
rect 19622 35254 19624 35306
rect 19624 35254 19676 35306
rect 19676 35254 19678 35306
rect 19622 35252 19678 35254
rect 19726 35306 19782 35308
rect 19726 35254 19728 35306
rect 19728 35254 19780 35306
rect 19780 35254 19782 35306
rect 19726 35252 19782 35254
rect 19830 35306 19886 35308
rect 19830 35254 19832 35306
rect 19832 35254 19884 35306
rect 19884 35254 19886 35306
rect 19830 35252 19886 35254
rect 19292 34860 19348 34916
rect 19516 34748 19572 34804
rect 19622 33738 19678 33740
rect 19622 33686 19624 33738
rect 19624 33686 19676 33738
rect 19676 33686 19678 33738
rect 19622 33684 19678 33686
rect 19726 33738 19782 33740
rect 19726 33686 19728 33738
rect 19728 33686 19780 33738
rect 19780 33686 19782 33738
rect 19726 33684 19782 33686
rect 19830 33738 19886 33740
rect 19830 33686 19832 33738
rect 19832 33686 19884 33738
rect 19884 33686 19886 33738
rect 19830 33684 19886 33686
rect 19852 33516 19908 33572
rect 19292 33458 19348 33460
rect 19292 33406 19294 33458
rect 19294 33406 19346 33458
rect 19346 33406 19348 33458
rect 19292 33404 19348 33406
rect 19852 33068 19908 33124
rect 19622 32170 19678 32172
rect 19622 32118 19624 32170
rect 19624 32118 19676 32170
rect 19676 32118 19678 32170
rect 19622 32116 19678 32118
rect 19726 32170 19782 32172
rect 19726 32118 19728 32170
rect 19728 32118 19780 32170
rect 19780 32118 19782 32170
rect 19726 32116 19782 32118
rect 19830 32170 19886 32172
rect 19830 32118 19832 32170
rect 19832 32118 19884 32170
rect 19884 32118 19886 32170
rect 19830 32116 19886 32118
rect 19292 31164 19348 31220
rect 19622 30602 19678 30604
rect 19622 30550 19624 30602
rect 19624 30550 19676 30602
rect 19676 30550 19678 30602
rect 19622 30548 19678 30550
rect 19726 30602 19782 30604
rect 19726 30550 19728 30602
rect 19728 30550 19780 30602
rect 19780 30550 19782 30602
rect 19726 30548 19782 30550
rect 19830 30602 19886 30604
rect 19830 30550 19832 30602
rect 19832 30550 19884 30602
rect 19884 30550 19886 30602
rect 19830 30548 19886 30550
rect 19622 29034 19678 29036
rect 19622 28982 19624 29034
rect 19624 28982 19676 29034
rect 19676 28982 19678 29034
rect 19622 28980 19678 28982
rect 19726 29034 19782 29036
rect 19726 28982 19728 29034
rect 19728 28982 19780 29034
rect 19780 28982 19782 29034
rect 19726 28980 19782 28982
rect 19830 29034 19886 29036
rect 19830 28982 19832 29034
rect 19832 28982 19884 29034
rect 19884 28982 19886 29034
rect 19830 28980 19886 28982
rect 19622 27466 19678 27468
rect 19622 27414 19624 27466
rect 19624 27414 19676 27466
rect 19676 27414 19678 27466
rect 19622 27412 19678 27414
rect 19726 27466 19782 27468
rect 19726 27414 19728 27466
rect 19728 27414 19780 27466
rect 19780 27414 19782 27466
rect 19726 27412 19782 27414
rect 19830 27466 19886 27468
rect 19830 27414 19832 27466
rect 19832 27414 19884 27466
rect 19884 27414 19886 27466
rect 19830 27412 19886 27414
rect 19622 25898 19678 25900
rect 19622 25846 19624 25898
rect 19624 25846 19676 25898
rect 19676 25846 19678 25898
rect 19622 25844 19678 25846
rect 19726 25898 19782 25900
rect 19726 25846 19728 25898
rect 19728 25846 19780 25898
rect 19780 25846 19782 25898
rect 19726 25844 19782 25846
rect 19830 25898 19886 25900
rect 19830 25846 19832 25898
rect 19832 25846 19884 25898
rect 19884 25846 19886 25898
rect 19830 25844 19886 25846
rect 19622 24330 19678 24332
rect 19622 24278 19624 24330
rect 19624 24278 19676 24330
rect 19676 24278 19678 24330
rect 19622 24276 19678 24278
rect 19726 24330 19782 24332
rect 19726 24278 19728 24330
rect 19728 24278 19780 24330
rect 19780 24278 19782 24330
rect 19726 24276 19782 24278
rect 19830 24330 19886 24332
rect 19830 24278 19832 24330
rect 19832 24278 19884 24330
rect 19884 24278 19886 24330
rect 19830 24276 19886 24278
rect 19622 22762 19678 22764
rect 19622 22710 19624 22762
rect 19624 22710 19676 22762
rect 19676 22710 19678 22762
rect 19622 22708 19678 22710
rect 19726 22762 19782 22764
rect 19726 22710 19728 22762
rect 19728 22710 19780 22762
rect 19780 22710 19782 22762
rect 19726 22708 19782 22710
rect 19830 22762 19886 22764
rect 19830 22710 19832 22762
rect 19832 22710 19884 22762
rect 19884 22710 19886 22762
rect 19830 22708 19886 22710
rect 19622 21194 19678 21196
rect 19622 21142 19624 21194
rect 19624 21142 19676 21194
rect 19676 21142 19678 21194
rect 19622 21140 19678 21142
rect 19726 21194 19782 21196
rect 19726 21142 19728 21194
rect 19728 21142 19780 21194
rect 19780 21142 19782 21194
rect 19726 21140 19782 21142
rect 19830 21194 19886 21196
rect 19830 21142 19832 21194
rect 19832 21142 19884 21194
rect 19884 21142 19886 21194
rect 19830 21140 19886 21142
rect 19622 19626 19678 19628
rect 19622 19574 19624 19626
rect 19624 19574 19676 19626
rect 19676 19574 19678 19626
rect 19622 19572 19678 19574
rect 19726 19626 19782 19628
rect 19726 19574 19728 19626
rect 19728 19574 19780 19626
rect 19780 19574 19782 19626
rect 19726 19572 19782 19574
rect 19830 19626 19886 19628
rect 19830 19574 19832 19626
rect 19832 19574 19884 19626
rect 19884 19574 19886 19626
rect 19830 19572 19886 19574
rect 19622 18058 19678 18060
rect 19622 18006 19624 18058
rect 19624 18006 19676 18058
rect 19676 18006 19678 18058
rect 19622 18004 19678 18006
rect 19726 18058 19782 18060
rect 19726 18006 19728 18058
rect 19728 18006 19780 18058
rect 19780 18006 19782 18058
rect 19726 18004 19782 18006
rect 19830 18058 19886 18060
rect 19830 18006 19832 18058
rect 19832 18006 19884 18058
rect 19884 18006 19886 18058
rect 19830 18004 19886 18006
rect 19622 16490 19678 16492
rect 19622 16438 19624 16490
rect 19624 16438 19676 16490
rect 19676 16438 19678 16490
rect 19622 16436 19678 16438
rect 19726 16490 19782 16492
rect 19726 16438 19728 16490
rect 19728 16438 19780 16490
rect 19780 16438 19782 16490
rect 19726 16436 19782 16438
rect 19830 16490 19886 16492
rect 19830 16438 19832 16490
rect 19832 16438 19884 16490
rect 19884 16438 19886 16490
rect 19830 16436 19886 16438
rect 19622 14922 19678 14924
rect 19622 14870 19624 14922
rect 19624 14870 19676 14922
rect 19676 14870 19678 14922
rect 19622 14868 19678 14870
rect 19726 14922 19782 14924
rect 19726 14870 19728 14922
rect 19728 14870 19780 14922
rect 19780 14870 19782 14922
rect 19726 14868 19782 14870
rect 19830 14922 19886 14924
rect 19830 14870 19832 14922
rect 19832 14870 19884 14922
rect 19884 14870 19886 14922
rect 19830 14868 19886 14870
rect 19622 13354 19678 13356
rect 19622 13302 19624 13354
rect 19624 13302 19676 13354
rect 19676 13302 19678 13354
rect 19622 13300 19678 13302
rect 19726 13354 19782 13356
rect 19726 13302 19728 13354
rect 19728 13302 19780 13354
rect 19780 13302 19782 13354
rect 19726 13300 19782 13302
rect 19830 13354 19886 13356
rect 19830 13302 19832 13354
rect 19832 13302 19884 13354
rect 19884 13302 19886 13354
rect 19830 13300 19886 13302
rect 19622 11786 19678 11788
rect 19622 11734 19624 11786
rect 19624 11734 19676 11786
rect 19676 11734 19678 11786
rect 19622 11732 19678 11734
rect 19726 11786 19782 11788
rect 19726 11734 19728 11786
rect 19728 11734 19780 11786
rect 19780 11734 19782 11786
rect 19726 11732 19782 11734
rect 19830 11786 19886 11788
rect 19830 11734 19832 11786
rect 19832 11734 19884 11786
rect 19884 11734 19886 11786
rect 19830 11732 19886 11734
rect 19622 10218 19678 10220
rect 19622 10166 19624 10218
rect 19624 10166 19676 10218
rect 19676 10166 19678 10218
rect 19622 10164 19678 10166
rect 19726 10218 19782 10220
rect 19726 10166 19728 10218
rect 19728 10166 19780 10218
rect 19780 10166 19782 10218
rect 19726 10164 19782 10166
rect 19830 10218 19886 10220
rect 19830 10166 19832 10218
rect 19832 10166 19884 10218
rect 19884 10166 19886 10218
rect 19830 10164 19886 10166
rect 19622 8650 19678 8652
rect 19622 8598 19624 8650
rect 19624 8598 19676 8650
rect 19676 8598 19678 8650
rect 19622 8596 19678 8598
rect 19726 8650 19782 8652
rect 19726 8598 19728 8650
rect 19728 8598 19780 8650
rect 19780 8598 19782 8650
rect 19726 8596 19782 8598
rect 19830 8650 19886 8652
rect 19830 8598 19832 8650
rect 19832 8598 19884 8650
rect 19884 8598 19886 8650
rect 19830 8596 19886 8598
rect 19292 7362 19348 7364
rect 19292 7310 19294 7362
rect 19294 7310 19346 7362
rect 19346 7310 19348 7362
rect 19292 7308 19348 7310
rect 19622 7082 19678 7084
rect 19622 7030 19624 7082
rect 19624 7030 19676 7082
rect 19676 7030 19678 7082
rect 19622 7028 19678 7030
rect 19726 7082 19782 7084
rect 19726 7030 19728 7082
rect 19728 7030 19780 7082
rect 19780 7030 19782 7082
rect 19726 7028 19782 7030
rect 19830 7082 19886 7084
rect 19830 7030 19832 7082
rect 19832 7030 19884 7082
rect 19884 7030 19886 7082
rect 19830 7028 19886 7030
rect 19628 6914 19684 6916
rect 19628 6862 19630 6914
rect 19630 6862 19682 6914
rect 19682 6862 19684 6914
rect 19628 6860 19684 6862
rect 20076 35308 20132 35364
rect 20076 34300 20132 34356
rect 20076 33628 20132 33684
rect 20412 35810 20468 35812
rect 20412 35758 20414 35810
rect 20414 35758 20466 35810
rect 20466 35758 20468 35810
rect 20412 35756 20468 35758
rect 20748 35308 20804 35364
rect 20300 34860 20356 34916
rect 21644 36540 21700 36596
rect 22204 36594 22260 36596
rect 22204 36542 22206 36594
rect 22206 36542 22258 36594
rect 22258 36542 22260 36594
rect 22204 36540 22260 36542
rect 22092 35308 22148 35364
rect 20412 34242 20468 34244
rect 20412 34190 20414 34242
rect 20414 34190 20466 34242
rect 20466 34190 20468 34242
rect 20412 34188 20468 34190
rect 21308 33852 21364 33908
rect 21756 33852 21812 33908
rect 20636 33628 20692 33684
rect 21756 33628 21812 33684
rect 20300 32396 20356 32452
rect 20300 7362 20356 7364
rect 20300 7310 20302 7362
rect 20302 7310 20354 7362
rect 20354 7310 20356 7362
rect 20300 7308 20356 7310
rect 19964 6860 20020 6916
rect 20524 6860 20580 6916
rect 18844 5852 18900 5908
rect 19628 6018 19684 6020
rect 19628 5966 19630 6018
rect 19630 5966 19682 6018
rect 19682 5966 19684 6018
rect 19628 5964 19684 5966
rect 21532 5906 21588 5908
rect 21532 5854 21534 5906
rect 21534 5854 21586 5906
rect 21586 5854 21588 5906
rect 21532 5852 21588 5854
rect 19622 5514 19678 5516
rect 19622 5462 19624 5514
rect 19624 5462 19676 5514
rect 19676 5462 19678 5514
rect 19622 5460 19678 5462
rect 19726 5514 19782 5516
rect 19726 5462 19728 5514
rect 19728 5462 19780 5514
rect 19780 5462 19782 5514
rect 19726 5460 19782 5462
rect 19830 5514 19886 5516
rect 19830 5462 19832 5514
rect 19832 5462 19884 5514
rect 19884 5462 19886 5514
rect 19830 5460 19886 5462
rect 19068 5292 19124 5348
rect 20300 5404 20356 5460
rect 20300 4844 20356 4900
rect 17612 4338 17668 4340
rect 17612 4286 17614 4338
rect 17614 4286 17666 4338
rect 17666 4286 17668 4338
rect 17612 4284 17668 4286
rect 17948 4284 18004 4340
rect 17612 3836 17668 3892
rect 18172 4172 18228 4228
rect 18732 4508 18788 4564
rect 20300 4172 20356 4228
rect 20748 5346 20804 5348
rect 20748 5294 20750 5346
rect 20750 5294 20802 5346
rect 20802 5294 20804 5346
rect 20748 5292 20804 5294
rect 20412 4396 20468 4452
rect 19622 3946 19678 3948
rect 19622 3894 19624 3946
rect 19624 3894 19676 3946
rect 19676 3894 19678 3946
rect 19622 3892 19678 3894
rect 19726 3946 19782 3948
rect 19726 3894 19728 3946
rect 19728 3894 19780 3946
rect 19780 3894 19782 3946
rect 19726 3892 19782 3894
rect 19830 3946 19886 3948
rect 19830 3894 19832 3946
rect 19832 3894 19884 3946
rect 19884 3894 19886 3946
rect 19830 3892 19886 3894
rect 18844 3442 18900 3444
rect 18844 3390 18846 3442
rect 18846 3390 18898 3442
rect 18898 3390 18900 3442
rect 18844 3388 18900 3390
rect 16716 3330 16772 3332
rect 16716 3278 16718 3330
rect 16718 3278 16770 3330
rect 16770 3278 16772 3330
rect 16716 3276 16772 3278
rect 20412 3612 20468 3668
rect 20524 4284 20580 4340
rect 20636 4172 20692 4228
rect 21532 5122 21588 5124
rect 21532 5070 21534 5122
rect 21534 5070 21586 5122
rect 21586 5070 21588 5122
rect 21532 5068 21588 5070
rect 23100 38444 23156 38500
rect 24220 36092 24276 36148
rect 23436 35532 23492 35588
rect 23100 35196 23156 35252
rect 23996 35308 24052 35364
rect 24332 35586 24388 35588
rect 24332 35534 24334 35586
rect 24334 35534 24386 35586
rect 24386 35534 24388 35586
rect 24332 35532 24388 35534
rect 22876 34524 22932 34580
rect 23324 34412 23380 34468
rect 22428 33740 22484 33796
rect 25788 36764 25844 36820
rect 25676 35420 25732 35476
rect 26572 37548 26628 37604
rect 25900 35420 25956 35476
rect 25452 34300 25508 34356
rect 24892 34076 24948 34132
rect 25004 34188 25060 34244
rect 25564 34130 25620 34132
rect 25564 34078 25566 34130
rect 25566 34078 25618 34130
rect 25618 34078 25620 34130
rect 25564 34076 25620 34078
rect 25004 30940 25060 30996
rect 25116 31164 25172 31220
rect 24332 25676 24388 25732
rect 25116 25564 25172 25620
rect 26236 35420 26292 35476
rect 27804 36594 27860 36596
rect 27804 36542 27806 36594
rect 27806 36542 27858 36594
rect 27858 36542 27860 36594
rect 27804 36540 27860 36542
rect 28364 37212 28420 37268
rect 26012 34354 26068 34356
rect 26012 34302 26014 34354
rect 26014 34302 26066 34354
rect 26066 34302 26068 34354
rect 26012 34300 26068 34302
rect 28140 34802 28196 34804
rect 28140 34750 28142 34802
rect 28142 34750 28194 34802
rect 28194 34750 28196 34802
rect 28140 34748 28196 34750
rect 28812 36540 28868 36596
rect 28476 36482 28532 36484
rect 28476 36430 28478 36482
rect 28478 36430 28530 36482
rect 28530 36430 28532 36482
rect 28476 36428 28532 36430
rect 29596 36428 29652 36484
rect 29372 35698 29428 35700
rect 29372 35646 29374 35698
rect 29374 35646 29426 35698
rect 29426 35646 29428 35698
rect 29372 35644 29428 35646
rect 28700 34748 28756 34804
rect 28700 34300 28756 34356
rect 27132 33516 27188 33572
rect 28364 33068 28420 33124
rect 26908 29372 26964 29428
rect 28364 27580 28420 27636
rect 26908 26460 26964 26516
rect 27804 26460 27860 26516
rect 25116 5122 25172 5124
rect 25116 5070 25118 5122
rect 25118 5070 25170 5122
rect 25170 5070 25172 5122
rect 25116 5068 25172 5070
rect 22092 4338 22148 4340
rect 22092 4286 22094 4338
rect 22094 4286 22146 4338
rect 22146 4286 22148 4338
rect 22092 4284 22148 4286
rect 22540 4338 22596 4340
rect 22540 4286 22542 4338
rect 22542 4286 22594 4338
rect 22594 4286 22596 4338
rect 22540 4284 22596 4286
rect 25004 4226 25060 4228
rect 25004 4174 25006 4226
rect 25006 4174 25058 4226
rect 25058 4174 25060 4226
rect 25004 4172 25060 4174
rect 24556 3388 24612 3444
rect 23772 3164 23828 3220
rect 25676 4060 25732 4116
rect 25900 4172 25956 4228
rect 25676 3442 25732 3444
rect 25676 3390 25678 3442
rect 25678 3390 25730 3442
rect 25730 3390 25732 3442
rect 25676 3388 25732 3390
rect 25116 3164 25172 3220
rect 26460 9212 26516 9268
rect 26572 7532 26628 7588
rect 26684 7474 26740 7476
rect 26684 7422 26686 7474
rect 26686 7422 26738 7474
rect 26738 7422 26740 7474
rect 26684 7420 26740 7422
rect 27244 7586 27300 7588
rect 27244 7534 27246 7586
rect 27246 7534 27298 7586
rect 27298 7534 27300 7586
rect 27244 7532 27300 7534
rect 26908 7308 26964 7364
rect 27132 7196 27188 7252
rect 27692 6636 27748 6692
rect 27356 6466 27412 6468
rect 27356 6414 27358 6466
rect 27358 6414 27410 6466
rect 27410 6414 27412 6466
rect 27356 6412 27412 6414
rect 27692 5964 27748 6020
rect 26572 5180 26628 5236
rect 27132 4508 27188 4564
rect 27468 4450 27524 4452
rect 27468 4398 27470 4450
rect 27470 4398 27522 4450
rect 27522 4398 27524 4450
rect 27468 4396 27524 4398
rect 27244 4060 27300 4116
rect 26236 3276 26292 3332
rect 28028 8034 28084 8036
rect 28028 7982 28030 8034
rect 28030 7982 28082 8034
rect 28082 7982 28084 8034
rect 28028 7980 28084 7982
rect 29372 34860 29428 34916
rect 29036 34636 29092 34692
rect 30156 37772 30212 37828
rect 30156 36706 30212 36708
rect 30156 36654 30158 36706
rect 30158 36654 30210 36706
rect 30210 36654 30212 36706
rect 30156 36652 30212 36654
rect 29708 35532 29764 35588
rect 29932 34914 29988 34916
rect 29932 34862 29934 34914
rect 29934 34862 29986 34914
rect 29986 34862 29988 34914
rect 29932 34860 29988 34862
rect 30156 34636 30212 34692
rect 30044 33404 30100 33460
rect 31724 36652 31780 36708
rect 30604 35084 30660 35140
rect 31500 35586 31556 35588
rect 31500 35534 31502 35586
rect 31502 35534 31554 35586
rect 31554 35534 31556 35586
rect 31500 35532 31556 35534
rect 31388 35084 31444 35140
rect 31836 36428 31892 36484
rect 32172 36482 32228 36484
rect 32172 36430 32174 36482
rect 32174 36430 32226 36482
rect 32226 36430 32228 36482
rect 32172 36428 32228 36430
rect 32396 35756 32452 35812
rect 32620 35644 32676 35700
rect 30604 33458 30660 33460
rect 30604 33406 30606 33458
rect 30606 33406 30658 33458
rect 30658 33406 30660 33458
rect 30604 33404 30660 33406
rect 31052 33458 31108 33460
rect 31052 33406 31054 33458
rect 31054 33406 31106 33458
rect 31106 33406 31108 33458
rect 31052 33404 31108 33406
rect 31164 33292 31220 33348
rect 28924 7980 28980 8036
rect 28028 7420 28084 7476
rect 28588 7474 28644 7476
rect 28588 7422 28590 7474
rect 28590 7422 28642 7474
rect 28642 7422 28644 7474
rect 28588 7420 28644 7422
rect 28364 7308 28420 7364
rect 28252 7250 28308 7252
rect 28252 7198 28254 7250
rect 28254 7198 28306 7250
rect 28306 7198 28308 7250
rect 28252 7196 28308 7198
rect 28812 7308 28868 7364
rect 27916 6524 27972 6580
rect 28252 6412 28308 6468
rect 32844 34914 32900 34916
rect 32844 34862 32846 34914
rect 32846 34862 32898 34914
rect 32898 34862 32900 34914
rect 32844 34860 32900 34862
rect 33852 36988 33908 37044
rect 33516 36540 33572 36596
rect 35084 36540 35140 36596
rect 36092 36594 36148 36596
rect 36092 36542 36094 36594
rect 36094 36542 36146 36594
rect 36146 36542 36148 36594
rect 36092 36540 36148 36542
rect 34524 35810 34580 35812
rect 34524 35758 34526 35810
rect 34526 35758 34578 35810
rect 34578 35758 34580 35810
rect 34524 35756 34580 35758
rect 33292 34860 33348 34916
rect 34188 33628 34244 33684
rect 36316 35868 36372 35924
rect 34524 33964 34580 34020
rect 33068 31836 33124 31892
rect 32620 26348 32676 26404
rect 32396 9212 32452 9268
rect 33516 9324 33572 9380
rect 30380 7474 30436 7476
rect 30380 7422 30382 7474
rect 30382 7422 30434 7474
rect 30434 7422 30436 7474
rect 30380 7420 30436 7422
rect 29932 7362 29988 7364
rect 29932 7310 29934 7362
rect 29934 7310 29986 7362
rect 29986 7310 29988 7362
rect 29932 7308 29988 7310
rect 29596 6578 29652 6580
rect 29596 6526 29598 6578
rect 29598 6526 29650 6578
rect 29650 6526 29652 6578
rect 29596 6524 29652 6526
rect 29372 6188 29428 6244
rect 31388 6188 31444 6244
rect 27916 5404 27972 5460
rect 29708 5346 29764 5348
rect 29708 5294 29710 5346
rect 29710 5294 29762 5346
rect 29762 5294 29764 5346
rect 29708 5292 29764 5294
rect 30604 5292 30660 5348
rect 28588 5234 28644 5236
rect 28588 5182 28590 5234
rect 28590 5182 28642 5234
rect 28642 5182 28644 5234
rect 28588 5180 28644 5182
rect 28700 5068 28756 5124
rect 29596 4844 29652 4900
rect 29148 4562 29204 4564
rect 29148 4510 29150 4562
rect 29150 4510 29202 4562
rect 29202 4510 29204 4562
rect 29148 4508 29204 4510
rect 28140 4450 28196 4452
rect 28140 4398 28142 4450
rect 28142 4398 28194 4450
rect 28194 4398 28196 4450
rect 28140 4396 28196 4398
rect 30156 4898 30212 4900
rect 30156 4846 30158 4898
rect 30158 4846 30210 4898
rect 30210 4846 30212 4898
rect 30156 4844 30212 4846
rect 29596 4450 29652 4452
rect 29596 4398 29598 4450
rect 29598 4398 29650 4450
rect 29650 4398 29652 4450
rect 29596 4396 29652 4398
rect 29148 4060 29204 4116
rect 31724 6018 31780 6020
rect 31724 5966 31726 6018
rect 31726 5966 31778 6018
rect 31778 5966 31780 6018
rect 31724 5964 31780 5966
rect 28588 3442 28644 3444
rect 28588 3390 28590 3442
rect 28590 3390 28642 3442
rect 28642 3390 28644 3442
rect 28588 3388 28644 3390
rect 29596 3442 29652 3444
rect 29596 3390 29598 3442
rect 29598 3390 29650 3442
rect 29650 3390 29652 3442
rect 29596 3388 29652 3390
rect 29932 3388 29988 3444
rect 29260 3330 29316 3332
rect 29260 3278 29262 3330
rect 29262 3278 29314 3330
rect 29314 3278 29316 3330
rect 29260 3276 29316 3278
rect 30492 3442 30548 3444
rect 30492 3390 30494 3442
rect 30494 3390 30546 3442
rect 30546 3390 30548 3442
rect 30492 3388 30548 3390
rect 31276 3388 31332 3444
rect 31836 3388 31892 3444
rect 32620 3388 32676 3444
rect 32284 3164 32340 3220
rect 32956 3388 33012 3444
rect 33180 3442 33236 3444
rect 33180 3390 33182 3442
rect 33182 3390 33234 3442
rect 33234 3390 33236 3442
rect 33180 3388 33236 3390
rect 35084 34018 35140 34020
rect 35084 33966 35086 34018
rect 35086 33966 35138 34018
rect 35138 33966 35140 34018
rect 35084 33964 35140 33966
rect 34860 29148 34916 29204
rect 38444 36482 38500 36484
rect 38444 36430 38446 36482
rect 38446 36430 38498 36482
rect 38498 36430 38500 36482
rect 38444 36428 38500 36430
rect 38032 36090 38088 36092
rect 38032 36038 38034 36090
rect 38034 36038 38086 36090
rect 38086 36038 38088 36090
rect 38032 36036 38088 36038
rect 38136 36090 38192 36092
rect 38136 36038 38138 36090
rect 38138 36038 38190 36090
rect 38190 36038 38192 36090
rect 38136 36036 38192 36038
rect 38240 36090 38296 36092
rect 38240 36038 38242 36090
rect 38242 36038 38294 36090
rect 38294 36038 38296 36090
rect 38240 36036 38296 36038
rect 39004 38332 39060 38388
rect 37548 35532 37604 35588
rect 38108 35586 38164 35588
rect 38108 35534 38110 35586
rect 38110 35534 38162 35586
rect 38162 35534 38164 35586
rect 38108 35532 38164 35534
rect 37772 34914 37828 34916
rect 37772 34862 37774 34914
rect 37774 34862 37826 34914
rect 37826 34862 37828 34914
rect 37772 34860 37828 34862
rect 39116 36428 39172 36484
rect 38332 34914 38388 34916
rect 38332 34862 38334 34914
rect 38334 34862 38386 34914
rect 38386 34862 38388 34914
rect 38332 34860 38388 34862
rect 38032 34522 38088 34524
rect 38032 34470 38034 34522
rect 38034 34470 38086 34522
rect 38086 34470 38088 34522
rect 38032 34468 38088 34470
rect 38136 34522 38192 34524
rect 38136 34470 38138 34522
rect 38138 34470 38190 34522
rect 38190 34470 38192 34522
rect 38136 34468 38192 34470
rect 38240 34522 38296 34524
rect 38240 34470 38242 34522
rect 38242 34470 38294 34522
rect 38294 34470 38296 34522
rect 38240 34468 38296 34470
rect 37548 34076 37604 34132
rect 36764 32508 36820 32564
rect 37436 33740 37492 33796
rect 36316 29260 36372 29316
rect 36092 11564 36148 11620
rect 36316 4172 36372 4228
rect 37212 4226 37268 4228
rect 37212 4174 37214 4226
rect 37214 4174 37266 4226
rect 37266 4174 37268 4226
rect 37212 4172 37268 4174
rect 37772 33180 37828 33236
rect 38556 33740 38612 33796
rect 38332 33180 38388 33236
rect 37996 33122 38052 33124
rect 37996 33070 37998 33122
rect 37998 33070 38050 33122
rect 38050 33070 38052 33122
rect 37996 33068 38052 33070
rect 38032 32954 38088 32956
rect 38032 32902 38034 32954
rect 38034 32902 38086 32954
rect 38086 32902 38088 32954
rect 38032 32900 38088 32902
rect 38136 32954 38192 32956
rect 38136 32902 38138 32954
rect 38138 32902 38190 32954
rect 38190 32902 38192 32954
rect 38136 32900 38192 32902
rect 38240 32954 38296 32956
rect 38240 32902 38242 32954
rect 38242 32902 38294 32954
rect 38294 32902 38296 32954
rect 38240 32900 38296 32902
rect 40236 36482 40292 36484
rect 40236 36430 40238 36482
rect 40238 36430 40290 36482
rect 40290 36430 40292 36482
rect 40236 36428 40292 36430
rect 41804 36764 41860 36820
rect 40908 36428 40964 36484
rect 39900 35810 39956 35812
rect 39900 35758 39902 35810
rect 39902 35758 39954 35810
rect 39954 35758 39956 35810
rect 39900 35756 39956 35758
rect 39340 35532 39396 35588
rect 39116 33740 39172 33796
rect 38668 33180 38724 33236
rect 38556 32844 38612 32900
rect 38032 31386 38088 31388
rect 38032 31334 38034 31386
rect 38034 31334 38086 31386
rect 38086 31334 38088 31386
rect 38032 31332 38088 31334
rect 38136 31386 38192 31388
rect 38136 31334 38138 31386
rect 38138 31334 38190 31386
rect 38190 31334 38192 31386
rect 38136 31332 38192 31334
rect 38240 31386 38296 31388
rect 38240 31334 38242 31386
rect 38242 31334 38294 31386
rect 38294 31334 38296 31386
rect 38240 31332 38296 31334
rect 38032 29818 38088 29820
rect 38032 29766 38034 29818
rect 38034 29766 38086 29818
rect 38086 29766 38088 29818
rect 38032 29764 38088 29766
rect 38136 29818 38192 29820
rect 38136 29766 38138 29818
rect 38138 29766 38190 29818
rect 38190 29766 38192 29818
rect 38136 29764 38192 29766
rect 38240 29818 38296 29820
rect 38240 29766 38242 29818
rect 38242 29766 38294 29818
rect 38294 29766 38296 29818
rect 38240 29764 38296 29766
rect 38032 28250 38088 28252
rect 38032 28198 38034 28250
rect 38034 28198 38086 28250
rect 38086 28198 38088 28250
rect 38032 28196 38088 28198
rect 38136 28250 38192 28252
rect 38136 28198 38138 28250
rect 38138 28198 38190 28250
rect 38190 28198 38192 28250
rect 38136 28196 38192 28198
rect 38240 28250 38296 28252
rect 38240 28198 38242 28250
rect 38242 28198 38294 28250
rect 38294 28198 38296 28250
rect 38240 28196 38296 28198
rect 38032 26682 38088 26684
rect 38032 26630 38034 26682
rect 38034 26630 38086 26682
rect 38086 26630 38088 26682
rect 38032 26628 38088 26630
rect 38136 26682 38192 26684
rect 38136 26630 38138 26682
rect 38138 26630 38190 26682
rect 38190 26630 38192 26682
rect 38136 26628 38192 26630
rect 38240 26682 38296 26684
rect 38240 26630 38242 26682
rect 38242 26630 38294 26682
rect 38294 26630 38296 26682
rect 38240 26628 38296 26630
rect 38032 25114 38088 25116
rect 38032 25062 38034 25114
rect 38034 25062 38086 25114
rect 38086 25062 38088 25114
rect 38032 25060 38088 25062
rect 38136 25114 38192 25116
rect 38136 25062 38138 25114
rect 38138 25062 38190 25114
rect 38190 25062 38192 25114
rect 38136 25060 38192 25062
rect 38240 25114 38296 25116
rect 38240 25062 38242 25114
rect 38242 25062 38294 25114
rect 38294 25062 38296 25114
rect 38240 25060 38296 25062
rect 38032 23546 38088 23548
rect 38032 23494 38034 23546
rect 38034 23494 38086 23546
rect 38086 23494 38088 23546
rect 38032 23492 38088 23494
rect 38136 23546 38192 23548
rect 38136 23494 38138 23546
rect 38138 23494 38190 23546
rect 38190 23494 38192 23546
rect 38136 23492 38192 23494
rect 38240 23546 38296 23548
rect 38240 23494 38242 23546
rect 38242 23494 38294 23546
rect 38294 23494 38296 23546
rect 38240 23492 38296 23494
rect 38032 21978 38088 21980
rect 38032 21926 38034 21978
rect 38034 21926 38086 21978
rect 38086 21926 38088 21978
rect 38032 21924 38088 21926
rect 38136 21978 38192 21980
rect 38136 21926 38138 21978
rect 38138 21926 38190 21978
rect 38190 21926 38192 21978
rect 38136 21924 38192 21926
rect 38240 21978 38296 21980
rect 38240 21926 38242 21978
rect 38242 21926 38294 21978
rect 38294 21926 38296 21978
rect 38240 21924 38296 21926
rect 38032 20410 38088 20412
rect 38032 20358 38034 20410
rect 38034 20358 38086 20410
rect 38086 20358 38088 20410
rect 38032 20356 38088 20358
rect 38136 20410 38192 20412
rect 38136 20358 38138 20410
rect 38138 20358 38190 20410
rect 38190 20358 38192 20410
rect 38136 20356 38192 20358
rect 38240 20410 38296 20412
rect 38240 20358 38242 20410
rect 38242 20358 38294 20410
rect 38294 20358 38296 20410
rect 38240 20356 38296 20358
rect 39564 35532 39620 35588
rect 39452 27244 39508 27300
rect 40796 35420 40852 35476
rect 41132 35756 41188 35812
rect 40684 33852 40740 33908
rect 40348 32284 40404 32340
rect 41804 35756 41860 35812
rect 43372 36428 43428 36484
rect 43260 36316 43316 36372
rect 42588 35868 42644 35924
rect 41132 28364 41188 28420
rect 42588 34412 42644 34468
rect 39900 22876 39956 22932
rect 41244 20972 41300 21028
rect 43932 35810 43988 35812
rect 43932 35758 43934 35810
rect 43934 35758 43986 35810
rect 43986 35758 43988 35810
rect 43932 35756 43988 35758
rect 44156 36482 44212 36484
rect 44156 36430 44158 36482
rect 44158 36430 44210 36482
rect 44210 36430 44212 36482
rect 44156 36428 44212 36430
rect 45724 36876 45780 36932
rect 45724 36316 45780 36372
rect 45276 36258 45332 36260
rect 45276 36206 45278 36258
rect 45278 36206 45330 36258
rect 45330 36206 45332 36258
rect 45276 36204 45332 36206
rect 44380 35420 44436 35476
rect 41916 33852 41972 33908
rect 38032 18842 38088 18844
rect 38032 18790 38034 18842
rect 38034 18790 38086 18842
rect 38086 18790 38088 18842
rect 38032 18788 38088 18790
rect 38136 18842 38192 18844
rect 38136 18790 38138 18842
rect 38138 18790 38190 18842
rect 38190 18790 38192 18842
rect 38136 18788 38192 18790
rect 38240 18842 38296 18844
rect 38240 18790 38242 18842
rect 38242 18790 38294 18842
rect 38294 18790 38296 18842
rect 38240 18788 38296 18790
rect 38032 17274 38088 17276
rect 38032 17222 38034 17274
rect 38034 17222 38086 17274
rect 38086 17222 38088 17274
rect 38032 17220 38088 17222
rect 38136 17274 38192 17276
rect 38136 17222 38138 17274
rect 38138 17222 38190 17274
rect 38190 17222 38192 17274
rect 38136 17220 38192 17222
rect 38240 17274 38296 17276
rect 38240 17222 38242 17274
rect 38242 17222 38294 17274
rect 38294 17222 38296 17274
rect 38240 17220 38296 17222
rect 38032 15706 38088 15708
rect 38032 15654 38034 15706
rect 38034 15654 38086 15706
rect 38086 15654 38088 15706
rect 38032 15652 38088 15654
rect 38136 15706 38192 15708
rect 38136 15654 38138 15706
rect 38138 15654 38190 15706
rect 38190 15654 38192 15706
rect 38136 15652 38192 15654
rect 38240 15706 38296 15708
rect 38240 15654 38242 15706
rect 38242 15654 38294 15706
rect 38294 15654 38296 15706
rect 38240 15652 38296 15654
rect 38032 14138 38088 14140
rect 38032 14086 38034 14138
rect 38034 14086 38086 14138
rect 38086 14086 38088 14138
rect 38032 14084 38088 14086
rect 38136 14138 38192 14140
rect 38136 14086 38138 14138
rect 38138 14086 38190 14138
rect 38190 14086 38192 14138
rect 38136 14084 38192 14086
rect 38240 14138 38296 14140
rect 38240 14086 38242 14138
rect 38242 14086 38294 14138
rect 38294 14086 38296 14138
rect 38240 14084 38296 14086
rect 38032 12570 38088 12572
rect 38032 12518 38034 12570
rect 38034 12518 38086 12570
rect 38086 12518 38088 12570
rect 38032 12516 38088 12518
rect 38136 12570 38192 12572
rect 38136 12518 38138 12570
rect 38138 12518 38190 12570
rect 38190 12518 38192 12570
rect 38136 12516 38192 12518
rect 38240 12570 38296 12572
rect 38240 12518 38242 12570
rect 38242 12518 38294 12570
rect 38294 12518 38296 12570
rect 38240 12516 38296 12518
rect 38032 11002 38088 11004
rect 38032 10950 38034 11002
rect 38034 10950 38086 11002
rect 38086 10950 38088 11002
rect 38032 10948 38088 10950
rect 38136 11002 38192 11004
rect 38136 10950 38138 11002
rect 38138 10950 38190 11002
rect 38190 10950 38192 11002
rect 38136 10948 38192 10950
rect 38240 11002 38296 11004
rect 38240 10950 38242 11002
rect 38242 10950 38294 11002
rect 38294 10950 38296 11002
rect 38240 10948 38296 10950
rect 38032 9434 38088 9436
rect 38032 9382 38034 9434
rect 38034 9382 38086 9434
rect 38086 9382 38088 9434
rect 38032 9380 38088 9382
rect 38136 9434 38192 9436
rect 38136 9382 38138 9434
rect 38138 9382 38190 9434
rect 38190 9382 38192 9434
rect 38136 9380 38192 9382
rect 38240 9434 38296 9436
rect 38240 9382 38242 9434
rect 38242 9382 38294 9434
rect 38294 9382 38296 9434
rect 38240 9380 38296 9382
rect 38032 7866 38088 7868
rect 38032 7814 38034 7866
rect 38034 7814 38086 7866
rect 38086 7814 38088 7866
rect 38032 7812 38088 7814
rect 38136 7866 38192 7868
rect 38136 7814 38138 7866
rect 38138 7814 38190 7866
rect 38190 7814 38192 7866
rect 38136 7812 38192 7814
rect 38240 7866 38296 7868
rect 38240 7814 38242 7866
rect 38242 7814 38294 7866
rect 38294 7814 38296 7866
rect 38240 7812 38296 7814
rect 38892 6524 38948 6580
rect 38032 6298 38088 6300
rect 38032 6246 38034 6298
rect 38034 6246 38086 6298
rect 38086 6246 38088 6298
rect 38032 6244 38088 6246
rect 38136 6298 38192 6300
rect 38136 6246 38138 6298
rect 38138 6246 38190 6298
rect 38190 6246 38192 6298
rect 38136 6244 38192 6246
rect 38240 6298 38296 6300
rect 38240 6246 38242 6298
rect 38242 6246 38294 6298
rect 38294 6246 38296 6298
rect 38240 6244 38296 6246
rect 39452 6524 39508 6580
rect 39452 5628 39508 5684
rect 38032 4730 38088 4732
rect 38032 4678 38034 4730
rect 38034 4678 38086 4730
rect 38086 4678 38088 4730
rect 38032 4676 38088 4678
rect 38136 4730 38192 4732
rect 38136 4678 38138 4730
rect 38138 4678 38190 4730
rect 38190 4678 38192 4730
rect 38136 4676 38192 4678
rect 38240 4730 38296 4732
rect 38240 4678 38242 4730
rect 38242 4678 38294 4730
rect 38294 4678 38296 4730
rect 38240 4676 38296 4678
rect 38032 3162 38088 3164
rect 38032 3110 38034 3162
rect 38034 3110 38086 3162
rect 38086 3110 38088 3162
rect 38032 3108 38088 3110
rect 38136 3162 38192 3164
rect 38136 3110 38138 3162
rect 38138 3110 38190 3162
rect 38190 3110 38192 3162
rect 38136 3108 38192 3110
rect 38240 3162 38296 3164
rect 38240 3110 38242 3162
rect 38242 3110 38294 3162
rect 38294 3110 38296 3162
rect 38240 3108 38296 3110
rect 43596 33964 43652 34020
rect 43036 32620 43092 32676
rect 43148 33068 43204 33124
rect 44492 33964 44548 34020
rect 44492 28812 44548 28868
rect 43596 27132 43652 27188
rect 44716 34130 44772 34132
rect 44716 34078 44718 34130
rect 44718 34078 44770 34130
rect 44770 34078 44772 34130
rect 44716 34076 44772 34078
rect 44716 33404 44772 33460
rect 44604 26124 44660 26180
rect 42924 19404 42980 19460
rect 39788 6130 39844 6132
rect 39788 6078 39790 6130
rect 39790 6078 39842 6130
rect 39842 6078 39844 6130
rect 39788 6076 39844 6078
rect 39788 5292 39844 5348
rect 41020 5122 41076 5124
rect 41020 5070 41022 5122
rect 41022 5070 41074 5122
rect 41074 5070 41076 5122
rect 41020 5068 41076 5070
rect 40236 4844 40292 4900
rect 40684 3500 40740 3556
rect 39564 3276 39620 3332
rect 41244 3554 41300 3556
rect 41244 3502 41246 3554
rect 41246 3502 41298 3554
rect 41298 3502 41300 3554
rect 41244 3500 41300 3502
rect 41020 3330 41076 3332
rect 41020 3278 41022 3330
rect 41022 3278 41074 3330
rect 41074 3278 41076 3330
rect 41020 3276 41076 3278
rect 44156 7308 44212 7364
rect 43372 6914 43428 6916
rect 43372 6862 43374 6914
rect 43374 6862 43426 6914
rect 43426 6862 43428 6914
rect 43372 6860 43428 6862
rect 43820 5906 43876 5908
rect 43820 5854 43822 5906
rect 43822 5854 43874 5906
rect 43874 5854 43876 5906
rect 43820 5852 43876 5854
rect 45612 35586 45668 35588
rect 45612 35534 45614 35586
rect 45614 35534 45666 35586
rect 45666 35534 45668 35586
rect 45612 35532 45668 35534
rect 45052 35084 45108 35140
rect 45724 35084 45780 35140
rect 47628 36876 47684 36932
rect 46732 36652 46788 36708
rect 47628 36652 47684 36708
rect 46060 35980 46116 36036
rect 46396 35810 46452 35812
rect 46396 35758 46398 35810
rect 46398 35758 46450 35810
rect 46450 35758 46452 35810
rect 46396 35756 46452 35758
rect 46172 35532 46228 35588
rect 46060 34242 46116 34244
rect 46060 34190 46062 34242
rect 46062 34190 46114 34242
rect 46114 34190 46116 34242
rect 46060 34188 46116 34190
rect 45276 34018 45332 34020
rect 45276 33966 45278 34018
rect 45278 33966 45330 34018
rect 45330 33966 45332 34018
rect 45276 33964 45332 33966
rect 45836 33404 45892 33460
rect 46956 35756 47012 35812
rect 46844 34636 46900 34692
rect 46284 33458 46340 33460
rect 46284 33406 46286 33458
rect 46286 33406 46338 33458
rect 46338 33406 46340 33458
rect 46284 33404 46340 33406
rect 47068 34300 47124 34356
rect 46956 33964 47012 34020
rect 45276 26908 45332 26964
rect 45164 7362 45220 7364
rect 45164 7310 45166 7362
rect 45166 7310 45218 7362
rect 45218 7310 45220 7362
rect 45164 7308 45220 7310
rect 44940 6860 44996 6916
rect 44604 6636 44660 6692
rect 44044 4844 44100 4900
rect 44156 5180 44212 5236
rect 44716 4844 44772 4900
rect 45052 4284 45108 4340
rect 43148 3164 43204 3220
rect 44156 3554 44212 3556
rect 44156 3502 44158 3554
rect 44158 3502 44210 3554
rect 44210 3502 44212 3554
rect 44156 3500 44212 3502
rect 45052 3500 45108 3556
rect 47516 36204 47572 36260
rect 48524 36540 48580 36596
rect 49308 37212 49364 37268
rect 47292 34300 47348 34356
rect 47740 34300 47796 34356
rect 47180 34076 47236 34132
rect 47404 34018 47460 34020
rect 47404 33966 47406 34018
rect 47406 33966 47458 34018
rect 47458 33966 47460 34018
rect 47404 33964 47460 33966
rect 48076 34690 48132 34692
rect 48076 34638 48078 34690
rect 48078 34638 48130 34690
rect 48130 34638 48132 34690
rect 48076 34636 48132 34638
rect 48524 34188 48580 34244
rect 48188 34130 48244 34132
rect 48188 34078 48190 34130
rect 48190 34078 48242 34130
rect 48242 34078 48244 34130
rect 48188 34076 48244 34078
rect 47068 26908 47124 26964
rect 48412 33964 48468 34020
rect 46060 17612 46116 17668
rect 46172 7308 46228 7364
rect 45948 6914 46004 6916
rect 45948 6862 45950 6914
rect 45950 6862 46002 6914
rect 46002 6862 46004 6914
rect 45948 6860 46004 6862
rect 45612 6690 45668 6692
rect 45612 6638 45614 6690
rect 45614 6638 45666 6690
rect 45666 6638 45668 6690
rect 45612 6636 45668 6638
rect 47180 7362 47236 7364
rect 47180 7310 47182 7362
rect 47182 7310 47234 7362
rect 47234 7310 47236 7362
rect 47180 7308 47236 7310
rect 48524 33180 48580 33236
rect 48412 24444 48468 24500
rect 49532 36594 49588 36596
rect 49532 36542 49534 36594
rect 49534 36542 49586 36594
rect 49586 36542 49588 36594
rect 49532 36540 49588 36542
rect 49196 35196 49252 35252
rect 48860 34354 48916 34356
rect 48860 34302 48862 34354
rect 48862 34302 48914 34354
rect 48914 34302 48916 34354
rect 48860 34300 48916 34302
rect 49532 35196 49588 35252
rect 51324 36594 51380 36596
rect 51324 36542 51326 36594
rect 51326 36542 51378 36594
rect 51378 36542 51380 36594
rect 51324 36540 51380 36542
rect 52892 37212 52948 37268
rect 52108 36540 52164 36596
rect 52668 36652 52724 36708
rect 51996 36092 52052 36148
rect 49980 35084 50036 35140
rect 49644 34300 49700 34356
rect 48636 11228 48692 11284
rect 47852 6860 47908 6916
rect 45948 5516 46004 5572
rect 45388 5122 45444 5124
rect 45388 5070 45390 5122
rect 45390 5070 45442 5122
rect 45442 5070 45444 5122
rect 45388 5068 45444 5070
rect 46508 5516 46564 5572
rect 47628 5906 47684 5908
rect 47628 5854 47630 5906
rect 47630 5854 47682 5906
rect 47682 5854 47684 5906
rect 47628 5852 47684 5854
rect 47740 5740 47796 5796
rect 47292 5516 47348 5572
rect 46396 5234 46452 5236
rect 46396 5182 46398 5234
rect 46398 5182 46450 5234
rect 46450 5182 46452 5234
rect 46396 5180 46452 5182
rect 46620 5180 46676 5236
rect 47180 5234 47236 5236
rect 47180 5182 47182 5234
rect 47182 5182 47234 5234
rect 47234 5182 47236 5234
rect 47180 5180 47236 5182
rect 48188 4562 48244 4564
rect 48188 4510 48190 4562
rect 48190 4510 48242 4562
rect 48242 4510 48244 4562
rect 48188 4508 48244 4510
rect 45948 4172 46004 4228
rect 46172 4172 46228 4228
rect 47180 4226 47236 4228
rect 47180 4174 47182 4226
rect 47182 4174 47234 4226
rect 47234 4174 47236 4226
rect 47180 4172 47236 4174
rect 45948 3330 46004 3332
rect 45948 3278 45950 3330
rect 45950 3278 46002 3330
rect 46002 3278 46004 3330
rect 45948 3276 46004 3278
rect 50316 34636 50372 34692
rect 49868 28028 49924 28084
rect 50988 34300 51044 34356
rect 51212 34018 51268 34020
rect 51212 33966 51214 34018
rect 51214 33966 51266 34018
rect 51266 33966 51268 34018
rect 51212 33964 51268 33966
rect 50316 26236 50372 26292
rect 50652 33516 50708 33572
rect 49532 26012 49588 26068
rect 50540 6466 50596 6468
rect 50540 6414 50542 6466
rect 50542 6414 50594 6466
rect 50594 6414 50596 6466
rect 50540 6412 50596 6414
rect 50540 5628 50596 5684
rect 49532 3276 49588 3332
rect 51212 33516 51268 33572
rect 53900 36652 53956 36708
rect 53788 35868 53844 35924
rect 53004 35474 53060 35476
rect 53004 35422 53006 35474
rect 53006 35422 53058 35474
rect 53058 35422 53060 35474
rect 53004 35420 53060 35422
rect 51548 33346 51604 33348
rect 51548 33294 51550 33346
rect 51550 33294 51602 33346
rect 51602 33294 51604 33346
rect 51548 33292 51604 33294
rect 51660 35308 51716 35364
rect 51660 34188 51716 34244
rect 52220 34412 52276 34468
rect 52332 33964 52388 34020
rect 52444 33292 52500 33348
rect 53116 34242 53172 34244
rect 53116 34190 53118 34242
rect 53118 34190 53170 34242
rect 53170 34190 53172 34242
rect 53116 34188 53172 34190
rect 53452 34242 53508 34244
rect 53452 34190 53454 34242
rect 53454 34190 53506 34242
rect 53506 34190 53508 34242
rect 53452 34188 53508 34190
rect 53340 33458 53396 33460
rect 53340 33406 53342 33458
rect 53342 33406 53394 33458
rect 53394 33406 53396 33458
rect 53340 33404 53396 33406
rect 52780 33346 52836 33348
rect 52780 33294 52782 33346
rect 52782 33294 52834 33346
rect 52834 33294 52836 33346
rect 52780 33292 52836 33294
rect 51996 30156 52052 30212
rect 53788 35532 53844 35588
rect 53676 35420 53732 35476
rect 53340 31052 53396 31108
rect 52444 29596 52500 29652
rect 51660 26012 51716 26068
rect 53004 14252 53060 14308
rect 51660 7308 51716 7364
rect 50988 6466 51044 6468
rect 50988 6414 50990 6466
rect 50990 6414 51042 6466
rect 51042 6414 51044 6466
rect 50988 6412 51044 6414
rect 51324 6300 51380 6356
rect 51436 4172 51492 4228
rect 51212 3442 51268 3444
rect 51212 3390 51214 3442
rect 51214 3390 51266 3442
rect 51266 3390 51268 3442
rect 51212 3388 51268 3390
rect 52556 7196 52612 7252
rect 52668 6300 52724 6356
rect 52892 5964 52948 6020
rect 51884 4226 51940 4228
rect 51884 4174 51886 4226
rect 51886 4174 51938 4226
rect 51938 4174 51940 4226
rect 51884 4172 51940 4174
rect 51996 3554 52052 3556
rect 51996 3502 51998 3554
rect 51998 3502 52050 3554
rect 52050 3502 52052 3554
rect 51996 3500 52052 3502
rect 52332 3500 52388 3556
rect 52780 3500 52836 3556
rect 53452 7196 53508 7252
rect 53116 6018 53172 6020
rect 53116 5966 53118 6018
rect 53118 5966 53170 6018
rect 53170 5966 53172 6018
rect 53116 5964 53172 5966
rect 54236 35532 54292 35588
rect 54012 34524 54068 34580
rect 54012 33404 54068 33460
rect 54572 36092 54628 36148
rect 54796 35868 54852 35924
rect 54908 35698 54964 35700
rect 54908 35646 54910 35698
rect 54910 35646 54962 35698
rect 54962 35646 54964 35698
rect 54908 35644 54964 35646
rect 54572 34914 54628 34916
rect 54572 34862 54574 34914
rect 54574 34862 54626 34914
rect 54626 34862 54628 34914
rect 54572 34860 54628 34862
rect 56924 38220 56980 38276
rect 55020 34914 55076 34916
rect 55020 34862 55022 34914
rect 55022 34862 55074 34914
rect 55074 34862 55076 34914
rect 55020 34860 55076 34862
rect 55244 35644 55300 35700
rect 54460 33346 54516 33348
rect 54460 33294 54462 33346
rect 54462 33294 54514 33346
rect 54514 33294 54516 33346
rect 54460 33292 54516 33294
rect 54348 31052 54404 31108
rect 54572 7196 54628 7252
rect 54012 6300 54068 6356
rect 53676 5234 53732 5236
rect 53676 5182 53678 5234
rect 53678 5182 53730 5234
rect 53730 5182 53732 5234
rect 53676 5180 53732 5182
rect 54460 5180 54516 5236
rect 53452 4338 53508 4340
rect 53452 4286 53454 4338
rect 53454 4286 53506 4338
rect 53506 4286 53508 4338
rect 53452 4284 53508 4286
rect 54012 4284 54068 4340
rect 56442 36874 56498 36876
rect 56442 36822 56444 36874
rect 56444 36822 56496 36874
rect 56496 36822 56498 36874
rect 56442 36820 56498 36822
rect 56546 36874 56602 36876
rect 56546 36822 56548 36874
rect 56548 36822 56600 36874
rect 56600 36822 56602 36874
rect 56546 36820 56602 36822
rect 56650 36874 56706 36876
rect 56650 36822 56652 36874
rect 56652 36822 56704 36874
rect 56704 36822 56706 36874
rect 56650 36820 56706 36822
rect 56700 35698 56756 35700
rect 56700 35646 56702 35698
rect 56702 35646 56754 35698
rect 56754 35646 56756 35698
rect 56700 35644 56756 35646
rect 56442 35306 56498 35308
rect 56442 35254 56444 35306
rect 56444 35254 56496 35306
rect 56496 35254 56498 35306
rect 56442 35252 56498 35254
rect 56546 35306 56602 35308
rect 56546 35254 56548 35306
rect 56548 35254 56600 35306
rect 56600 35254 56602 35306
rect 56546 35252 56602 35254
rect 56650 35306 56706 35308
rect 56650 35254 56652 35306
rect 56652 35254 56704 35306
rect 56704 35254 56706 35306
rect 56650 35252 56706 35254
rect 56028 34860 56084 34916
rect 56476 34802 56532 34804
rect 56476 34750 56478 34802
rect 56478 34750 56530 34802
rect 56530 34750 56532 34802
rect 56476 34748 56532 34750
rect 56028 34188 56084 34244
rect 55804 33516 55860 33572
rect 56140 34018 56196 34020
rect 56140 33966 56142 34018
rect 56142 33966 56194 34018
rect 56194 33966 56196 34018
rect 56140 33964 56196 33966
rect 56476 33964 56532 34020
rect 57148 37996 57204 38052
rect 57596 36428 57652 36484
rect 57484 35644 57540 35700
rect 57372 34914 57428 34916
rect 57372 34862 57374 34914
rect 57374 34862 57426 34914
rect 57426 34862 57428 34914
rect 57372 34860 57428 34862
rect 56588 33852 56644 33908
rect 56442 33738 56498 33740
rect 56028 31164 56084 31220
rect 56252 33628 56308 33684
rect 56442 33686 56444 33738
rect 56444 33686 56496 33738
rect 56496 33686 56498 33738
rect 56442 33684 56498 33686
rect 56546 33738 56602 33740
rect 56546 33686 56548 33738
rect 56548 33686 56600 33738
rect 56600 33686 56602 33738
rect 56546 33684 56602 33686
rect 56650 33738 56706 33740
rect 56650 33686 56652 33738
rect 56652 33686 56704 33738
rect 56704 33686 56706 33738
rect 56650 33684 56706 33686
rect 55356 29932 55412 29988
rect 55244 19292 55300 19348
rect 56442 32170 56498 32172
rect 56442 32118 56444 32170
rect 56444 32118 56496 32170
rect 56496 32118 56498 32170
rect 56442 32116 56498 32118
rect 56546 32170 56602 32172
rect 56546 32118 56548 32170
rect 56548 32118 56600 32170
rect 56600 32118 56602 32170
rect 56546 32116 56602 32118
rect 56650 32170 56706 32172
rect 56650 32118 56652 32170
rect 56652 32118 56704 32170
rect 56704 32118 56706 32170
rect 56650 32116 56706 32118
rect 56442 30602 56498 30604
rect 56442 30550 56444 30602
rect 56444 30550 56496 30602
rect 56496 30550 56498 30602
rect 56442 30548 56498 30550
rect 56546 30602 56602 30604
rect 56546 30550 56548 30602
rect 56548 30550 56600 30602
rect 56600 30550 56602 30602
rect 56546 30548 56602 30550
rect 56650 30602 56706 30604
rect 56650 30550 56652 30602
rect 56652 30550 56704 30602
rect 56704 30550 56706 30602
rect 56650 30548 56706 30550
rect 57708 31500 57764 31556
rect 58940 38556 58996 38612
rect 58828 36482 58884 36484
rect 58828 36430 58830 36482
rect 58830 36430 58882 36482
rect 58882 36430 58884 36482
rect 58828 36428 58884 36430
rect 58716 36204 58772 36260
rect 58604 35810 58660 35812
rect 58604 35758 58606 35810
rect 58606 35758 58658 35810
rect 58658 35758 58660 35810
rect 58604 35756 58660 35758
rect 57484 29484 57540 29540
rect 56442 29034 56498 29036
rect 56442 28982 56444 29034
rect 56444 28982 56496 29034
rect 56496 28982 56498 29034
rect 56442 28980 56498 28982
rect 56546 29034 56602 29036
rect 56546 28982 56548 29034
rect 56548 28982 56600 29034
rect 56600 28982 56602 29034
rect 56546 28980 56602 28982
rect 56650 29034 56706 29036
rect 56650 28982 56652 29034
rect 56652 28982 56704 29034
rect 56704 28982 56706 29034
rect 56650 28980 56706 28982
rect 56442 27466 56498 27468
rect 56442 27414 56444 27466
rect 56444 27414 56496 27466
rect 56496 27414 56498 27466
rect 56442 27412 56498 27414
rect 56546 27466 56602 27468
rect 56546 27414 56548 27466
rect 56548 27414 56600 27466
rect 56600 27414 56602 27466
rect 56546 27412 56602 27414
rect 56650 27466 56706 27468
rect 56650 27414 56652 27466
rect 56652 27414 56704 27466
rect 56704 27414 56706 27466
rect 56650 27412 56706 27414
rect 56442 25898 56498 25900
rect 56442 25846 56444 25898
rect 56444 25846 56496 25898
rect 56496 25846 56498 25898
rect 56442 25844 56498 25846
rect 56546 25898 56602 25900
rect 56546 25846 56548 25898
rect 56548 25846 56600 25898
rect 56600 25846 56602 25898
rect 56546 25844 56602 25846
rect 56650 25898 56706 25900
rect 56650 25846 56652 25898
rect 56652 25846 56704 25898
rect 56704 25846 56706 25898
rect 56650 25844 56706 25846
rect 56442 24330 56498 24332
rect 56442 24278 56444 24330
rect 56444 24278 56496 24330
rect 56496 24278 56498 24330
rect 56442 24276 56498 24278
rect 56546 24330 56602 24332
rect 56546 24278 56548 24330
rect 56548 24278 56600 24330
rect 56600 24278 56602 24330
rect 56546 24276 56602 24278
rect 56650 24330 56706 24332
rect 56650 24278 56652 24330
rect 56652 24278 56704 24330
rect 56704 24278 56706 24330
rect 56650 24276 56706 24278
rect 56442 22762 56498 22764
rect 56442 22710 56444 22762
rect 56444 22710 56496 22762
rect 56496 22710 56498 22762
rect 56442 22708 56498 22710
rect 56546 22762 56602 22764
rect 56546 22710 56548 22762
rect 56548 22710 56600 22762
rect 56600 22710 56602 22762
rect 56546 22708 56602 22710
rect 56650 22762 56706 22764
rect 56650 22710 56652 22762
rect 56652 22710 56704 22762
rect 56704 22710 56706 22762
rect 56650 22708 56706 22710
rect 56442 21194 56498 21196
rect 56442 21142 56444 21194
rect 56444 21142 56496 21194
rect 56496 21142 56498 21194
rect 56442 21140 56498 21142
rect 56546 21194 56602 21196
rect 56546 21142 56548 21194
rect 56548 21142 56600 21194
rect 56600 21142 56602 21194
rect 56546 21140 56602 21142
rect 56650 21194 56706 21196
rect 56650 21142 56652 21194
rect 56652 21142 56704 21194
rect 56704 21142 56706 21194
rect 56650 21140 56706 21142
rect 56442 19626 56498 19628
rect 56442 19574 56444 19626
rect 56444 19574 56496 19626
rect 56496 19574 56498 19626
rect 56442 19572 56498 19574
rect 56546 19626 56602 19628
rect 56546 19574 56548 19626
rect 56548 19574 56600 19626
rect 56600 19574 56602 19626
rect 56546 19572 56602 19574
rect 56650 19626 56706 19628
rect 56650 19574 56652 19626
rect 56652 19574 56704 19626
rect 56704 19574 56706 19626
rect 56650 19572 56706 19574
rect 56442 18058 56498 18060
rect 56442 18006 56444 18058
rect 56444 18006 56496 18058
rect 56496 18006 56498 18058
rect 56442 18004 56498 18006
rect 56546 18058 56602 18060
rect 56546 18006 56548 18058
rect 56548 18006 56600 18058
rect 56600 18006 56602 18058
rect 56546 18004 56602 18006
rect 56650 18058 56706 18060
rect 56650 18006 56652 18058
rect 56652 18006 56704 18058
rect 56704 18006 56706 18058
rect 56650 18004 56706 18006
rect 56442 16490 56498 16492
rect 56442 16438 56444 16490
rect 56444 16438 56496 16490
rect 56496 16438 56498 16490
rect 56442 16436 56498 16438
rect 56546 16490 56602 16492
rect 56546 16438 56548 16490
rect 56548 16438 56600 16490
rect 56600 16438 56602 16490
rect 56546 16436 56602 16438
rect 56650 16490 56706 16492
rect 56650 16438 56652 16490
rect 56652 16438 56704 16490
rect 56704 16438 56706 16490
rect 56650 16436 56706 16438
rect 56442 14922 56498 14924
rect 56442 14870 56444 14922
rect 56444 14870 56496 14922
rect 56496 14870 56498 14922
rect 56442 14868 56498 14870
rect 56546 14922 56602 14924
rect 56546 14870 56548 14922
rect 56548 14870 56600 14922
rect 56600 14870 56602 14922
rect 56546 14868 56602 14870
rect 56650 14922 56706 14924
rect 56650 14870 56652 14922
rect 56652 14870 56704 14922
rect 56704 14870 56706 14922
rect 56650 14868 56706 14870
rect 56442 13354 56498 13356
rect 56442 13302 56444 13354
rect 56444 13302 56496 13354
rect 56496 13302 56498 13354
rect 56442 13300 56498 13302
rect 56546 13354 56602 13356
rect 56546 13302 56548 13354
rect 56548 13302 56600 13354
rect 56600 13302 56602 13354
rect 56546 13300 56602 13302
rect 56650 13354 56706 13356
rect 56650 13302 56652 13354
rect 56652 13302 56704 13354
rect 56704 13302 56706 13354
rect 56650 13300 56706 13302
rect 59612 37324 59668 37380
rect 59164 36428 59220 36484
rect 58716 32732 58772 32788
rect 58156 30156 58212 30212
rect 58940 30044 58996 30100
rect 59052 33964 59108 34020
rect 57820 12684 57876 12740
rect 56442 11786 56498 11788
rect 56442 11734 56444 11786
rect 56444 11734 56496 11786
rect 56496 11734 56498 11786
rect 56442 11732 56498 11734
rect 56546 11786 56602 11788
rect 56546 11734 56548 11786
rect 56548 11734 56600 11786
rect 56600 11734 56602 11786
rect 56546 11732 56602 11734
rect 56650 11786 56706 11788
rect 56650 11734 56652 11786
rect 56652 11734 56704 11786
rect 56704 11734 56706 11786
rect 56650 11732 56706 11734
rect 56442 10218 56498 10220
rect 56442 10166 56444 10218
rect 56444 10166 56496 10218
rect 56496 10166 56498 10218
rect 56442 10164 56498 10166
rect 56546 10218 56602 10220
rect 56546 10166 56548 10218
rect 56548 10166 56600 10218
rect 56600 10166 56602 10218
rect 56546 10164 56602 10166
rect 56650 10218 56706 10220
rect 56650 10166 56652 10218
rect 56652 10166 56704 10218
rect 56704 10166 56706 10218
rect 56650 10164 56706 10166
rect 56442 8650 56498 8652
rect 56442 8598 56444 8650
rect 56444 8598 56496 8650
rect 56496 8598 56498 8650
rect 56442 8596 56498 8598
rect 56546 8650 56602 8652
rect 56546 8598 56548 8650
rect 56548 8598 56600 8650
rect 56600 8598 56602 8650
rect 56546 8596 56602 8598
rect 56650 8650 56706 8652
rect 56650 8598 56652 8650
rect 56652 8598 56704 8650
rect 56704 8598 56706 8650
rect 56650 8596 56706 8598
rect 58156 8092 58212 8148
rect 56252 7308 56308 7364
rect 57708 7532 57764 7588
rect 56442 7082 56498 7084
rect 56442 7030 56444 7082
rect 56444 7030 56496 7082
rect 56496 7030 56498 7082
rect 56442 7028 56498 7030
rect 56546 7082 56602 7084
rect 56546 7030 56548 7082
rect 56548 7030 56600 7082
rect 56600 7030 56602 7082
rect 56546 7028 56602 7030
rect 56650 7082 56706 7084
rect 56650 7030 56652 7082
rect 56652 7030 56704 7082
rect 56704 7030 56706 7082
rect 56650 7028 56706 7030
rect 54684 5180 54740 5236
rect 54012 3612 54068 3668
rect 53788 3500 53844 3556
rect 53340 3442 53396 3444
rect 53340 3390 53342 3442
rect 53342 3390 53394 3442
rect 53394 3390 53396 3442
rect 53340 3388 53396 3390
rect 54124 3388 54180 3444
rect 53788 2940 53844 2996
rect 55244 6076 55300 6132
rect 55692 6076 55748 6132
rect 55356 5852 55412 5908
rect 57148 5852 57204 5908
rect 57820 5906 57876 5908
rect 57820 5854 57822 5906
rect 57822 5854 57874 5906
rect 57874 5854 57876 5906
rect 57820 5852 57876 5854
rect 55692 5628 55748 5684
rect 56442 5514 56498 5516
rect 56442 5462 56444 5514
rect 56444 5462 56496 5514
rect 56496 5462 56498 5514
rect 56442 5460 56498 5462
rect 56546 5514 56602 5516
rect 56546 5462 56548 5514
rect 56548 5462 56600 5514
rect 56600 5462 56602 5514
rect 56546 5460 56602 5462
rect 56650 5514 56706 5516
rect 56650 5462 56652 5514
rect 56652 5462 56704 5514
rect 56704 5462 56706 5514
rect 56650 5460 56706 5462
rect 55692 5180 55748 5236
rect 55244 4508 55300 4564
rect 56812 4508 56868 4564
rect 55132 3778 55188 3780
rect 55132 3726 55134 3778
rect 55134 3726 55186 3778
rect 55186 3726 55188 3778
rect 55132 3724 55188 3726
rect 56364 4060 56420 4116
rect 57484 4956 57540 5012
rect 57932 5404 57988 5460
rect 56442 3946 56498 3948
rect 56442 3894 56444 3946
rect 56444 3894 56496 3946
rect 56496 3894 56498 3946
rect 56442 3892 56498 3894
rect 56546 3946 56602 3948
rect 56546 3894 56548 3946
rect 56548 3894 56600 3946
rect 56600 3894 56602 3946
rect 56546 3892 56602 3894
rect 56650 3946 56706 3948
rect 56650 3894 56652 3946
rect 56652 3894 56704 3946
rect 56704 3894 56706 3946
rect 56650 3892 56706 3894
rect 55916 3554 55972 3556
rect 55916 3502 55918 3554
rect 55918 3502 55970 3554
rect 55970 3502 55972 3554
rect 55916 3500 55972 3502
rect 55468 3388 55524 3444
rect 57596 3724 57652 3780
rect 58268 5794 58324 5796
rect 58268 5742 58270 5794
rect 58270 5742 58322 5794
rect 58322 5742 58324 5794
rect 58268 5740 58324 5742
rect 58268 5180 58324 5236
rect 58156 4956 58212 5012
rect 57036 3442 57092 3444
rect 57036 3390 57038 3442
rect 57038 3390 57090 3442
rect 57090 3390 57092 3442
rect 57036 3388 57092 3390
rect 56924 2940 56980 2996
rect 59500 36204 59556 36260
rect 59276 35756 59332 35812
rect 59612 34860 59668 34916
rect 59836 34018 59892 34020
rect 59836 33966 59838 34018
rect 59838 33966 59890 34018
rect 59890 33966 59892 34018
rect 59836 33964 59892 33966
rect 60172 35756 60228 35812
rect 60732 37660 60788 37716
rect 61404 37884 61460 37940
rect 61292 36764 61348 36820
rect 60060 34076 60116 34132
rect 60620 34076 60676 34132
rect 60172 34018 60228 34020
rect 60172 33966 60174 34018
rect 60174 33966 60226 34018
rect 60226 33966 60228 34018
rect 60172 33964 60228 33966
rect 60284 33458 60340 33460
rect 60284 33406 60286 33458
rect 60286 33406 60338 33458
rect 60338 33406 60340 33458
rect 60284 33404 60340 33406
rect 61404 36428 61460 36484
rect 61292 35532 61348 35588
rect 61180 34130 61236 34132
rect 61180 34078 61182 34130
rect 61182 34078 61234 34130
rect 61234 34078 61236 34130
rect 61180 34076 61236 34078
rect 60732 33404 60788 33460
rect 61292 33292 61348 33348
rect 61404 33628 61460 33684
rect 59948 27804 60004 27860
rect 60284 32396 60340 32452
rect 60284 26796 60340 26852
rect 59052 14252 59108 14308
rect 60284 14252 60340 14308
rect 59052 11564 59108 11620
rect 58492 4508 58548 4564
rect 60284 11564 60340 11620
rect 59612 9212 59668 9268
rect 59164 7586 59220 7588
rect 59164 7534 59166 7586
rect 59166 7534 59218 7586
rect 59218 7534 59220 7586
rect 59164 7532 59220 7534
rect 59500 7474 59556 7476
rect 59500 7422 59502 7474
rect 59502 7422 59554 7474
rect 59554 7422 59556 7474
rect 59500 7420 59556 7422
rect 58828 5516 58884 5572
rect 59052 4844 59108 4900
rect 59388 5794 59444 5796
rect 59388 5742 59390 5794
rect 59390 5742 59442 5794
rect 59442 5742 59444 5794
rect 59388 5740 59444 5742
rect 59276 5180 59332 5236
rect 59276 5010 59332 5012
rect 59276 4958 59278 5010
rect 59278 4958 59330 5010
rect 59330 4958 59332 5010
rect 59276 4956 59332 4958
rect 61740 33458 61796 33460
rect 61740 33406 61742 33458
rect 61742 33406 61794 33458
rect 61794 33406 61796 33458
rect 61740 33404 61796 33406
rect 61628 32732 61684 32788
rect 62636 37324 62692 37380
rect 62524 36988 62580 37044
rect 62188 34914 62244 34916
rect 62188 34862 62190 34914
rect 62190 34862 62242 34914
rect 62242 34862 62244 34914
rect 62188 34860 62244 34862
rect 62300 34130 62356 34132
rect 62300 34078 62302 34130
rect 62302 34078 62354 34130
rect 62354 34078 62356 34130
rect 62300 34076 62356 34078
rect 61964 33404 62020 33460
rect 61852 32396 61908 32452
rect 62076 33068 62132 33124
rect 62636 34354 62692 34356
rect 62636 34302 62638 34354
rect 62638 34302 62690 34354
rect 62690 34302 62692 34354
rect 62636 34300 62692 34302
rect 62860 34972 62916 35028
rect 63084 34300 63140 34356
rect 62748 33292 62804 33348
rect 62412 33068 62468 33124
rect 62636 31948 62692 32004
rect 62972 32786 63028 32788
rect 62972 32734 62974 32786
rect 62974 32734 63026 32786
rect 63026 32734 63028 32786
rect 62972 32732 63028 32734
rect 62076 31836 62132 31892
rect 63420 35026 63476 35028
rect 63420 34974 63422 35026
rect 63422 34974 63474 35026
rect 63474 34974 63476 35026
rect 63420 34972 63476 34974
rect 63532 33628 63588 33684
rect 63420 33404 63476 33460
rect 63308 33292 63364 33348
rect 63196 32732 63252 32788
rect 62972 27916 63028 27972
rect 59948 6578 60004 6580
rect 59948 6526 59950 6578
rect 59950 6526 60002 6578
rect 60002 6526 60004 6578
rect 59948 6524 60004 6526
rect 59836 5906 59892 5908
rect 59836 5854 59838 5906
rect 59838 5854 59890 5906
rect 59890 5854 59892 5906
rect 59836 5852 59892 5854
rect 62188 8428 62244 8484
rect 60956 7474 61012 7476
rect 60956 7422 60958 7474
rect 60958 7422 61010 7474
rect 61010 7422 61012 7474
rect 60956 7420 61012 7422
rect 61628 7196 61684 7252
rect 60284 6412 60340 6468
rect 60732 5964 60788 6020
rect 61292 6466 61348 6468
rect 61292 6414 61294 6466
rect 61294 6414 61346 6466
rect 61346 6414 61348 6466
rect 61292 6412 61348 6414
rect 60284 5852 60340 5908
rect 60508 5404 60564 5460
rect 60620 5010 60676 5012
rect 60620 4958 60622 5010
rect 60622 4958 60674 5010
rect 60674 4958 60676 5010
rect 60620 4956 60676 4958
rect 59612 4732 59668 4788
rect 58940 3612 58996 3668
rect 60844 3612 60900 3668
rect 59836 3554 59892 3556
rect 59836 3502 59838 3554
rect 59838 3502 59890 3554
rect 59890 3502 59892 3554
rect 59836 3500 59892 3502
rect 59612 3388 59668 3444
rect 58604 3164 58660 3220
rect 59500 2940 59556 2996
rect 58604 2716 58660 2772
rect 58380 2604 58436 2660
rect 62076 7474 62132 7476
rect 62076 7422 62078 7474
rect 62078 7422 62130 7474
rect 62130 7422 62132 7474
rect 62076 7420 62132 7422
rect 61852 6578 61908 6580
rect 61852 6526 61854 6578
rect 61854 6526 61906 6578
rect 61906 6526 61908 6578
rect 61852 6524 61908 6526
rect 62412 6412 62468 6468
rect 62860 7586 62916 7588
rect 62860 7534 62862 7586
rect 62862 7534 62914 7586
rect 62914 7534 62916 7586
rect 62860 7532 62916 7534
rect 63084 6076 63140 6132
rect 61740 5964 61796 6020
rect 64316 37436 64372 37492
rect 63868 34748 63924 34804
rect 63868 34354 63924 34356
rect 63868 34302 63870 34354
rect 63870 34302 63922 34354
rect 63922 34302 63924 34354
rect 63868 34300 63924 34302
rect 64652 37212 64708 37268
rect 64540 36594 64596 36596
rect 64540 36542 64542 36594
rect 64542 36542 64594 36594
rect 64594 36542 64596 36594
rect 64540 36540 64596 36542
rect 64988 36482 65044 36484
rect 64988 36430 64990 36482
rect 64990 36430 65042 36482
rect 65042 36430 65044 36482
rect 64988 36428 65044 36430
rect 65548 36428 65604 36484
rect 65324 36370 65380 36372
rect 65324 36318 65326 36370
rect 65326 36318 65378 36370
rect 65378 36318 65380 36370
rect 65324 36316 65380 36318
rect 65436 34412 65492 34468
rect 64764 34188 64820 34244
rect 63756 33346 63812 33348
rect 63756 33294 63758 33346
rect 63758 33294 63810 33346
rect 63810 33294 63812 33346
rect 63756 33292 63812 33294
rect 64204 32732 64260 32788
rect 65100 33458 65156 33460
rect 65100 33406 65102 33458
rect 65102 33406 65154 33458
rect 65154 33406 65156 33458
rect 65100 33404 65156 33406
rect 65660 38108 65716 38164
rect 66108 36540 66164 36596
rect 66444 36540 66500 36596
rect 65660 36316 65716 36372
rect 65772 34412 65828 34468
rect 66780 36482 66836 36484
rect 66780 36430 66782 36482
rect 66782 36430 66834 36482
rect 66834 36430 66836 36482
rect 66780 36428 66836 36430
rect 66108 35698 66164 35700
rect 66108 35646 66110 35698
rect 66110 35646 66162 35698
rect 66162 35646 66164 35698
rect 66108 35644 66164 35646
rect 66668 35644 66724 35700
rect 66556 35474 66612 35476
rect 66556 35422 66558 35474
rect 66558 35422 66610 35474
rect 66610 35422 66612 35474
rect 66556 35420 66612 35422
rect 66668 35026 66724 35028
rect 66668 34974 66670 35026
rect 66670 34974 66722 35026
rect 66722 34974 66724 35026
rect 66668 34972 66724 34974
rect 65884 32844 65940 32900
rect 66332 34076 66388 34132
rect 64764 30828 64820 30884
rect 66444 31612 66500 31668
rect 64540 8428 64596 8484
rect 63644 8204 63700 8260
rect 63420 7474 63476 7476
rect 63420 7422 63422 7474
rect 63422 7422 63474 7474
rect 63474 7422 63476 7474
rect 63420 7420 63476 7422
rect 63532 7196 63588 7252
rect 63308 5740 63364 5796
rect 62860 5122 62916 5124
rect 62860 5070 62862 5122
rect 62862 5070 62914 5122
rect 62914 5070 62916 5122
rect 62860 5068 62916 5070
rect 62188 4956 62244 5012
rect 60956 3442 61012 3444
rect 60956 3390 60958 3442
rect 60958 3390 61010 3442
rect 61010 3390 61012 3442
rect 60956 3388 61012 3390
rect 62412 3554 62468 3556
rect 62412 3502 62414 3554
rect 62414 3502 62466 3554
rect 62466 3502 62468 3554
rect 62412 3500 62468 3502
rect 62748 3500 62804 3556
rect 63532 3724 63588 3780
rect 64540 8258 64596 8260
rect 64540 8206 64542 8258
rect 64542 8206 64594 8258
rect 64594 8206 64596 8258
rect 64540 8204 64596 8206
rect 63980 8146 64036 8148
rect 63980 8094 63982 8146
rect 63982 8094 64034 8146
rect 64034 8094 64036 8146
rect 63980 8092 64036 8094
rect 63868 7420 63924 7476
rect 64204 7532 64260 7588
rect 63980 6130 64036 6132
rect 63980 6078 63982 6130
rect 63982 6078 64034 6130
rect 64034 6078 64036 6130
rect 63980 6076 64036 6078
rect 64652 6636 64708 6692
rect 65772 8316 65828 8372
rect 65436 8092 65492 8148
rect 65996 7980 66052 8036
rect 65548 7474 65604 7476
rect 65548 7422 65550 7474
rect 65550 7422 65602 7474
rect 65602 7422 65604 7474
rect 65548 7420 65604 7422
rect 63980 5234 64036 5236
rect 63980 5182 63982 5234
rect 63982 5182 64034 5234
rect 64034 5182 64036 5234
rect 63980 5180 64036 5182
rect 63868 5068 63924 5124
rect 66556 8146 66612 8148
rect 66556 8094 66558 8146
rect 66558 8094 66610 8146
rect 66610 8094 66612 8146
rect 66556 8092 66612 8094
rect 66444 7644 66500 7700
rect 67116 34914 67172 34916
rect 67116 34862 67118 34914
rect 67118 34862 67170 34914
rect 67170 34862 67172 34914
rect 67116 34860 67172 34862
rect 68236 36876 68292 36932
rect 68796 37772 68852 37828
rect 67900 36540 67956 36596
rect 67676 36428 67732 36484
rect 67340 34860 67396 34916
rect 67452 35420 67508 35476
rect 67004 34076 67060 34132
rect 67564 34914 67620 34916
rect 67564 34862 67566 34914
rect 67566 34862 67618 34914
rect 67618 34862 67620 34914
rect 67564 34860 67620 34862
rect 67788 36370 67844 36372
rect 67788 36318 67790 36370
rect 67790 36318 67842 36370
rect 67842 36318 67844 36370
rect 67788 36316 67844 36318
rect 68796 36540 68852 36596
rect 68908 36876 68964 36932
rect 68572 36092 68628 36148
rect 67452 32508 67508 32564
rect 68684 35026 68740 35028
rect 68684 34974 68686 35026
rect 68686 34974 68738 35026
rect 68738 34974 68740 35026
rect 68684 34972 68740 34974
rect 68572 33740 68628 33796
rect 69692 37772 69748 37828
rect 70028 36876 70084 36932
rect 70588 36876 70644 36932
rect 69692 36316 69748 36372
rect 70812 36092 70868 36148
rect 70476 35810 70532 35812
rect 70476 35758 70478 35810
rect 70478 35758 70530 35810
rect 70530 35758 70532 35810
rect 70476 35756 70532 35758
rect 70924 35756 70980 35812
rect 69916 35644 69972 35700
rect 69580 35196 69636 35252
rect 70140 35196 70196 35252
rect 69132 34972 69188 35028
rect 72492 37100 72548 37156
rect 71596 35196 71652 35252
rect 72044 35026 72100 35028
rect 72044 34974 72046 35026
rect 72046 34974 72098 35026
rect 72098 34974 72100 35026
rect 72044 34972 72100 34974
rect 68012 30156 68068 30212
rect 72156 33964 72212 34020
rect 72604 36204 72660 36260
rect 72828 38668 72884 38724
rect 73836 37100 73892 37156
rect 72828 36092 72884 36148
rect 73724 36092 73780 36148
rect 72716 34972 72772 35028
rect 73276 35308 73332 35364
rect 74396 36764 74452 36820
rect 75068 36876 75124 36932
rect 74508 36092 74564 36148
rect 74284 35532 74340 35588
rect 73164 34524 73220 34580
rect 73836 34524 73892 34580
rect 73948 34354 74004 34356
rect 73948 34302 73950 34354
rect 73950 34302 74002 34354
rect 74002 34302 74004 34354
rect 73948 34300 74004 34302
rect 74172 34188 74228 34244
rect 72716 33404 72772 33460
rect 74396 34748 74452 34804
rect 74620 36764 74676 36820
rect 74852 36090 74908 36092
rect 74852 36038 74854 36090
rect 74854 36038 74906 36090
rect 74906 36038 74908 36090
rect 74852 36036 74908 36038
rect 74956 36090 75012 36092
rect 74956 36038 74958 36090
rect 74958 36038 75010 36090
rect 75010 36038 75012 36090
rect 74956 36036 75012 36038
rect 75060 36090 75116 36092
rect 75060 36038 75062 36090
rect 75062 36038 75114 36090
rect 75114 36038 75116 36090
rect 75060 36036 75116 36038
rect 74620 35532 74676 35588
rect 74732 35308 74788 35364
rect 74732 34914 74788 34916
rect 74732 34862 74734 34914
rect 74734 34862 74786 34914
rect 74786 34862 74788 34914
rect 74732 34860 74788 34862
rect 74732 34636 74788 34692
rect 75404 35474 75460 35476
rect 75404 35422 75406 35474
rect 75406 35422 75458 35474
rect 75458 35422 75460 35474
rect 75404 35420 75460 35422
rect 75292 34860 75348 34916
rect 75404 34748 75460 34804
rect 74852 34522 74908 34524
rect 74852 34470 74854 34522
rect 74854 34470 74906 34522
rect 74906 34470 74908 34522
rect 74852 34468 74908 34470
rect 74956 34522 75012 34524
rect 74956 34470 74958 34522
rect 74958 34470 75010 34522
rect 75010 34470 75012 34522
rect 74956 34468 75012 34470
rect 75060 34522 75116 34524
rect 75060 34470 75062 34522
rect 75062 34470 75114 34522
rect 75114 34470 75116 34522
rect 75060 34468 75116 34470
rect 75404 34524 75460 34580
rect 74852 32954 74908 32956
rect 74852 32902 74854 32954
rect 74854 32902 74906 32954
rect 74906 32902 74908 32954
rect 74852 32900 74908 32902
rect 74956 32954 75012 32956
rect 74956 32902 74958 32954
rect 74958 32902 75010 32954
rect 75010 32902 75012 32954
rect 74956 32900 75012 32902
rect 75060 32954 75116 32956
rect 75060 32902 75062 32954
rect 75062 32902 75114 32954
rect 75114 32902 75116 32954
rect 75060 32900 75116 32902
rect 72156 32284 72212 32340
rect 69692 31836 69748 31892
rect 74852 31386 74908 31388
rect 74852 31334 74854 31386
rect 74854 31334 74906 31386
rect 74906 31334 74908 31386
rect 74852 31332 74908 31334
rect 74956 31386 75012 31388
rect 74956 31334 74958 31386
rect 74958 31334 75010 31386
rect 75010 31334 75012 31386
rect 74956 31332 75012 31334
rect 75060 31386 75116 31388
rect 75060 31334 75062 31386
rect 75062 31334 75114 31386
rect 75114 31334 75116 31386
rect 75060 31332 75116 31334
rect 74852 29818 74908 29820
rect 74852 29766 74854 29818
rect 74854 29766 74906 29818
rect 74906 29766 74908 29818
rect 74852 29764 74908 29766
rect 74956 29818 75012 29820
rect 74956 29766 74958 29818
rect 74958 29766 75010 29818
rect 75010 29766 75012 29818
rect 74956 29764 75012 29766
rect 75060 29818 75116 29820
rect 75060 29766 75062 29818
rect 75062 29766 75114 29818
rect 75114 29766 75116 29818
rect 75060 29764 75116 29766
rect 69020 28476 69076 28532
rect 74852 28250 74908 28252
rect 74852 28198 74854 28250
rect 74854 28198 74906 28250
rect 74906 28198 74908 28250
rect 74852 28196 74908 28198
rect 74956 28250 75012 28252
rect 74956 28198 74958 28250
rect 74958 28198 75010 28250
rect 75010 28198 75012 28250
rect 74956 28196 75012 28198
rect 75060 28250 75116 28252
rect 75060 28198 75062 28250
rect 75062 28198 75114 28250
rect 75114 28198 75116 28250
rect 75060 28196 75116 28198
rect 74852 26682 74908 26684
rect 74852 26630 74854 26682
rect 74854 26630 74906 26682
rect 74906 26630 74908 26682
rect 74852 26628 74908 26630
rect 74956 26682 75012 26684
rect 74956 26630 74958 26682
rect 74958 26630 75010 26682
rect 75010 26630 75012 26682
rect 74956 26628 75012 26630
rect 75060 26682 75116 26684
rect 75060 26630 75062 26682
rect 75062 26630 75114 26682
rect 75114 26630 75116 26682
rect 75060 26628 75116 26630
rect 67900 25452 67956 25508
rect 74852 25114 74908 25116
rect 74852 25062 74854 25114
rect 74854 25062 74906 25114
rect 74906 25062 74908 25114
rect 74852 25060 74908 25062
rect 74956 25114 75012 25116
rect 74956 25062 74958 25114
rect 74958 25062 75010 25114
rect 75010 25062 75012 25114
rect 74956 25060 75012 25062
rect 75060 25114 75116 25116
rect 75060 25062 75062 25114
rect 75062 25062 75114 25114
rect 75114 25062 75116 25114
rect 75060 25060 75116 25062
rect 75852 35532 75908 35588
rect 75628 34860 75684 34916
rect 75516 24668 75572 24724
rect 73052 24556 73108 24612
rect 68796 22876 68852 22932
rect 69804 20972 69860 21028
rect 68908 17724 68964 17780
rect 67340 15372 67396 15428
rect 67004 8258 67060 8260
rect 67004 8206 67006 8258
rect 67006 8206 67058 8258
rect 67058 8206 67060 8258
rect 67004 8204 67060 8206
rect 67228 7698 67284 7700
rect 67228 7646 67230 7698
rect 67230 7646 67282 7698
rect 67282 7646 67284 7698
rect 67228 7644 67284 7646
rect 66892 7532 66948 7588
rect 66108 7196 66164 7252
rect 66332 6636 66388 6692
rect 65996 6300 66052 6356
rect 66108 6130 66164 6132
rect 66108 6078 66110 6130
rect 66110 6078 66162 6130
rect 66162 6078 66164 6130
rect 66108 6076 66164 6078
rect 66108 5404 66164 5460
rect 63644 3554 63700 3556
rect 63644 3502 63646 3554
rect 63646 3502 63698 3554
rect 63698 3502 63700 3554
rect 63644 3500 63700 3502
rect 63532 3388 63588 3444
rect 64988 3500 65044 3556
rect 64876 3442 64932 3444
rect 64876 3390 64878 3442
rect 64878 3390 64930 3442
rect 64930 3390 64932 3442
rect 64876 3388 64932 3390
rect 67116 5122 67172 5124
rect 67116 5070 67118 5122
rect 67118 5070 67170 5122
rect 67170 5070 67172 5122
rect 67116 5068 67172 5070
rect 66892 4284 66948 4340
rect 66556 4172 66612 4228
rect 66556 3612 66612 3668
rect 68796 15372 68852 15428
rect 68348 8316 68404 8372
rect 67676 6690 67732 6692
rect 67676 6638 67678 6690
rect 67678 6638 67730 6690
rect 67730 6638 67732 6690
rect 67676 6636 67732 6638
rect 67564 6076 67620 6132
rect 67676 5404 67732 5460
rect 68124 6690 68180 6692
rect 68124 6638 68126 6690
rect 68126 6638 68178 6690
rect 68178 6638 68180 6690
rect 68124 6636 68180 6638
rect 68572 6636 68628 6692
rect 69356 6690 69412 6692
rect 69356 6638 69358 6690
rect 69358 6638 69410 6690
rect 69410 6638 69412 6690
rect 69356 6636 69412 6638
rect 68348 4338 68404 4340
rect 68348 4286 68350 4338
rect 68350 4286 68402 4338
rect 68402 4286 68404 4338
rect 68348 4284 68404 4286
rect 67564 3554 67620 3556
rect 67564 3502 67566 3554
rect 67566 3502 67618 3554
rect 67618 3502 67620 3554
rect 67564 3500 67620 3502
rect 67676 3388 67732 3444
rect 6412 28 6468 84
rect 69356 5292 69412 5348
rect 68908 5180 68964 5236
rect 69692 5234 69748 5236
rect 69692 5182 69694 5234
rect 69694 5182 69746 5234
rect 69746 5182 69748 5234
rect 69692 5180 69748 5182
rect 71372 20972 71428 21028
rect 69804 4956 69860 5012
rect 70140 5628 70196 5684
rect 68796 3442 68852 3444
rect 68796 3390 68798 3442
rect 68798 3390 68850 3442
rect 68850 3390 68852 3442
rect 68796 3388 68852 3390
rect 68572 28 68628 84
rect 70700 5068 70756 5124
rect 70252 4562 70308 4564
rect 70252 4510 70254 4562
rect 70254 4510 70306 4562
rect 70306 4510 70308 4562
rect 70252 4508 70308 4510
rect 71372 4732 71428 4788
rect 70700 4338 70756 4340
rect 70700 4286 70702 4338
rect 70702 4286 70754 4338
rect 70754 4286 70756 4338
rect 70700 4284 70756 4286
rect 74852 23546 74908 23548
rect 74852 23494 74854 23546
rect 74854 23494 74906 23546
rect 74906 23494 74908 23546
rect 74852 23492 74908 23494
rect 74956 23546 75012 23548
rect 74956 23494 74958 23546
rect 74958 23494 75010 23546
rect 75010 23494 75012 23546
rect 74956 23492 75012 23494
rect 75060 23546 75116 23548
rect 75060 23494 75062 23546
rect 75062 23494 75114 23546
rect 75114 23494 75116 23546
rect 75060 23492 75116 23494
rect 74852 21978 74908 21980
rect 74852 21926 74854 21978
rect 74854 21926 74906 21978
rect 74906 21926 74908 21978
rect 74852 21924 74908 21926
rect 74956 21978 75012 21980
rect 74956 21926 74958 21978
rect 74958 21926 75010 21978
rect 75010 21926 75012 21978
rect 74956 21924 75012 21926
rect 75060 21978 75116 21980
rect 75060 21926 75062 21978
rect 75062 21926 75114 21978
rect 75114 21926 75116 21978
rect 75060 21924 75116 21926
rect 74852 20410 74908 20412
rect 74852 20358 74854 20410
rect 74854 20358 74906 20410
rect 74906 20358 74908 20410
rect 74852 20356 74908 20358
rect 74956 20410 75012 20412
rect 74956 20358 74958 20410
rect 74958 20358 75010 20410
rect 75010 20358 75012 20410
rect 74956 20356 75012 20358
rect 75060 20410 75116 20412
rect 75060 20358 75062 20410
rect 75062 20358 75114 20410
rect 75114 20358 75116 20410
rect 75060 20356 75116 20358
rect 73052 4956 73108 5012
rect 74172 19404 74228 19460
rect 72604 4338 72660 4340
rect 72604 4286 72606 4338
rect 72606 4286 72658 4338
rect 72658 4286 72660 4338
rect 72604 4284 72660 4286
rect 70252 4172 70308 4228
rect 70588 3554 70644 3556
rect 70588 3502 70590 3554
rect 70590 3502 70642 3554
rect 70642 3502 70644 3554
rect 70588 3500 70644 3502
rect 71708 3554 71764 3556
rect 71708 3502 71710 3554
rect 71710 3502 71762 3554
rect 71762 3502 71764 3554
rect 71708 3500 71764 3502
rect 73612 3554 73668 3556
rect 73612 3502 73614 3554
rect 73614 3502 73666 3554
rect 73666 3502 73668 3554
rect 73612 3500 73668 3502
rect 71596 3388 71652 3444
rect 72716 3442 72772 3444
rect 72716 3390 72718 3442
rect 72718 3390 72770 3442
rect 72770 3390 72772 3442
rect 72716 3388 72772 3390
rect 72940 3388 72996 3444
rect 74852 18842 74908 18844
rect 74852 18790 74854 18842
rect 74854 18790 74906 18842
rect 74906 18790 74908 18842
rect 74852 18788 74908 18790
rect 74956 18842 75012 18844
rect 74956 18790 74958 18842
rect 74958 18790 75010 18842
rect 75010 18790 75012 18842
rect 74956 18788 75012 18790
rect 75060 18842 75116 18844
rect 75060 18790 75062 18842
rect 75062 18790 75114 18842
rect 75114 18790 75116 18842
rect 75060 18788 75116 18790
rect 74852 17274 74908 17276
rect 74852 17222 74854 17274
rect 74854 17222 74906 17274
rect 74906 17222 74908 17274
rect 74852 17220 74908 17222
rect 74956 17274 75012 17276
rect 74956 17222 74958 17274
rect 74958 17222 75010 17274
rect 75010 17222 75012 17274
rect 74956 17220 75012 17222
rect 75060 17274 75116 17276
rect 75060 17222 75062 17274
rect 75062 17222 75114 17274
rect 75114 17222 75116 17274
rect 75060 17220 75116 17222
rect 74852 15706 74908 15708
rect 74852 15654 74854 15706
rect 74854 15654 74906 15706
rect 74906 15654 74908 15706
rect 74852 15652 74908 15654
rect 74956 15706 75012 15708
rect 74956 15654 74958 15706
rect 74958 15654 75010 15706
rect 75010 15654 75012 15706
rect 74956 15652 75012 15654
rect 75060 15706 75116 15708
rect 75060 15654 75062 15706
rect 75062 15654 75114 15706
rect 75114 15654 75116 15706
rect 75060 15652 75116 15654
rect 74852 14138 74908 14140
rect 74852 14086 74854 14138
rect 74854 14086 74906 14138
rect 74906 14086 74908 14138
rect 74852 14084 74908 14086
rect 74956 14138 75012 14140
rect 74956 14086 74958 14138
rect 74958 14086 75010 14138
rect 75010 14086 75012 14138
rect 74956 14084 75012 14086
rect 75060 14138 75116 14140
rect 75060 14086 75062 14138
rect 75062 14086 75114 14138
rect 75114 14086 75116 14138
rect 75060 14084 75116 14086
rect 74852 12570 74908 12572
rect 74852 12518 74854 12570
rect 74854 12518 74906 12570
rect 74906 12518 74908 12570
rect 74852 12516 74908 12518
rect 74956 12570 75012 12572
rect 74956 12518 74958 12570
rect 74958 12518 75010 12570
rect 75010 12518 75012 12570
rect 74956 12516 75012 12518
rect 75060 12570 75116 12572
rect 75060 12518 75062 12570
rect 75062 12518 75114 12570
rect 75114 12518 75116 12570
rect 75060 12516 75116 12518
rect 76300 34972 76356 35028
rect 75964 34300 76020 34356
rect 76188 34914 76244 34916
rect 76188 34862 76190 34914
rect 76190 34862 76242 34914
rect 76242 34862 76244 34914
rect 76188 34860 76244 34862
rect 76636 34690 76692 34692
rect 76636 34638 76638 34690
rect 76638 34638 76690 34690
rect 76690 34638 76692 34690
rect 76636 34636 76692 34638
rect 76748 35420 76804 35476
rect 76076 32620 76132 32676
rect 78092 36764 78148 36820
rect 77196 35532 77252 35588
rect 77308 34914 77364 34916
rect 77308 34862 77310 34914
rect 77310 34862 77362 34914
rect 77362 34862 77364 34914
rect 77308 34860 77364 34862
rect 78764 36370 78820 36372
rect 78764 36318 78766 36370
rect 78766 36318 78818 36370
rect 78818 36318 78820 36370
rect 78764 36316 78820 36318
rect 77532 35980 77588 36036
rect 77420 34300 77476 34356
rect 76860 33964 76916 34020
rect 77196 34018 77252 34020
rect 77196 33966 77198 34018
rect 77198 33966 77250 34018
rect 77250 33966 77252 34018
rect 77196 33964 77252 33966
rect 76748 31724 76804 31780
rect 75740 11116 75796 11172
rect 74852 11002 74908 11004
rect 74852 10950 74854 11002
rect 74854 10950 74906 11002
rect 74906 10950 74908 11002
rect 74852 10948 74908 10950
rect 74956 11002 75012 11004
rect 74956 10950 74958 11002
rect 74958 10950 75010 11002
rect 75010 10950 75012 11002
rect 74956 10948 75012 10950
rect 75060 11002 75116 11004
rect 75060 10950 75062 11002
rect 75062 10950 75114 11002
rect 75114 10950 75116 11002
rect 75060 10948 75116 10950
rect 74852 9434 74908 9436
rect 74852 9382 74854 9434
rect 74854 9382 74906 9434
rect 74906 9382 74908 9434
rect 74852 9380 74908 9382
rect 74956 9434 75012 9436
rect 74956 9382 74958 9434
rect 74958 9382 75010 9434
rect 75010 9382 75012 9434
rect 74956 9380 75012 9382
rect 75060 9434 75116 9436
rect 75060 9382 75062 9434
rect 75062 9382 75114 9434
rect 75114 9382 75116 9434
rect 75060 9380 75116 9382
rect 74852 7866 74908 7868
rect 74852 7814 74854 7866
rect 74854 7814 74906 7866
rect 74906 7814 74908 7866
rect 74852 7812 74908 7814
rect 74956 7866 75012 7868
rect 74956 7814 74958 7866
rect 74958 7814 75010 7866
rect 75010 7814 75012 7866
rect 74956 7812 75012 7814
rect 75060 7866 75116 7868
rect 75060 7814 75062 7866
rect 75062 7814 75114 7866
rect 75114 7814 75116 7866
rect 75060 7812 75116 7814
rect 75628 6802 75684 6804
rect 75628 6750 75630 6802
rect 75630 6750 75682 6802
rect 75682 6750 75684 6802
rect 75628 6748 75684 6750
rect 74852 6298 74908 6300
rect 74852 6246 74854 6298
rect 74854 6246 74906 6298
rect 74906 6246 74908 6298
rect 74852 6244 74908 6246
rect 74956 6298 75012 6300
rect 74956 6246 74958 6298
rect 74958 6246 75010 6298
rect 75010 6246 75012 6298
rect 74956 6244 75012 6246
rect 75060 6298 75116 6300
rect 75060 6246 75062 6298
rect 75062 6246 75114 6298
rect 75114 6246 75116 6298
rect 75060 6244 75116 6246
rect 76412 7084 76468 7140
rect 77084 7474 77140 7476
rect 77084 7422 77086 7474
rect 77086 7422 77138 7474
rect 77138 7422 77140 7474
rect 77084 7420 77140 7422
rect 76860 7084 76916 7140
rect 78428 36258 78484 36260
rect 78428 36206 78430 36258
rect 78430 36206 78482 36258
rect 78482 36206 78484 36258
rect 78428 36204 78484 36206
rect 78540 35698 78596 35700
rect 78540 35646 78542 35698
rect 78542 35646 78594 35698
rect 78594 35646 78596 35698
rect 78540 35644 78596 35646
rect 78092 35084 78148 35140
rect 78428 35084 78484 35140
rect 77980 35026 78036 35028
rect 77980 34974 77982 35026
rect 77982 34974 78034 35026
rect 78034 34974 78036 35026
rect 77980 34972 78036 34974
rect 78204 34354 78260 34356
rect 78204 34302 78206 34354
rect 78206 34302 78258 34354
rect 78258 34302 78260 34354
rect 78204 34300 78260 34302
rect 78764 34354 78820 34356
rect 78764 34302 78766 34354
rect 78766 34302 78818 34354
rect 78818 34302 78820 34354
rect 78764 34300 78820 34302
rect 79436 36316 79492 36372
rect 79100 35644 79156 35700
rect 79212 35586 79268 35588
rect 79212 35534 79214 35586
rect 79214 35534 79266 35586
rect 79266 35534 79268 35586
rect 79212 35532 79268 35534
rect 80332 38780 80388 38836
rect 80556 37548 80612 37604
rect 80332 35980 80388 36036
rect 79884 35196 79940 35252
rect 79436 34636 79492 34692
rect 78988 34300 79044 34356
rect 79436 34300 79492 34356
rect 78204 34076 78260 34132
rect 78204 12684 78260 12740
rect 77756 6748 77812 6804
rect 77980 7084 78036 7140
rect 75740 5682 75796 5684
rect 75740 5630 75742 5682
rect 75742 5630 75794 5682
rect 75794 5630 75796 5682
rect 75740 5628 75796 5630
rect 76300 6412 76356 6468
rect 75516 5234 75572 5236
rect 75516 5182 75518 5234
rect 75518 5182 75570 5234
rect 75570 5182 75572 5234
rect 75516 5180 75572 5182
rect 75292 5068 75348 5124
rect 74852 4730 74908 4732
rect 74852 4678 74854 4730
rect 74854 4678 74906 4730
rect 74906 4678 74908 4730
rect 74852 4676 74908 4678
rect 74956 4730 75012 4732
rect 74956 4678 74958 4730
rect 74958 4678 75010 4730
rect 75010 4678 75012 4730
rect 74956 4676 75012 4678
rect 75060 4730 75116 4732
rect 75060 4678 75062 4730
rect 75062 4678 75114 4730
rect 75114 4678 75116 4730
rect 75060 4676 75116 4678
rect 74844 4338 74900 4340
rect 74844 4286 74846 4338
rect 74846 4286 74898 4338
rect 74898 4286 74900 4338
rect 74844 4284 74900 4286
rect 75628 3666 75684 3668
rect 75628 3614 75630 3666
rect 75630 3614 75682 3666
rect 75682 3614 75684 3666
rect 75628 3612 75684 3614
rect 76524 6018 76580 6020
rect 76524 5966 76526 6018
rect 76526 5966 76578 6018
rect 76578 5966 76580 6018
rect 76524 5964 76580 5966
rect 77644 5852 77700 5908
rect 77420 5180 77476 5236
rect 77756 5122 77812 5124
rect 77756 5070 77758 5122
rect 77758 5070 77810 5122
rect 77810 5070 77812 5122
rect 77756 5068 77812 5070
rect 76300 3500 76356 3556
rect 77532 3612 77588 3668
rect 74508 3442 74564 3444
rect 74508 3390 74510 3442
rect 74510 3390 74562 3442
rect 74562 3390 74564 3442
rect 74508 3388 74564 3390
rect 74956 3442 75012 3444
rect 74956 3390 74958 3442
rect 74958 3390 75010 3442
rect 75010 3390 75012 3442
rect 74956 3388 75012 3390
rect 75628 3388 75684 3444
rect 74852 3162 74908 3164
rect 74852 3110 74854 3162
rect 74854 3110 74906 3162
rect 74906 3110 74908 3162
rect 74852 3108 74908 3110
rect 74956 3162 75012 3164
rect 74956 3110 74958 3162
rect 74958 3110 75010 3162
rect 75010 3110 75012 3162
rect 74956 3108 75012 3110
rect 75060 3162 75116 3164
rect 75060 3110 75062 3162
rect 75062 3110 75114 3162
rect 75114 3110 75116 3162
rect 75060 3108 75116 3110
rect 74172 2828 74228 2884
rect 76636 3442 76692 3444
rect 76636 3390 76638 3442
rect 76638 3390 76690 3442
rect 76690 3390 76692 3442
rect 76636 3388 76692 3390
rect 76972 3388 77028 3444
rect 79772 32620 79828 32676
rect 79212 27580 79268 27636
rect 80556 35644 80612 35700
rect 80892 36764 80948 36820
rect 80780 35532 80836 35588
rect 81340 35698 81396 35700
rect 81340 35646 81342 35698
rect 81342 35646 81394 35698
rect 81394 35646 81396 35698
rect 81340 35644 81396 35646
rect 80668 34690 80724 34692
rect 80668 34638 80670 34690
rect 80670 34638 80722 34690
rect 80722 34638 80724 34690
rect 80668 34636 80724 34638
rect 82012 38444 82068 38500
rect 82012 35586 82068 35588
rect 82012 35534 82014 35586
rect 82014 35534 82066 35586
rect 82066 35534 82068 35586
rect 82012 35532 82068 35534
rect 81676 34972 81732 35028
rect 83468 36764 83524 36820
rect 84812 36764 84868 36820
rect 80444 34188 80500 34244
rect 83468 35810 83524 35812
rect 83468 35758 83470 35810
rect 83470 35758 83522 35810
rect 83522 35758 83524 35810
rect 83468 35756 83524 35758
rect 82684 35196 82740 35252
rect 82572 35026 82628 35028
rect 82572 34974 82574 35026
rect 82574 34974 82626 35026
rect 82626 34974 82628 35026
rect 82572 34972 82628 34974
rect 82348 34188 82404 34244
rect 81452 30940 81508 30996
rect 83132 34242 83188 34244
rect 83132 34190 83134 34242
rect 83134 34190 83186 34242
rect 83186 34190 83188 34242
rect 83132 34188 83188 34190
rect 83692 33516 83748 33572
rect 84028 34412 84084 34468
rect 83916 29260 83972 29316
rect 86940 37324 86996 37380
rect 85260 36764 85316 36820
rect 86156 36764 86212 36820
rect 85260 34860 85316 34916
rect 84364 29148 84420 29204
rect 84588 34412 84644 34468
rect 83804 26460 83860 26516
rect 82796 25676 82852 25732
rect 83132 26012 83188 26068
rect 80108 14252 80164 14308
rect 81452 24444 81508 24500
rect 81452 12684 81508 12740
rect 78428 7420 78484 7476
rect 78540 6748 78596 6804
rect 79100 6466 79156 6468
rect 79100 6414 79102 6466
rect 79102 6414 79154 6466
rect 79154 6414 79156 6466
rect 79100 6412 79156 6414
rect 80892 6412 80948 6468
rect 79884 6018 79940 6020
rect 79884 5966 79886 6018
rect 79886 5966 79938 6018
rect 79938 5966 79940 6018
rect 79884 5964 79940 5966
rect 78764 5906 78820 5908
rect 78764 5854 78766 5906
rect 78766 5854 78818 5906
rect 78818 5854 78820 5906
rect 78764 5852 78820 5854
rect 79436 5906 79492 5908
rect 79436 5854 79438 5906
rect 79438 5854 79490 5906
rect 79490 5854 79492 5906
rect 79436 5852 79492 5854
rect 80444 5852 80500 5908
rect 78988 5180 79044 5236
rect 78428 5068 78484 5124
rect 80444 5068 80500 5124
rect 81340 4956 81396 5012
rect 79884 4450 79940 4452
rect 79884 4398 79886 4450
rect 79886 4398 79938 4450
rect 79938 4398 79940 4450
rect 79884 4396 79940 4398
rect 80444 4450 80500 4452
rect 80444 4398 80446 4450
rect 80446 4398 80498 4450
rect 80498 4398 80500 4450
rect 80444 4396 80500 4398
rect 81340 4396 81396 4452
rect 79100 4338 79156 4340
rect 79100 4286 79102 4338
rect 79102 4286 79154 4338
rect 79154 4286 79156 4338
rect 79100 4284 79156 4286
rect 81452 3554 81508 3556
rect 81452 3502 81454 3554
rect 81454 3502 81506 3554
rect 81506 3502 81508 3554
rect 81452 3500 81508 3502
rect 78428 3442 78484 3444
rect 78428 3390 78430 3442
rect 78430 3390 78482 3442
rect 78482 3390 78484 3442
rect 78428 3388 78484 3390
rect 79324 3442 79380 3444
rect 79324 3390 79326 3442
rect 79326 3390 79378 3442
rect 79378 3390 79380 3442
rect 79324 3388 79380 3390
rect 79660 3388 79716 3444
rect 78204 3164 78260 3220
rect 80556 3442 80612 3444
rect 80556 3390 80558 3442
rect 80558 3390 80610 3442
rect 80610 3390 80612 3442
rect 80556 3388 80612 3390
rect 81004 3388 81060 3444
rect 81788 3388 81844 3444
rect 82012 3442 82068 3444
rect 82012 3390 82014 3442
rect 82014 3390 82066 3442
rect 82066 3390 82068 3442
rect 82012 3388 82068 3390
rect 82908 8092 82964 8148
rect 82908 3554 82964 3556
rect 82908 3502 82910 3554
rect 82910 3502 82962 3554
rect 82962 3502 82964 3554
rect 82908 3500 82964 3502
rect 86044 34188 86100 34244
rect 86940 36482 86996 36484
rect 86940 36430 86942 36482
rect 86942 36430 86994 36482
rect 86994 36430 86996 36482
rect 86940 36428 86996 36430
rect 87052 35532 87108 35588
rect 87276 37100 87332 37156
rect 86380 26348 86436 26404
rect 88172 38332 88228 38388
rect 87948 36482 88004 36484
rect 87948 36430 87950 36482
rect 87950 36430 88002 36482
rect 88002 36430 88004 36482
rect 87948 36428 88004 36430
rect 87388 35756 87444 35812
rect 87948 35586 88004 35588
rect 87948 35534 87950 35586
rect 87950 35534 88002 35586
rect 88002 35534 88004 35586
rect 87948 35532 88004 35534
rect 88060 35084 88116 35140
rect 89068 37548 89124 37604
rect 87388 34524 87444 34580
rect 87948 34524 88004 34580
rect 88508 33516 88564 33572
rect 89068 36876 89124 36932
rect 88956 36482 89012 36484
rect 88956 36430 88958 36482
rect 88958 36430 89010 36482
rect 89010 36430 89012 36482
rect 88956 36428 89012 36430
rect 89516 36204 89572 36260
rect 88732 34972 88788 35028
rect 88844 35084 88900 35140
rect 89292 34524 89348 34580
rect 89628 35084 89684 35140
rect 89740 36204 89796 36260
rect 89404 33628 89460 33684
rect 86604 20972 86660 21028
rect 85820 17612 85876 17668
rect 85820 11676 85876 11732
rect 85484 7980 85540 8036
rect 84588 6076 84644 6132
rect 84476 4508 84532 4564
rect 85596 5010 85652 5012
rect 85596 4958 85598 5010
rect 85598 4958 85650 5010
rect 85650 4958 85652 5010
rect 85596 4956 85652 4958
rect 85260 4508 85316 4564
rect 85372 3612 85428 3668
rect 83132 3164 83188 3220
rect 83692 3388 83748 3444
rect 84476 3442 84532 3444
rect 84476 3390 84478 3442
rect 84478 3390 84530 3442
rect 84530 3390 84532 3442
rect 84476 3388 84532 3390
rect 85036 3388 85092 3444
rect 86044 7980 86100 8036
rect 86268 7420 86324 7476
rect 85932 5068 85988 5124
rect 87052 7532 87108 7588
rect 86492 7084 86548 7140
rect 87052 6690 87108 6692
rect 87052 6638 87054 6690
rect 87054 6638 87106 6690
rect 87106 6638 87108 6690
rect 87052 6636 87108 6638
rect 86380 5122 86436 5124
rect 86380 5070 86382 5122
rect 86382 5070 86434 5122
rect 86434 5070 86436 5122
rect 86380 5068 86436 5070
rect 89068 11228 89124 11284
rect 87948 8258 88004 8260
rect 87948 8206 87950 8258
rect 87950 8206 88002 8258
rect 88002 8206 88004 8258
rect 87948 8204 88004 8206
rect 87724 7644 87780 7700
rect 87836 7586 87892 7588
rect 87836 7534 87838 7586
rect 87838 7534 87890 7586
rect 87890 7534 87892 7586
rect 87836 7532 87892 7534
rect 88508 8146 88564 8148
rect 88508 8094 88510 8146
rect 88510 8094 88562 8146
rect 88562 8094 88564 8146
rect 88508 8092 88564 8094
rect 88284 7532 88340 7588
rect 88396 7308 88452 7364
rect 86828 5180 86884 5236
rect 88508 4562 88564 4564
rect 88508 4510 88510 4562
rect 88510 4510 88562 4562
rect 88562 4510 88564 4562
rect 88508 4508 88564 4510
rect 86268 3612 86324 3668
rect 86268 3442 86324 3444
rect 86268 3390 86270 3442
rect 86270 3390 86322 3442
rect 86322 3390 86324 3442
rect 86268 3388 86324 3390
rect 86716 3442 86772 3444
rect 86716 3390 86718 3442
rect 86718 3390 86770 3442
rect 86770 3390 86772 3442
rect 86716 3388 86772 3390
rect 87724 3388 87780 3444
rect 88396 3442 88452 3444
rect 88396 3390 88398 3442
rect 88398 3390 88450 3442
rect 88450 3390 88452 3442
rect 88396 3388 88452 3390
rect 89516 33234 89572 33236
rect 89516 33182 89518 33234
rect 89518 33182 89570 33234
rect 89570 33182 89572 33234
rect 89516 33180 89572 33182
rect 89964 35810 90020 35812
rect 89964 35758 89966 35810
rect 89966 35758 90018 35810
rect 90018 35758 90020 35810
rect 89964 35756 90020 35758
rect 90188 35698 90244 35700
rect 90188 35646 90190 35698
rect 90190 35646 90242 35698
rect 90242 35646 90244 35698
rect 90188 35644 90244 35646
rect 90636 35980 90692 36036
rect 90412 35420 90468 35476
rect 90188 35026 90244 35028
rect 90188 34974 90190 35026
rect 90190 34974 90242 35026
rect 90242 34974 90244 35026
rect 90188 34972 90244 34974
rect 90300 34018 90356 34020
rect 90300 33966 90302 34018
rect 90302 33966 90354 34018
rect 90354 33966 90356 34018
rect 90300 33964 90356 33966
rect 89628 26124 89684 26180
rect 91196 36370 91252 36372
rect 91196 36318 91198 36370
rect 91198 36318 91250 36370
rect 91250 36318 91252 36370
rect 91196 36316 91252 36318
rect 90972 35420 91028 35476
rect 90636 33964 90692 34020
rect 92316 38220 92372 38276
rect 91980 36540 92036 36596
rect 91868 35980 91924 36036
rect 91532 34300 91588 34356
rect 90524 33628 90580 33684
rect 91868 35084 91924 35140
rect 92316 35980 92372 36036
rect 93262 36874 93318 36876
rect 93262 36822 93264 36874
rect 93264 36822 93316 36874
rect 93316 36822 93318 36874
rect 93262 36820 93318 36822
rect 93366 36874 93422 36876
rect 93366 36822 93368 36874
rect 93368 36822 93420 36874
rect 93420 36822 93422 36874
rect 93366 36820 93422 36822
rect 93470 36874 93526 36876
rect 93470 36822 93472 36874
rect 93472 36822 93524 36874
rect 93524 36822 93526 36874
rect 93470 36820 93526 36822
rect 92988 36428 93044 36484
rect 92764 36258 92820 36260
rect 92764 36206 92766 36258
rect 92766 36206 92818 36258
rect 92818 36206 92820 36258
rect 92764 36204 92820 36206
rect 92988 35644 93044 35700
rect 93100 36092 93156 36148
rect 92428 34972 92484 35028
rect 92428 34524 92484 34580
rect 92652 34300 92708 34356
rect 92092 33404 92148 33460
rect 93772 36092 93828 36148
rect 93548 35756 93604 35812
rect 93262 35306 93318 35308
rect 93262 35254 93264 35306
rect 93264 35254 93316 35306
rect 93316 35254 93318 35306
rect 93262 35252 93318 35254
rect 93366 35306 93422 35308
rect 93366 35254 93368 35306
rect 93368 35254 93420 35306
rect 93420 35254 93422 35306
rect 93366 35252 93422 35254
rect 93470 35306 93526 35308
rect 93470 35254 93472 35306
rect 93472 35254 93524 35306
rect 93524 35254 93526 35306
rect 93470 35252 93526 35254
rect 94220 36540 94276 36596
rect 94332 36316 94388 36372
rect 94332 35698 94388 35700
rect 94332 35646 94334 35698
rect 94334 35646 94386 35698
rect 94386 35646 94388 35698
rect 94332 35644 94388 35646
rect 93884 35196 93940 35252
rect 93996 35026 94052 35028
rect 93996 34974 93998 35026
rect 93998 34974 94050 35026
rect 94050 34974 94052 35026
rect 93996 34972 94052 34974
rect 93324 34636 93380 34692
rect 93436 34524 93492 34580
rect 93262 33738 93318 33740
rect 93262 33686 93264 33738
rect 93264 33686 93316 33738
rect 93316 33686 93318 33738
rect 93262 33684 93318 33686
rect 93366 33738 93422 33740
rect 93366 33686 93368 33738
rect 93368 33686 93420 33738
rect 93420 33686 93422 33738
rect 93366 33684 93422 33686
rect 93470 33738 93526 33740
rect 93470 33686 93472 33738
rect 93472 33686 93524 33738
rect 93524 33686 93526 33738
rect 93470 33684 93526 33686
rect 93262 32170 93318 32172
rect 93262 32118 93264 32170
rect 93264 32118 93316 32170
rect 93316 32118 93318 32170
rect 93262 32116 93318 32118
rect 93366 32170 93422 32172
rect 93366 32118 93368 32170
rect 93368 32118 93420 32170
rect 93420 32118 93422 32170
rect 93366 32116 93422 32118
rect 93470 32170 93526 32172
rect 93470 32118 93472 32170
rect 93472 32118 93524 32170
rect 93524 32118 93526 32170
rect 93470 32116 93526 32118
rect 93262 30602 93318 30604
rect 93262 30550 93264 30602
rect 93264 30550 93316 30602
rect 93316 30550 93318 30602
rect 93262 30548 93318 30550
rect 93366 30602 93422 30604
rect 93366 30550 93368 30602
rect 93368 30550 93420 30602
rect 93420 30550 93422 30602
rect 93366 30548 93422 30550
rect 93470 30602 93526 30604
rect 93470 30550 93472 30602
rect 93472 30550 93524 30602
rect 93524 30550 93526 30602
rect 93470 30548 93526 30550
rect 93262 29034 93318 29036
rect 93262 28982 93264 29034
rect 93264 28982 93316 29034
rect 93316 28982 93318 29034
rect 93262 28980 93318 28982
rect 93366 29034 93422 29036
rect 93366 28982 93368 29034
rect 93368 28982 93420 29034
rect 93420 28982 93422 29034
rect 93366 28980 93422 28982
rect 93470 29034 93526 29036
rect 93470 28982 93472 29034
rect 93472 28982 93524 29034
rect 93524 28982 93526 29034
rect 93470 28980 93526 28982
rect 91196 28812 91252 28868
rect 90860 27804 90916 27860
rect 93262 27466 93318 27468
rect 93262 27414 93264 27466
rect 93264 27414 93316 27466
rect 93316 27414 93318 27466
rect 93262 27412 93318 27414
rect 93366 27466 93422 27468
rect 93366 27414 93368 27466
rect 93368 27414 93420 27466
rect 93420 27414 93422 27466
rect 93366 27412 93422 27414
rect 93470 27466 93526 27468
rect 93470 27414 93472 27466
rect 93472 27414 93524 27466
rect 93524 27414 93526 27466
rect 93470 27412 93526 27414
rect 93884 27244 93940 27300
rect 90300 25564 90356 25620
rect 91532 26124 91588 26180
rect 93262 25898 93318 25900
rect 93262 25846 93264 25898
rect 93264 25846 93316 25898
rect 93316 25846 93318 25898
rect 93262 25844 93318 25846
rect 93366 25898 93422 25900
rect 93366 25846 93368 25898
rect 93368 25846 93420 25898
rect 93420 25846 93422 25898
rect 93366 25844 93422 25846
rect 93470 25898 93526 25900
rect 93470 25846 93472 25898
rect 93472 25846 93524 25898
rect 93524 25846 93526 25898
rect 93470 25844 93526 25846
rect 93262 24330 93318 24332
rect 93262 24278 93264 24330
rect 93264 24278 93316 24330
rect 93316 24278 93318 24330
rect 93262 24276 93318 24278
rect 93366 24330 93422 24332
rect 93366 24278 93368 24330
rect 93368 24278 93420 24330
rect 93420 24278 93422 24330
rect 93366 24276 93422 24278
rect 93470 24330 93526 24332
rect 93470 24278 93472 24330
rect 93472 24278 93524 24330
rect 93524 24278 93526 24330
rect 93470 24276 93526 24278
rect 93262 22762 93318 22764
rect 93262 22710 93264 22762
rect 93264 22710 93316 22762
rect 93316 22710 93318 22762
rect 93262 22708 93318 22710
rect 93366 22762 93422 22764
rect 93366 22710 93368 22762
rect 93368 22710 93420 22762
rect 93420 22710 93422 22762
rect 93366 22708 93422 22710
rect 93470 22762 93526 22764
rect 93470 22710 93472 22762
rect 93472 22710 93524 22762
rect 93524 22710 93526 22762
rect 93470 22708 93526 22710
rect 93262 21194 93318 21196
rect 93262 21142 93264 21194
rect 93264 21142 93316 21194
rect 93316 21142 93318 21194
rect 93262 21140 93318 21142
rect 93366 21194 93422 21196
rect 93366 21142 93368 21194
rect 93368 21142 93420 21194
rect 93420 21142 93422 21194
rect 93366 21140 93422 21142
rect 93470 21194 93526 21196
rect 93470 21142 93472 21194
rect 93472 21142 93524 21194
rect 93524 21142 93526 21194
rect 93470 21140 93526 21142
rect 93262 19626 93318 19628
rect 93262 19574 93264 19626
rect 93264 19574 93316 19626
rect 93316 19574 93318 19626
rect 93262 19572 93318 19574
rect 93366 19626 93422 19628
rect 93366 19574 93368 19626
rect 93368 19574 93420 19626
rect 93420 19574 93422 19626
rect 93366 19572 93422 19574
rect 93470 19626 93526 19628
rect 93470 19574 93472 19626
rect 93472 19574 93524 19626
rect 93524 19574 93526 19626
rect 93470 19572 93526 19574
rect 93262 18058 93318 18060
rect 93262 18006 93264 18058
rect 93264 18006 93316 18058
rect 93316 18006 93318 18058
rect 93262 18004 93318 18006
rect 93366 18058 93422 18060
rect 93366 18006 93368 18058
rect 93368 18006 93420 18058
rect 93420 18006 93422 18058
rect 93366 18004 93422 18006
rect 93470 18058 93526 18060
rect 93470 18006 93472 18058
rect 93472 18006 93524 18058
rect 93524 18006 93526 18058
rect 93470 18004 93526 18006
rect 93262 16490 93318 16492
rect 93262 16438 93264 16490
rect 93264 16438 93316 16490
rect 93316 16438 93318 16490
rect 93262 16436 93318 16438
rect 93366 16490 93422 16492
rect 93366 16438 93368 16490
rect 93368 16438 93420 16490
rect 93420 16438 93422 16490
rect 93366 16436 93422 16438
rect 93470 16490 93526 16492
rect 93470 16438 93472 16490
rect 93472 16438 93524 16490
rect 93524 16438 93526 16490
rect 93470 16436 93526 16438
rect 93262 14922 93318 14924
rect 93262 14870 93264 14922
rect 93264 14870 93316 14922
rect 93316 14870 93318 14922
rect 93262 14868 93318 14870
rect 93366 14922 93422 14924
rect 93366 14870 93368 14922
rect 93368 14870 93420 14922
rect 93420 14870 93422 14922
rect 93366 14868 93422 14870
rect 93470 14922 93526 14924
rect 93470 14870 93472 14922
rect 93472 14870 93524 14922
rect 93524 14870 93526 14922
rect 93470 14868 93526 14870
rect 93262 13354 93318 13356
rect 93262 13302 93264 13354
rect 93264 13302 93316 13354
rect 93316 13302 93318 13354
rect 93262 13300 93318 13302
rect 93366 13354 93422 13356
rect 93366 13302 93368 13354
rect 93368 13302 93420 13354
rect 93420 13302 93422 13354
rect 93366 13300 93422 13302
rect 93470 13354 93526 13356
rect 93470 13302 93472 13354
rect 93472 13302 93524 13354
rect 93524 13302 93526 13354
rect 93470 13300 93526 13302
rect 91532 11676 91588 11732
rect 93262 11786 93318 11788
rect 93262 11734 93264 11786
rect 93264 11734 93316 11786
rect 93316 11734 93318 11786
rect 93262 11732 93318 11734
rect 93366 11786 93422 11788
rect 93366 11734 93368 11786
rect 93368 11734 93420 11786
rect 93420 11734 93422 11786
rect 93366 11732 93422 11734
rect 93470 11786 93526 11788
rect 93470 11734 93472 11786
rect 93472 11734 93524 11786
rect 93524 11734 93526 11786
rect 93470 11732 93526 11734
rect 93262 10218 93318 10220
rect 93262 10166 93264 10218
rect 93264 10166 93316 10218
rect 93316 10166 93318 10218
rect 93262 10164 93318 10166
rect 93366 10218 93422 10220
rect 93366 10166 93368 10218
rect 93368 10166 93420 10218
rect 93420 10166 93422 10218
rect 93366 10164 93422 10166
rect 93470 10218 93526 10220
rect 93470 10166 93472 10218
rect 93472 10166 93524 10218
rect 93524 10166 93526 10218
rect 93470 10164 93526 10166
rect 93262 8650 93318 8652
rect 93262 8598 93264 8650
rect 93264 8598 93316 8650
rect 93316 8598 93318 8650
rect 93262 8596 93318 8598
rect 93366 8650 93422 8652
rect 93366 8598 93368 8650
rect 93368 8598 93420 8650
rect 93420 8598 93422 8650
rect 93366 8596 93422 8598
rect 93470 8650 93526 8652
rect 93470 8598 93472 8650
rect 93472 8598 93524 8650
rect 93524 8598 93526 8650
rect 93470 8596 93526 8598
rect 89404 8258 89460 8260
rect 89404 8206 89406 8258
rect 89406 8206 89458 8258
rect 89458 8206 89460 8258
rect 89404 8204 89460 8206
rect 90748 8204 90804 8260
rect 89852 8146 89908 8148
rect 89852 8094 89854 8146
rect 89854 8094 89906 8146
rect 89906 8094 89908 8146
rect 89852 8092 89908 8094
rect 90076 8092 90132 8148
rect 89180 7698 89236 7700
rect 89180 7646 89182 7698
rect 89182 7646 89234 7698
rect 89234 7646 89236 7698
rect 89180 7644 89236 7646
rect 89628 7362 89684 7364
rect 89628 7310 89630 7362
rect 89630 7310 89682 7362
rect 89682 7310 89684 7362
rect 89628 7308 89684 7310
rect 89404 4956 89460 5012
rect 89628 5628 89684 5684
rect 89292 4508 89348 4564
rect 89964 4956 90020 5012
rect 89852 3724 89908 3780
rect 95900 36316 95956 36372
rect 95116 35084 95172 35140
rect 95564 35196 95620 35252
rect 96572 36594 96628 36596
rect 96572 36542 96574 36594
rect 96574 36542 96626 36594
rect 96626 36542 96628 36594
rect 96572 36540 96628 36542
rect 96908 36540 96964 36596
rect 97244 36876 97300 36932
rect 96012 35084 96068 35140
rect 96124 34972 96180 35028
rect 96236 34636 96292 34692
rect 98364 36594 98420 36596
rect 98364 36542 98366 36594
rect 98366 36542 98418 36594
rect 98418 36542 98420 36594
rect 98364 36540 98420 36542
rect 97244 35644 97300 35700
rect 97356 34972 97412 35028
rect 95452 33852 95508 33908
rect 96012 33180 96068 33236
rect 96348 31164 96404 31220
rect 95116 28364 95172 28420
rect 96572 27692 96628 27748
rect 94780 8258 94836 8260
rect 94780 8206 94782 8258
rect 94782 8206 94834 8258
rect 94834 8206 94836 8258
rect 94780 8204 94836 8206
rect 93772 8146 93828 8148
rect 93772 8094 93774 8146
rect 93774 8094 93826 8146
rect 93826 8094 93828 8146
rect 93772 8092 93828 8094
rect 92540 7980 92596 8036
rect 93100 7980 93156 8036
rect 94892 8092 94948 8148
rect 93262 7082 93318 7084
rect 93262 7030 93264 7082
rect 93264 7030 93316 7082
rect 93316 7030 93318 7082
rect 93262 7028 93318 7030
rect 93366 7082 93422 7084
rect 93366 7030 93368 7082
rect 93368 7030 93420 7082
rect 93420 7030 93422 7082
rect 93366 7028 93422 7030
rect 93470 7082 93526 7084
rect 93470 7030 93472 7082
rect 93472 7030 93524 7082
rect 93524 7030 93526 7082
rect 93470 7028 93526 7030
rect 94444 7420 94500 7476
rect 96124 8258 96180 8260
rect 96124 8206 96126 8258
rect 96126 8206 96178 8258
rect 96178 8206 96180 8258
rect 96124 8204 96180 8206
rect 95564 8092 95620 8148
rect 95340 7980 95396 8036
rect 95116 7644 95172 7700
rect 96012 7698 96068 7700
rect 96012 7646 96014 7698
rect 96014 7646 96066 7698
rect 96066 7646 96068 7698
rect 96012 7644 96068 7646
rect 96460 7474 96516 7476
rect 96460 7422 96462 7474
rect 96462 7422 96514 7474
rect 96514 7422 96516 7474
rect 96460 7420 96516 7422
rect 93262 5514 93318 5516
rect 93262 5462 93264 5514
rect 93264 5462 93316 5514
rect 93316 5462 93318 5514
rect 93262 5460 93318 5462
rect 93366 5514 93422 5516
rect 93366 5462 93368 5514
rect 93368 5462 93420 5514
rect 93420 5462 93422 5514
rect 93366 5460 93422 5462
rect 93470 5514 93526 5516
rect 93470 5462 93472 5514
rect 93472 5462 93524 5514
rect 93524 5462 93526 5514
rect 93470 5460 93526 5462
rect 93884 5122 93940 5124
rect 93884 5070 93886 5122
rect 93886 5070 93938 5122
rect 93938 5070 93940 5122
rect 93884 5068 93940 5070
rect 94556 5122 94612 5124
rect 94556 5070 94558 5122
rect 94558 5070 94610 5122
rect 94610 5070 94612 5122
rect 94556 5068 94612 5070
rect 95452 6690 95508 6692
rect 95452 6638 95454 6690
rect 95454 6638 95506 6690
rect 95506 6638 95508 6690
rect 95452 6636 95508 6638
rect 95676 6636 95732 6692
rect 95340 6412 95396 6468
rect 95564 6076 95620 6132
rect 95788 6412 95844 6468
rect 90412 4956 90468 5012
rect 90860 4898 90916 4900
rect 90860 4846 90862 4898
rect 90862 4846 90914 4898
rect 90914 4846 90916 4898
rect 90860 4844 90916 4846
rect 93262 3946 93318 3948
rect 93262 3894 93264 3946
rect 93264 3894 93316 3946
rect 93316 3894 93318 3946
rect 93262 3892 93318 3894
rect 93366 3946 93422 3948
rect 93366 3894 93368 3946
rect 93368 3894 93420 3946
rect 93420 3894 93422 3946
rect 93366 3892 93422 3894
rect 93470 3946 93526 3948
rect 93470 3894 93472 3946
rect 93472 3894 93524 3946
rect 93524 3894 93526 3946
rect 93470 3892 93526 3894
rect 93212 3612 93268 3668
rect 89068 3276 89124 3332
rect 89180 3388 89236 3444
rect 90188 3442 90244 3444
rect 90188 3390 90190 3442
rect 90190 3390 90242 3442
rect 90242 3390 90244 3442
rect 90188 3388 90244 3390
rect 90636 3442 90692 3444
rect 90636 3390 90638 3442
rect 90638 3390 90690 3442
rect 90690 3390 90692 3442
rect 90636 3388 90692 3390
rect 91756 3388 91812 3444
rect 89852 3330 89908 3332
rect 89852 3278 89854 3330
rect 89854 3278 89906 3330
rect 89906 3278 89908 3330
rect 89852 3276 89908 3278
rect 89852 2492 89908 2548
rect 92316 3442 92372 3444
rect 92316 3390 92318 3442
rect 92318 3390 92370 3442
rect 92370 3390 92372 3442
rect 92316 3388 92372 3390
rect 93100 3388 93156 3444
rect 94668 3666 94724 3668
rect 94668 3614 94670 3666
rect 94670 3614 94722 3666
rect 94722 3614 94724 3666
rect 94668 3612 94724 3614
rect 93772 3442 93828 3444
rect 93772 3390 93774 3442
rect 93774 3390 93826 3442
rect 93826 3390 93828 3442
rect 93772 3388 93828 3390
rect 97132 27132 97188 27188
rect 100492 36540 100548 36596
rect 101052 36652 101108 36708
rect 100604 35980 100660 36036
rect 99820 35922 99876 35924
rect 99820 35870 99822 35922
rect 99822 35870 99874 35922
rect 99874 35870 99876 35922
rect 99820 35868 99876 35870
rect 102172 36988 102228 37044
rect 101052 35756 101108 35812
rect 98812 35196 98868 35252
rect 99596 35196 99652 35252
rect 100044 35196 100100 35252
rect 98364 29596 98420 29652
rect 99932 34636 99988 34692
rect 98028 26236 98084 26292
rect 98140 19292 98196 19348
rect 98140 11788 98196 11844
rect 96684 8034 96740 8036
rect 96684 7982 96686 8034
rect 96686 7982 96738 8034
rect 96738 7982 96740 8034
rect 96684 7980 96740 7982
rect 98028 7980 98084 8036
rect 95564 3276 95620 3332
rect 95788 3388 95844 3444
rect 94108 3164 94164 3220
rect 94108 2604 94164 2660
rect 96348 3442 96404 3444
rect 96348 3390 96350 3442
rect 96350 3390 96402 3442
rect 96402 3390 96404 3442
rect 96348 3388 96404 3390
rect 96572 5628 96628 5684
rect 97244 5628 97300 5684
rect 97244 3554 97300 3556
rect 97244 3502 97246 3554
rect 97246 3502 97298 3554
rect 97298 3502 97300 3554
rect 97244 3500 97300 3502
rect 96460 3164 96516 3220
rect 97132 3388 97188 3444
rect 97580 3388 97636 3444
rect 97804 3442 97860 3444
rect 97804 3390 97806 3442
rect 97806 3390 97858 3442
rect 97858 3390 97860 3442
rect 97804 3388 97860 3390
rect 98924 7420 98980 7476
rect 98364 5628 98420 5684
rect 98924 5628 98980 5684
rect 98700 3554 98756 3556
rect 98700 3502 98702 3554
rect 98702 3502 98754 3554
rect 98754 3502 98756 3554
rect 98700 3500 98756 3502
rect 99820 3388 99876 3444
rect 101612 35810 101668 35812
rect 101612 35758 101614 35810
rect 101614 35758 101666 35810
rect 101666 35758 101668 35810
rect 101612 35756 101668 35758
rect 101612 34690 101668 34692
rect 101612 34638 101614 34690
rect 101614 34638 101666 34690
rect 101666 34638 101668 34690
rect 101612 34636 101668 34638
rect 100716 33740 100772 33796
rect 100716 32732 100772 32788
rect 101164 28028 101220 28084
rect 101612 32732 101668 32788
rect 102396 36594 102452 36596
rect 102396 36542 102398 36594
rect 102398 36542 102450 36594
rect 102450 36542 102452 36594
rect 102396 36540 102452 36542
rect 103740 37996 103796 38052
rect 103180 36540 103236 36596
rect 103516 37100 103572 37156
rect 102284 35756 102340 35812
rect 102844 35810 102900 35812
rect 102844 35758 102846 35810
rect 102846 35758 102898 35810
rect 102898 35758 102900 35810
rect 102844 35756 102900 35758
rect 102172 34188 102228 34244
rect 103292 34802 103348 34804
rect 103292 34750 103294 34802
rect 103294 34750 103346 34802
rect 103346 34750 103348 34802
rect 103292 34748 103348 34750
rect 102956 34636 103012 34692
rect 103740 35756 103796 35812
rect 102508 33628 102564 33684
rect 102508 33292 102564 33348
rect 102620 33068 102676 33124
rect 104188 37100 104244 37156
rect 104412 36594 104468 36596
rect 104412 36542 104414 36594
rect 104414 36542 104466 36594
rect 104466 36542 104468 36594
rect 104412 36540 104468 36542
rect 104972 34972 105028 35028
rect 104300 33740 104356 33796
rect 103740 31052 103796 31108
rect 102060 29484 102116 29540
rect 103292 24668 103348 24724
rect 105196 32620 105252 32676
rect 105532 35420 105588 35476
rect 106204 36428 106260 36484
rect 106428 36316 106484 36372
rect 107212 36316 107268 36372
rect 106316 35810 106372 35812
rect 106316 35758 106318 35810
rect 106318 35758 106370 35810
rect 106370 35758 106372 35810
rect 106316 35756 106372 35758
rect 105532 34412 105588 34468
rect 105084 30828 105140 30884
rect 105868 35026 105924 35028
rect 105868 34974 105870 35026
rect 105870 34974 105922 35026
rect 105922 34974 105924 35026
rect 105868 34972 105924 34974
rect 105644 34188 105700 34244
rect 106092 33628 106148 33684
rect 105756 33516 105812 33572
rect 106540 35532 106596 35588
rect 106428 34242 106484 34244
rect 106428 34190 106430 34242
rect 106430 34190 106482 34242
rect 106482 34190 106484 34242
rect 106428 34188 106484 34190
rect 106204 33516 106260 33572
rect 105532 29932 105588 29988
rect 106652 24556 106708 24612
rect 104412 17724 104468 17780
rect 104188 17612 104244 17668
rect 104188 11788 104244 11844
rect 103292 8876 103348 8932
rect 101276 3724 101332 3780
rect 100380 3442 100436 3444
rect 100380 3390 100382 3442
rect 100382 3390 100434 3442
rect 100434 3390 100436 3442
rect 100380 3388 100436 3390
rect 101164 3388 101220 3444
rect 99932 2716 99988 2772
rect 102956 7980 103012 8036
rect 102508 6636 102564 6692
rect 102508 5852 102564 5908
rect 103964 8034 104020 8036
rect 103964 7982 103966 8034
rect 103966 7982 104018 8034
rect 104018 7982 104020 8034
rect 103964 7980 104020 7982
rect 104076 7586 104132 7588
rect 104076 7534 104078 7586
rect 104078 7534 104130 7586
rect 104130 7534 104132 7586
rect 104076 7532 104132 7534
rect 102732 5628 102788 5684
rect 102620 5122 102676 5124
rect 102620 5070 102622 5122
rect 102622 5070 102674 5122
rect 102674 5070 102676 5122
rect 102620 5068 102676 5070
rect 102732 3724 102788 3780
rect 103068 7308 103124 7364
rect 103516 7362 103572 7364
rect 103516 7310 103518 7362
rect 103518 7310 103570 7362
rect 103570 7310 103572 7362
rect 103516 7308 103572 7310
rect 104412 6636 104468 6692
rect 105756 8258 105812 8260
rect 105756 8206 105758 8258
rect 105758 8206 105810 8258
rect 105810 8206 105812 8258
rect 105756 8204 105812 8206
rect 106652 8204 106708 8260
rect 105532 8092 105588 8148
rect 105980 8146 106036 8148
rect 105980 8094 105982 8146
rect 105982 8094 106034 8146
rect 106034 8094 106036 8146
rect 105980 8092 106036 8094
rect 105420 7532 105476 7588
rect 106316 7980 106372 8036
rect 105980 7644 106036 7700
rect 105756 7474 105812 7476
rect 105756 7422 105758 7474
rect 105758 7422 105810 7474
rect 105810 7422 105812 7474
rect 105756 7420 105812 7422
rect 106988 35084 107044 35140
rect 106988 34748 107044 34804
rect 107324 35586 107380 35588
rect 107324 35534 107326 35586
rect 107326 35534 107378 35586
rect 107378 35534 107380 35586
rect 107324 35532 107380 35534
rect 107324 35196 107380 35252
rect 107548 35756 107604 35812
rect 108668 36482 108724 36484
rect 108668 36430 108670 36482
rect 108670 36430 108722 36482
rect 108722 36430 108724 36482
rect 108668 36428 108724 36430
rect 106764 7420 106820 7476
rect 106876 33068 106932 33124
rect 106316 7308 106372 7364
rect 105980 6690 106036 6692
rect 105980 6638 105982 6690
rect 105982 6638 106034 6690
rect 106034 6638 106036 6690
rect 105980 6636 106036 6638
rect 104748 6524 104804 6580
rect 106092 6524 106148 6580
rect 105756 6412 105812 6468
rect 103740 6076 103796 6132
rect 104412 6130 104468 6132
rect 104412 6078 104414 6130
rect 104414 6078 104466 6130
rect 104466 6078 104468 6130
rect 104412 6076 104468 6078
rect 104524 5852 104580 5908
rect 103180 5628 103236 5684
rect 103628 5628 103684 5684
rect 104300 5628 104356 5684
rect 103964 5068 104020 5124
rect 105308 5906 105364 5908
rect 105308 5854 105310 5906
rect 105310 5854 105362 5906
rect 105362 5854 105364 5906
rect 105308 5852 105364 5854
rect 105308 5068 105364 5124
rect 106652 5852 106708 5908
rect 106764 5122 106820 5124
rect 106764 5070 106766 5122
rect 106766 5070 106818 5122
rect 106818 5070 106820 5122
rect 106764 5068 106820 5070
rect 105756 4338 105812 4340
rect 105756 4286 105758 4338
rect 105758 4286 105810 4338
rect 105810 4286 105812 4338
rect 105756 4284 105812 4286
rect 103068 3612 103124 3668
rect 102956 3500 103012 3556
rect 105308 3554 105364 3556
rect 105308 3502 105310 3554
rect 105310 3502 105362 3554
rect 105362 3502 105364 3554
rect 105308 3500 105364 3502
rect 101612 3388 101668 3444
rect 101836 3442 101892 3444
rect 101836 3390 101838 3442
rect 101838 3390 101890 3442
rect 101890 3390 101892 3442
rect 101836 3388 101892 3390
rect 103852 3388 103908 3444
rect 102172 3330 102228 3332
rect 102172 3278 102174 3330
rect 102174 3278 102226 3330
rect 102226 3278 102228 3330
rect 102172 3276 102228 3278
rect 101500 2828 101556 2884
rect 104412 3442 104468 3444
rect 104412 3390 104414 3442
rect 104414 3390 104466 3442
rect 104466 3390 104468 3442
rect 104412 3388 104468 3390
rect 105196 3388 105252 3444
rect 106204 3442 106260 3444
rect 106204 3390 106206 3442
rect 106206 3390 106258 3442
rect 106258 3390 106260 3442
rect 106204 3388 106260 3390
rect 106652 3442 106708 3444
rect 106652 3390 106654 3442
rect 106654 3390 106706 3442
rect 106706 3390 106708 3442
rect 106652 3388 106708 3390
rect 108332 35308 108388 35364
rect 108668 36092 108724 36148
rect 108556 34636 108612 34692
rect 108780 35084 108836 35140
rect 109340 36482 109396 36484
rect 109340 36430 109342 36482
rect 109342 36430 109394 36482
rect 109394 36430 109396 36482
rect 109340 36428 109396 36430
rect 109228 36092 109284 36148
rect 109004 35084 109060 35140
rect 109228 35420 109284 35476
rect 109228 34412 109284 34468
rect 108780 33852 108836 33908
rect 110236 37884 110292 37940
rect 110124 36428 110180 36484
rect 109452 34412 109508 34468
rect 107996 33122 108052 33124
rect 107996 33070 107998 33122
rect 107998 33070 108050 33122
rect 108050 33070 108052 33122
rect 107996 33068 108052 33070
rect 108332 33516 108388 33572
rect 109452 33516 109508 33572
rect 107548 32508 107604 32564
rect 109116 31500 109172 31556
rect 107100 8258 107156 8260
rect 107100 8206 107102 8258
rect 107102 8206 107154 8258
rect 107154 8206 107156 8258
rect 107100 8204 107156 8206
rect 107100 7698 107156 7700
rect 107100 7646 107102 7698
rect 107102 7646 107154 7698
rect 107154 7646 107156 7698
rect 107100 7644 107156 7646
rect 107548 7474 107604 7476
rect 107548 7422 107550 7474
rect 107550 7422 107602 7474
rect 107602 7422 107604 7474
rect 107548 7420 107604 7422
rect 107100 6466 107156 6468
rect 107100 6414 107102 6466
rect 107102 6414 107154 6466
rect 107154 6414 107156 6466
rect 107100 6412 107156 6414
rect 107212 4284 107268 4340
rect 108220 6130 108276 6132
rect 108220 6078 108222 6130
rect 108222 6078 108274 6130
rect 108274 6078 108276 6130
rect 108220 6076 108276 6078
rect 109228 6130 109284 6132
rect 109228 6078 109230 6130
rect 109230 6078 109282 6130
rect 109282 6078 109284 6130
rect 109228 6076 109284 6078
rect 108332 5964 108388 6020
rect 107548 5180 107604 5236
rect 109340 6018 109396 6020
rect 109340 5966 109342 6018
rect 109342 5966 109394 6018
rect 109394 5966 109396 6018
rect 109340 5964 109396 5966
rect 108444 4508 108500 4564
rect 107436 3724 107492 3780
rect 107884 4172 107940 4228
rect 108108 3778 108164 3780
rect 108108 3726 108110 3778
rect 108110 3726 108162 3778
rect 108162 3726 108164 3778
rect 108108 3724 108164 3726
rect 108780 3836 108836 3892
rect 109788 35084 109844 35140
rect 109900 34412 109956 34468
rect 110012 33404 110068 33460
rect 110348 36652 110404 36708
rect 111132 38780 111188 38836
rect 110348 35474 110404 35476
rect 110348 35422 110350 35474
rect 110350 35422 110402 35474
rect 110402 35422 110404 35474
rect 110348 35420 110404 35422
rect 110124 33292 110180 33348
rect 110796 34690 110852 34692
rect 110796 34638 110798 34690
rect 110798 34638 110850 34690
rect 110850 34638 110852 34690
rect 110796 34636 110852 34638
rect 110796 33404 110852 33460
rect 112140 36540 112196 36596
rect 112252 36652 112308 36708
rect 111356 35922 111412 35924
rect 111356 35870 111358 35922
rect 111358 35870 111410 35922
rect 111410 35870 111412 35922
rect 111356 35868 111412 35870
rect 111672 36090 111728 36092
rect 111672 36038 111674 36090
rect 111674 36038 111726 36090
rect 111726 36038 111728 36090
rect 111672 36036 111728 36038
rect 111776 36090 111832 36092
rect 111776 36038 111778 36090
rect 111778 36038 111830 36090
rect 111830 36038 111832 36090
rect 111776 36036 111832 36038
rect 111880 36090 111936 36092
rect 111880 36038 111882 36090
rect 111882 36038 111934 36090
rect 111934 36038 111936 36090
rect 111880 36036 111936 36038
rect 112252 35810 112308 35812
rect 112252 35758 112254 35810
rect 112254 35758 112306 35810
rect 112306 35758 112308 35810
rect 112252 35756 112308 35758
rect 111468 35196 111524 35252
rect 111580 34636 111636 34692
rect 111244 34524 111300 34580
rect 111672 34522 111728 34524
rect 111672 34470 111674 34522
rect 111674 34470 111726 34522
rect 111726 34470 111728 34522
rect 111672 34468 111728 34470
rect 111776 34522 111832 34524
rect 111776 34470 111778 34522
rect 111778 34470 111830 34522
rect 111830 34470 111832 34522
rect 111776 34468 111832 34470
rect 111880 34522 111936 34524
rect 111880 34470 111882 34522
rect 111882 34470 111934 34522
rect 111934 34470 111936 34522
rect 111880 34468 111936 34470
rect 112812 35420 112868 35476
rect 111020 33516 111076 33572
rect 110908 33068 110964 33124
rect 111020 32732 111076 32788
rect 109676 25452 109732 25508
rect 110236 6018 110292 6020
rect 110236 5966 110238 6018
rect 110238 5966 110290 6018
rect 110290 5966 110292 6018
rect 110236 5964 110292 5966
rect 109228 5234 109284 5236
rect 109228 5182 109230 5234
rect 109230 5182 109282 5234
rect 109282 5182 109284 5234
rect 109228 5180 109284 5182
rect 109564 5180 109620 5236
rect 110236 5628 110292 5684
rect 109452 4226 109508 4228
rect 109452 4174 109454 4226
rect 109454 4174 109506 4226
rect 109506 4174 109508 4226
rect 109452 4172 109508 4174
rect 110124 3836 110180 3892
rect 109004 3500 109060 3556
rect 109228 3554 109284 3556
rect 109228 3502 109230 3554
rect 109230 3502 109282 3554
rect 109282 3502 109284 3554
rect 109228 3500 109284 3502
rect 109900 3442 109956 3444
rect 109900 3390 109902 3442
rect 109902 3390 109954 3442
rect 109954 3390 109956 3442
rect 109900 3388 109956 3390
rect 112252 33516 112308 33572
rect 111672 32954 111728 32956
rect 111672 32902 111674 32954
rect 111674 32902 111726 32954
rect 111726 32902 111728 32954
rect 111672 32900 111728 32902
rect 111776 32954 111832 32956
rect 111776 32902 111778 32954
rect 111778 32902 111830 32954
rect 111830 32902 111832 32954
rect 111776 32900 111832 32902
rect 111880 32954 111936 32956
rect 111880 32902 111882 32954
rect 111882 32902 111934 32954
rect 111934 32902 111936 32954
rect 111880 32900 111936 32902
rect 111672 31386 111728 31388
rect 111672 31334 111674 31386
rect 111674 31334 111726 31386
rect 111726 31334 111728 31386
rect 111672 31332 111728 31334
rect 111776 31386 111832 31388
rect 111776 31334 111778 31386
rect 111778 31334 111830 31386
rect 111830 31334 111832 31386
rect 111776 31332 111832 31334
rect 111880 31386 111936 31388
rect 111880 31334 111882 31386
rect 111882 31334 111934 31386
rect 111934 31334 111936 31386
rect 111880 31332 111936 31334
rect 111672 29818 111728 29820
rect 111672 29766 111674 29818
rect 111674 29766 111726 29818
rect 111726 29766 111728 29818
rect 111672 29764 111728 29766
rect 111776 29818 111832 29820
rect 111776 29766 111778 29818
rect 111778 29766 111830 29818
rect 111830 29766 111832 29818
rect 111776 29764 111832 29766
rect 111880 29818 111936 29820
rect 111880 29766 111882 29818
rect 111882 29766 111934 29818
rect 111934 29766 111936 29818
rect 111880 29764 111936 29766
rect 111672 28250 111728 28252
rect 111672 28198 111674 28250
rect 111674 28198 111726 28250
rect 111726 28198 111728 28250
rect 111672 28196 111728 28198
rect 111776 28250 111832 28252
rect 111776 28198 111778 28250
rect 111778 28198 111830 28250
rect 111830 28198 111832 28250
rect 111776 28196 111832 28198
rect 111880 28250 111936 28252
rect 111880 28198 111882 28250
rect 111882 28198 111934 28250
rect 111934 28198 111936 28250
rect 111880 28196 111936 28198
rect 111672 26682 111728 26684
rect 111672 26630 111674 26682
rect 111674 26630 111726 26682
rect 111726 26630 111728 26682
rect 111672 26628 111728 26630
rect 111776 26682 111832 26684
rect 111776 26630 111778 26682
rect 111778 26630 111830 26682
rect 111830 26630 111832 26682
rect 111776 26628 111832 26630
rect 111880 26682 111936 26684
rect 111880 26630 111882 26682
rect 111882 26630 111934 26682
rect 111934 26630 111936 26682
rect 111880 26628 111936 26630
rect 111468 26012 111524 26068
rect 111672 25114 111728 25116
rect 111672 25062 111674 25114
rect 111674 25062 111726 25114
rect 111726 25062 111728 25114
rect 111672 25060 111728 25062
rect 111776 25114 111832 25116
rect 111776 25062 111778 25114
rect 111778 25062 111830 25114
rect 111830 25062 111832 25114
rect 111776 25060 111832 25062
rect 111880 25114 111936 25116
rect 111880 25062 111882 25114
rect 111882 25062 111934 25114
rect 111934 25062 111936 25114
rect 111880 25060 111936 25062
rect 111672 23546 111728 23548
rect 111672 23494 111674 23546
rect 111674 23494 111726 23546
rect 111726 23494 111728 23546
rect 111672 23492 111728 23494
rect 111776 23546 111832 23548
rect 111776 23494 111778 23546
rect 111778 23494 111830 23546
rect 111830 23494 111832 23546
rect 111776 23492 111832 23494
rect 111880 23546 111936 23548
rect 111880 23494 111882 23546
rect 111882 23494 111934 23546
rect 111934 23494 111936 23546
rect 111880 23492 111936 23494
rect 111672 21978 111728 21980
rect 111672 21926 111674 21978
rect 111674 21926 111726 21978
rect 111726 21926 111728 21978
rect 111672 21924 111728 21926
rect 111776 21978 111832 21980
rect 111776 21926 111778 21978
rect 111778 21926 111830 21978
rect 111830 21926 111832 21978
rect 111776 21924 111832 21926
rect 111880 21978 111936 21980
rect 111880 21926 111882 21978
rect 111882 21926 111934 21978
rect 111934 21926 111936 21978
rect 111880 21924 111936 21926
rect 111672 20410 111728 20412
rect 111672 20358 111674 20410
rect 111674 20358 111726 20410
rect 111726 20358 111728 20410
rect 111672 20356 111728 20358
rect 111776 20410 111832 20412
rect 111776 20358 111778 20410
rect 111778 20358 111830 20410
rect 111830 20358 111832 20410
rect 111776 20356 111832 20358
rect 111880 20410 111936 20412
rect 111880 20358 111882 20410
rect 111882 20358 111934 20410
rect 111934 20358 111936 20410
rect 111880 20356 111936 20358
rect 111672 18842 111728 18844
rect 111672 18790 111674 18842
rect 111674 18790 111726 18842
rect 111726 18790 111728 18842
rect 111672 18788 111728 18790
rect 111776 18842 111832 18844
rect 111776 18790 111778 18842
rect 111778 18790 111830 18842
rect 111830 18790 111832 18842
rect 111776 18788 111832 18790
rect 111880 18842 111936 18844
rect 111880 18790 111882 18842
rect 111882 18790 111934 18842
rect 111934 18790 111936 18842
rect 111880 18788 111936 18790
rect 111672 17274 111728 17276
rect 111672 17222 111674 17274
rect 111674 17222 111726 17274
rect 111726 17222 111728 17274
rect 111672 17220 111728 17222
rect 111776 17274 111832 17276
rect 111776 17222 111778 17274
rect 111778 17222 111830 17274
rect 111830 17222 111832 17274
rect 111776 17220 111832 17222
rect 111880 17274 111936 17276
rect 111880 17222 111882 17274
rect 111882 17222 111934 17274
rect 111934 17222 111936 17274
rect 111880 17220 111936 17222
rect 111672 15706 111728 15708
rect 111672 15654 111674 15706
rect 111674 15654 111726 15706
rect 111726 15654 111728 15706
rect 111672 15652 111728 15654
rect 111776 15706 111832 15708
rect 111776 15654 111778 15706
rect 111778 15654 111830 15706
rect 111830 15654 111832 15706
rect 111776 15652 111832 15654
rect 111880 15706 111936 15708
rect 111880 15654 111882 15706
rect 111882 15654 111934 15706
rect 111934 15654 111936 15706
rect 111880 15652 111936 15654
rect 111672 14138 111728 14140
rect 111672 14086 111674 14138
rect 111674 14086 111726 14138
rect 111726 14086 111728 14138
rect 111672 14084 111728 14086
rect 111776 14138 111832 14140
rect 111776 14086 111778 14138
rect 111778 14086 111830 14138
rect 111830 14086 111832 14138
rect 111776 14084 111832 14086
rect 111880 14138 111936 14140
rect 111880 14086 111882 14138
rect 111882 14086 111934 14138
rect 111934 14086 111936 14138
rect 111880 14084 111936 14086
rect 111672 12570 111728 12572
rect 111672 12518 111674 12570
rect 111674 12518 111726 12570
rect 111726 12518 111728 12570
rect 111672 12516 111728 12518
rect 111776 12570 111832 12572
rect 111776 12518 111778 12570
rect 111778 12518 111830 12570
rect 111830 12518 111832 12570
rect 111776 12516 111832 12518
rect 111880 12570 111936 12572
rect 111880 12518 111882 12570
rect 111882 12518 111934 12570
rect 111934 12518 111936 12570
rect 111880 12516 111936 12518
rect 111672 11002 111728 11004
rect 111672 10950 111674 11002
rect 111674 10950 111726 11002
rect 111726 10950 111728 11002
rect 111672 10948 111728 10950
rect 111776 11002 111832 11004
rect 111776 10950 111778 11002
rect 111778 10950 111830 11002
rect 111830 10950 111832 11002
rect 111776 10948 111832 10950
rect 111880 11002 111936 11004
rect 111880 10950 111882 11002
rect 111882 10950 111934 11002
rect 111934 10950 111936 11002
rect 111880 10948 111936 10950
rect 111672 9434 111728 9436
rect 111672 9382 111674 9434
rect 111674 9382 111726 9434
rect 111726 9382 111728 9434
rect 111672 9380 111728 9382
rect 111776 9434 111832 9436
rect 111776 9382 111778 9434
rect 111778 9382 111830 9434
rect 111830 9382 111832 9434
rect 111776 9380 111832 9382
rect 111880 9434 111936 9436
rect 111880 9382 111882 9434
rect 111882 9382 111934 9434
rect 111934 9382 111936 9434
rect 111880 9380 111936 9382
rect 111672 7866 111728 7868
rect 111672 7814 111674 7866
rect 111674 7814 111726 7866
rect 111726 7814 111728 7866
rect 111672 7812 111728 7814
rect 111776 7866 111832 7868
rect 111776 7814 111778 7866
rect 111778 7814 111830 7866
rect 111830 7814 111832 7866
rect 111776 7812 111832 7814
rect 111880 7866 111936 7868
rect 111880 7814 111882 7866
rect 111882 7814 111934 7866
rect 111934 7814 111936 7866
rect 111880 7812 111936 7814
rect 111672 6298 111728 6300
rect 111672 6246 111674 6298
rect 111674 6246 111726 6298
rect 111726 6246 111728 6298
rect 111672 6244 111728 6246
rect 111776 6298 111832 6300
rect 111776 6246 111778 6298
rect 111778 6246 111830 6298
rect 111830 6246 111832 6298
rect 111776 6244 111832 6246
rect 111880 6298 111936 6300
rect 111880 6246 111882 6298
rect 111882 6246 111934 6298
rect 111934 6246 111936 6298
rect 111880 6244 111936 6246
rect 110796 6076 110852 6132
rect 110908 5628 110964 5684
rect 112364 5906 112420 5908
rect 112364 5854 112366 5906
rect 112366 5854 112418 5906
rect 112418 5854 112420 5906
rect 112364 5852 112420 5854
rect 111580 5794 111636 5796
rect 111580 5742 111582 5794
rect 111582 5742 111634 5794
rect 111634 5742 111636 5794
rect 111580 5740 111636 5742
rect 111020 5292 111076 5348
rect 110460 4396 110516 4452
rect 111356 5234 111412 5236
rect 111356 5182 111358 5234
rect 111358 5182 111410 5234
rect 111410 5182 111412 5234
rect 111356 5180 111412 5182
rect 111672 4730 111728 4732
rect 111672 4678 111674 4730
rect 111674 4678 111726 4730
rect 111726 4678 111728 4730
rect 111672 4676 111728 4678
rect 111776 4730 111832 4732
rect 111776 4678 111778 4730
rect 111778 4678 111830 4730
rect 111830 4678 111832 4730
rect 111776 4676 111832 4678
rect 111880 4730 111936 4732
rect 111880 4678 111882 4730
rect 111882 4678 111934 4730
rect 111934 4678 111936 4730
rect 111880 4676 111936 4678
rect 110908 4562 110964 4564
rect 110908 4510 110910 4562
rect 110910 4510 110962 4562
rect 110962 4510 110964 4562
rect 110908 4508 110964 4510
rect 113148 37660 113204 37716
rect 113372 35868 113428 35924
rect 113484 35698 113540 35700
rect 113484 35646 113486 35698
rect 113486 35646 113538 35698
rect 113538 35646 113540 35698
rect 113484 35644 113540 35646
rect 114044 36594 114100 36596
rect 114044 36542 114046 36594
rect 114046 36542 114098 36594
rect 114098 36542 114100 36594
rect 114044 36540 114100 36542
rect 115724 36540 115780 36596
rect 116620 36594 116676 36596
rect 116620 36542 116622 36594
rect 116622 36542 116674 36594
rect 116674 36542 116676 36594
rect 116620 36540 116676 36542
rect 114268 35756 114324 35812
rect 113932 35532 113988 35588
rect 114828 35586 114884 35588
rect 114828 35534 114830 35586
rect 114830 35534 114882 35586
rect 114882 35534 114884 35586
rect 114828 35532 114884 35534
rect 115052 35420 115108 35476
rect 113036 35084 113092 35140
rect 114380 35084 114436 35140
rect 114380 34802 114436 34804
rect 114380 34750 114382 34802
rect 114382 34750 114434 34802
rect 114434 34750 114436 34802
rect 114380 34748 114436 34750
rect 113484 34690 113540 34692
rect 113484 34638 113486 34690
rect 113486 34638 113538 34690
rect 113538 34638 113540 34690
rect 113484 34636 113540 34638
rect 115500 35644 115556 35700
rect 115500 35084 115556 35140
rect 115836 34802 115892 34804
rect 115836 34750 115838 34802
rect 115838 34750 115890 34802
rect 115890 34750 115892 34802
rect 115836 34748 115892 34750
rect 116844 36204 116900 36260
rect 116284 35810 116340 35812
rect 116284 35758 116286 35810
rect 116286 35758 116338 35810
rect 116338 35758 116340 35810
rect 116284 35756 116340 35758
rect 115948 34636 116004 34692
rect 117516 35532 117572 35588
rect 117628 36204 117684 36260
rect 117516 35084 117572 35140
rect 114044 34188 114100 34244
rect 113932 33740 113988 33796
rect 114380 33740 114436 33796
rect 113596 27916 113652 27972
rect 116284 26124 116340 26180
rect 113148 12684 113204 12740
rect 113372 12572 113428 12628
rect 113260 5906 113316 5908
rect 113260 5854 113262 5906
rect 113262 5854 113314 5906
rect 113314 5854 113316 5906
rect 113260 5852 113316 5854
rect 112812 4508 112868 4564
rect 111356 4450 111412 4452
rect 111356 4398 111358 4450
rect 111358 4398 111410 4450
rect 111410 4398 111412 4450
rect 111356 4396 111412 4398
rect 115388 7532 115444 7588
rect 116620 7586 116676 7588
rect 116620 7534 116622 7586
rect 116622 7534 116674 7586
rect 116674 7534 116676 7586
rect 116620 7532 116676 7534
rect 116396 7474 116452 7476
rect 116396 7422 116398 7474
rect 116398 7422 116450 7474
rect 116450 7422 116452 7474
rect 116396 7420 116452 7422
rect 115052 7196 115108 7252
rect 114268 6748 114324 6804
rect 113708 6412 113764 6468
rect 110684 3500 110740 3556
rect 111468 3442 111524 3444
rect 111468 3390 111470 3442
rect 111470 3390 111522 3442
rect 111522 3390 111524 3442
rect 111468 3388 111524 3390
rect 111672 3162 111728 3164
rect 111672 3110 111674 3162
rect 111674 3110 111726 3162
rect 111726 3110 111728 3162
rect 111672 3108 111728 3110
rect 111776 3162 111832 3164
rect 111776 3110 111778 3162
rect 111778 3110 111830 3162
rect 111830 3110 111832 3162
rect 111776 3108 111832 3110
rect 111880 3162 111936 3164
rect 111880 3110 111882 3162
rect 111882 3110 111934 3162
rect 111934 3110 111936 3162
rect 111880 3108 111936 3110
rect 113372 4060 113428 4116
rect 113260 2492 113316 2548
rect 114716 6466 114772 6468
rect 114716 6414 114718 6466
rect 114718 6414 114770 6466
rect 114770 6414 114772 6466
rect 114716 6412 114772 6414
rect 114940 5964 114996 6020
rect 116956 7308 117012 7364
rect 116060 7250 116116 7252
rect 116060 7198 116062 7250
rect 116062 7198 116114 7250
rect 116114 7198 116116 7250
rect 116060 7196 116116 7198
rect 115388 5740 115444 5796
rect 118076 36428 118132 36484
rect 118748 37772 118804 37828
rect 117740 35756 117796 35812
rect 118412 35586 118468 35588
rect 118412 35534 118414 35586
rect 118414 35534 118466 35586
rect 118466 35534 118468 35586
rect 118412 35532 118468 35534
rect 117852 35084 117908 35140
rect 118076 34412 118132 34468
rect 118076 33740 118132 33796
rect 118188 32956 118244 33012
rect 118636 35084 118692 35140
rect 119532 36482 119588 36484
rect 119532 36430 119534 36482
rect 119534 36430 119586 36482
rect 119586 36430 119588 36482
rect 119532 36428 119588 36430
rect 119868 35922 119924 35924
rect 119868 35870 119870 35922
rect 119870 35870 119922 35922
rect 119922 35870 119924 35922
rect 119868 35868 119924 35870
rect 121548 37436 121604 37492
rect 121100 36764 121156 36820
rect 121324 35868 121380 35924
rect 119532 35420 119588 35476
rect 119308 33740 119364 33796
rect 118524 12572 118580 12628
rect 117740 7474 117796 7476
rect 117740 7422 117742 7474
rect 117742 7422 117794 7474
rect 117794 7422 117796 7474
rect 117740 7420 117796 7422
rect 117516 6748 117572 6804
rect 117180 6300 117236 6356
rect 114940 5234 114996 5236
rect 114940 5182 114942 5234
rect 114942 5182 114994 5234
rect 114994 5182 114996 5234
rect 114940 5180 114996 5182
rect 114380 5068 114436 5124
rect 115500 5234 115556 5236
rect 115500 5182 115502 5234
rect 115502 5182 115554 5234
rect 115554 5182 115556 5234
rect 115500 5180 115556 5182
rect 116284 5234 116340 5236
rect 116284 5182 116286 5234
rect 116286 5182 116338 5234
rect 116338 5182 116340 5234
rect 116284 5180 116340 5182
rect 115612 5068 115668 5124
rect 114380 4338 114436 4340
rect 114380 4286 114382 4338
rect 114382 4286 114434 4338
rect 114434 4286 114436 4338
rect 114380 4284 114436 4286
rect 114828 4956 114884 5012
rect 116172 5122 116228 5124
rect 116172 5070 116174 5122
rect 116174 5070 116226 5122
rect 116226 5070 116228 5122
rect 116172 5068 116228 5070
rect 116956 5234 117012 5236
rect 116956 5182 116958 5234
rect 116958 5182 117010 5234
rect 117010 5182 117012 5234
rect 116956 5180 117012 5182
rect 116732 4396 116788 4452
rect 114828 4060 114884 4116
rect 117068 3948 117124 4004
rect 115724 3666 115780 3668
rect 115724 3614 115726 3666
rect 115726 3614 115778 3666
rect 115778 3614 115780 3666
rect 115724 3612 115780 3614
rect 115948 3388 116004 3444
rect 116508 3442 116564 3444
rect 116508 3390 116510 3442
rect 116510 3390 116562 3442
rect 116562 3390 116564 3442
rect 116508 3388 116564 3390
rect 118300 7532 118356 7588
rect 118188 7362 118244 7364
rect 118188 7310 118190 7362
rect 118190 7310 118242 7362
rect 118242 7310 118244 7362
rect 118188 7308 118244 7310
rect 117852 5180 117908 5236
rect 117740 5010 117796 5012
rect 117740 4958 117742 5010
rect 117742 4958 117794 5010
rect 117794 4958 117796 5010
rect 117740 4956 117796 4958
rect 117180 3612 117236 3668
rect 117068 2940 117124 2996
rect 118524 5346 118580 5348
rect 118524 5294 118526 5346
rect 118526 5294 118578 5346
rect 118578 5294 118580 5346
rect 118524 5292 118580 5294
rect 119868 35084 119924 35140
rect 119644 33180 119700 33236
rect 120428 35084 120484 35140
rect 121996 35532 122052 35588
rect 121884 34636 121940 34692
rect 120316 27692 120372 27748
rect 122892 36540 122948 36596
rect 123116 38556 123172 38612
rect 122444 36316 122500 36372
rect 122332 35922 122388 35924
rect 122332 35870 122334 35922
rect 122334 35870 122386 35922
rect 122386 35870 122388 35922
rect 122332 35868 122388 35870
rect 122108 34860 122164 34916
rect 123452 36258 123508 36260
rect 123452 36206 123454 36258
rect 123454 36206 123506 36258
rect 123506 36206 123508 36258
rect 123452 36204 123508 36206
rect 123116 35756 123172 35812
rect 123676 35644 123732 35700
rect 122780 35586 122836 35588
rect 122780 35534 122782 35586
rect 122782 35534 122834 35586
rect 122834 35534 122836 35586
rect 122780 35532 122836 35534
rect 123564 35474 123620 35476
rect 123564 35422 123566 35474
rect 123566 35422 123618 35474
rect 123618 35422 123620 35474
rect 123564 35420 123620 35422
rect 122668 34914 122724 34916
rect 122668 34862 122670 34914
rect 122670 34862 122722 34914
rect 122722 34862 122724 34914
rect 122668 34860 122724 34862
rect 122108 34636 122164 34692
rect 123004 34354 123060 34356
rect 123004 34302 123006 34354
rect 123006 34302 123058 34354
rect 123058 34302 123060 34354
rect 123004 34300 123060 34302
rect 123340 34300 123396 34356
rect 123900 35474 123956 35476
rect 123900 35422 123902 35474
rect 123902 35422 123954 35474
rect 123954 35422 123956 35474
rect 123900 35420 123956 35422
rect 124012 34860 124068 34916
rect 124124 35756 124180 35812
rect 123788 34076 123844 34132
rect 123564 34018 123620 34020
rect 123564 33966 123566 34018
rect 123566 33966 123618 34018
rect 123618 33966 123620 34018
rect 123564 33964 123620 33966
rect 124460 35810 124516 35812
rect 124460 35758 124462 35810
rect 124462 35758 124514 35810
rect 124514 35758 124516 35810
rect 124460 35756 124516 35758
rect 125244 35868 125300 35924
rect 124684 35756 124740 35812
rect 125356 35698 125412 35700
rect 125356 35646 125358 35698
rect 125358 35646 125410 35698
rect 125410 35646 125412 35698
rect 125356 35644 125412 35646
rect 124572 35532 124628 35588
rect 125132 35420 125188 35476
rect 124796 34860 124852 34916
rect 124348 33964 124404 34020
rect 125244 34914 125300 34916
rect 125244 34862 125246 34914
rect 125246 34862 125298 34914
rect 125298 34862 125300 34914
rect 125244 34860 125300 34862
rect 126028 36594 126084 36596
rect 126028 36542 126030 36594
rect 126030 36542 126082 36594
rect 126082 36542 126084 36594
rect 126028 36540 126084 36542
rect 126476 36540 126532 36596
rect 126252 35810 126308 35812
rect 126252 35758 126254 35810
rect 126254 35758 126306 35810
rect 126306 35758 126308 35810
rect 126252 35756 126308 35758
rect 127932 36594 127988 36596
rect 127932 36542 127934 36594
rect 127934 36542 127986 36594
rect 127986 36542 127988 36594
rect 127932 36540 127988 36542
rect 128268 36540 128324 36596
rect 128156 36204 128212 36260
rect 127372 35586 127428 35588
rect 127372 35534 127374 35586
rect 127374 35534 127426 35586
rect 127426 35534 127428 35586
rect 127372 35532 127428 35534
rect 127260 35308 127316 35364
rect 125580 34860 125636 34916
rect 126588 34860 126644 34916
rect 125580 34130 125636 34132
rect 125580 34078 125582 34130
rect 125582 34078 125634 34130
rect 125634 34078 125636 34130
rect 125580 34076 125636 34078
rect 125020 33852 125076 33908
rect 125916 31612 125972 31668
rect 123564 30044 123620 30100
rect 126476 33964 126532 34020
rect 126476 33516 126532 33572
rect 126140 28476 126196 28532
rect 121996 17612 122052 17668
rect 120764 11116 120820 11172
rect 120764 8316 120820 8372
rect 121884 8370 121940 8372
rect 121884 8318 121886 8370
rect 121886 8318 121938 8370
rect 121938 8318 121940 8370
rect 121884 8316 121940 8318
rect 123116 8930 123172 8932
rect 123116 8878 123118 8930
rect 123118 8878 123170 8930
rect 123170 8878 123172 8930
rect 123116 8876 123172 8878
rect 124124 8930 124180 8932
rect 124124 8878 124126 8930
rect 124126 8878 124178 8930
rect 124178 8878 124180 8930
rect 124124 8876 124180 8878
rect 124348 8876 124404 8932
rect 123564 8428 123620 8484
rect 122780 8370 122836 8372
rect 122780 8318 122782 8370
rect 122782 8318 122834 8370
rect 122834 8318 122836 8370
rect 122780 8316 122836 8318
rect 124124 8428 124180 8484
rect 124908 8876 124964 8932
rect 125468 8930 125524 8932
rect 125468 8878 125470 8930
rect 125470 8878 125522 8930
rect 125522 8878 125524 8930
rect 125468 8876 125524 8878
rect 124796 8316 124852 8372
rect 125916 8316 125972 8372
rect 123788 8204 123844 8260
rect 125244 8258 125300 8260
rect 125244 8206 125246 8258
rect 125246 8206 125298 8258
rect 125298 8206 125300 8258
rect 125244 8204 125300 8206
rect 123452 8146 123508 8148
rect 123452 8094 123454 8146
rect 123454 8094 123506 8146
rect 123506 8094 123508 8146
rect 123452 8092 123508 8094
rect 124348 8092 124404 8148
rect 123116 7980 123172 8036
rect 122668 6636 122724 6692
rect 120204 5852 120260 5908
rect 121996 5906 122052 5908
rect 121996 5854 121998 5906
rect 121998 5854 122050 5906
rect 122050 5854 122052 5906
rect 121996 5852 122052 5854
rect 119532 5292 119588 5348
rect 121212 5292 121268 5348
rect 120204 4956 120260 5012
rect 121324 5068 121380 5124
rect 120876 4956 120932 5012
rect 118524 4338 118580 4340
rect 118524 4286 118526 4338
rect 118526 4286 118578 4338
rect 118578 4286 118580 4338
rect 118524 4284 118580 4286
rect 120876 4284 120932 4340
rect 121548 4284 121604 4340
rect 122220 4338 122276 4340
rect 122220 4286 122222 4338
rect 122222 4286 122274 4338
rect 122274 4286 122276 4338
rect 122220 4284 122276 4286
rect 118300 3948 118356 4004
rect 119308 3948 119364 4004
rect 121436 3612 121492 3668
rect 119980 3388 120036 3444
rect 120540 3442 120596 3444
rect 120540 3390 120542 3442
rect 120542 3390 120594 3442
rect 120594 3390 120596 3442
rect 120540 3388 120596 3390
rect 121324 3388 121380 3444
rect 121772 3388 121828 3444
rect 121996 3442 122052 3444
rect 121996 3390 121998 3442
rect 121998 3390 122050 3442
rect 122050 3390 122052 3442
rect 121996 3388 122052 3390
rect 122444 5906 122500 5908
rect 122444 5854 122446 5906
rect 122446 5854 122498 5906
rect 122498 5854 122500 5906
rect 122444 5852 122500 5854
rect 123340 7868 123396 7924
rect 123340 7084 123396 7140
rect 122892 4338 122948 4340
rect 122892 4286 122894 4338
rect 122894 4286 122946 4338
rect 122946 4286 122948 4338
rect 122892 4284 122948 4286
rect 125020 8034 125076 8036
rect 125020 7982 125022 8034
rect 125022 7982 125074 8034
rect 125074 7982 125076 8034
rect 125020 7980 125076 7982
rect 125916 8034 125972 8036
rect 125916 7982 125918 8034
rect 125918 7982 125970 8034
rect 125970 7982 125972 8034
rect 125916 7980 125972 7982
rect 125916 7756 125972 7812
rect 125804 7698 125860 7700
rect 125804 7646 125806 7698
rect 125806 7646 125858 7698
rect 125858 7646 125860 7698
rect 125804 7644 125860 7646
rect 126140 6860 126196 6916
rect 124908 6690 124964 6692
rect 124908 6638 124910 6690
rect 124910 6638 124962 6690
rect 124962 6638 124964 6690
rect 124908 6636 124964 6638
rect 123788 6466 123844 6468
rect 123788 6414 123790 6466
rect 123790 6414 123842 6466
rect 123842 6414 123844 6466
rect 123788 6412 123844 6414
rect 125244 5852 125300 5908
rect 123900 5292 123956 5348
rect 123788 4508 123844 4564
rect 123340 3666 123396 3668
rect 123340 3614 123342 3666
rect 123342 3614 123394 3666
rect 123394 3614 123396 3666
rect 123340 3612 123396 3614
rect 124348 5234 124404 5236
rect 124348 5182 124350 5234
rect 124350 5182 124402 5234
rect 124402 5182 124404 5234
rect 124348 5180 124404 5182
rect 124908 5122 124964 5124
rect 124908 5070 124910 5122
rect 124910 5070 124962 5122
rect 124962 5070 124964 5122
rect 124908 5068 124964 5070
rect 125244 5068 125300 5124
rect 125580 6130 125636 6132
rect 125580 6078 125582 6130
rect 125582 6078 125634 6130
rect 125634 6078 125636 6130
rect 125580 6076 125636 6078
rect 126364 7250 126420 7252
rect 126364 7198 126366 7250
rect 126366 7198 126418 7250
rect 126418 7198 126420 7250
rect 126364 7196 126420 7198
rect 126252 6636 126308 6692
rect 125804 5628 125860 5684
rect 125468 4732 125524 4788
rect 126364 4226 126420 4228
rect 126364 4174 126366 4226
rect 126366 4174 126418 4226
rect 126418 4174 126420 4226
rect 126364 4172 126420 4174
rect 125692 3724 125748 3780
rect 125356 3500 125412 3556
rect 124012 3388 124068 3444
rect 124572 3442 124628 3444
rect 124572 3390 124574 3442
rect 124574 3390 124626 3442
rect 124626 3390 124628 3442
rect 124572 3388 124628 3390
rect 126140 3554 126196 3556
rect 126140 3502 126142 3554
rect 126142 3502 126194 3554
rect 126194 3502 126196 3554
rect 126140 3500 126196 3502
rect 127036 34914 127092 34916
rect 127036 34862 127038 34914
rect 127038 34862 127090 34914
rect 127090 34862 127092 34914
rect 127036 34860 127092 34862
rect 126924 34018 126980 34020
rect 126924 33966 126926 34018
rect 126926 33966 126978 34018
rect 126978 33966 126980 34018
rect 126924 33964 126980 33966
rect 127484 34860 127540 34916
rect 127932 35698 127988 35700
rect 127932 35646 127934 35698
rect 127934 35646 127986 35698
rect 127986 35646 127988 35698
rect 127932 35644 127988 35646
rect 127708 34636 127764 34692
rect 127372 33516 127428 33572
rect 126812 33292 126868 33348
rect 128044 35084 128100 35140
rect 129052 35698 129108 35700
rect 129052 35646 129054 35698
rect 129054 35646 129106 35698
rect 129106 35646 129108 35698
rect 129052 35644 129108 35646
rect 128828 34914 128884 34916
rect 128828 34862 128830 34914
rect 128830 34862 128882 34914
rect 128882 34862 128884 34914
rect 128828 34860 128884 34862
rect 130844 37212 130900 37268
rect 129724 36594 129780 36596
rect 129724 36542 129726 36594
rect 129726 36542 129778 36594
rect 129778 36542 129780 36594
rect 129724 36540 129780 36542
rect 129388 34914 129444 34916
rect 129388 34862 129390 34914
rect 129390 34862 129442 34914
rect 129442 34862 129444 34914
rect 129388 34860 129444 34862
rect 129612 36316 129668 36372
rect 130082 36874 130138 36876
rect 130082 36822 130084 36874
rect 130084 36822 130136 36874
rect 130136 36822 130138 36874
rect 130082 36820 130138 36822
rect 130186 36874 130242 36876
rect 130186 36822 130188 36874
rect 130188 36822 130240 36874
rect 130240 36822 130242 36874
rect 130186 36820 130242 36822
rect 130290 36874 130346 36876
rect 130290 36822 130292 36874
rect 130292 36822 130344 36874
rect 130344 36822 130346 36874
rect 130290 36820 130346 36822
rect 131852 36876 131908 36932
rect 131292 36204 131348 36260
rect 130844 35810 130900 35812
rect 130844 35758 130846 35810
rect 130846 35758 130898 35810
rect 130898 35758 130900 35810
rect 130844 35756 130900 35758
rect 130060 35698 130116 35700
rect 130060 35646 130062 35698
rect 130062 35646 130114 35698
rect 130114 35646 130116 35698
rect 130060 35644 130116 35646
rect 130082 35306 130138 35308
rect 130082 35254 130084 35306
rect 130084 35254 130136 35306
rect 130136 35254 130138 35306
rect 130082 35252 130138 35254
rect 130186 35306 130242 35308
rect 130186 35254 130188 35306
rect 130188 35254 130240 35306
rect 130240 35254 130242 35306
rect 130186 35252 130242 35254
rect 130290 35306 130346 35308
rect 130290 35254 130292 35306
rect 130292 35254 130344 35306
rect 130344 35254 130346 35306
rect 130290 35252 130346 35254
rect 131068 35196 131124 35252
rect 131292 35644 131348 35700
rect 129948 34860 130004 34916
rect 130284 34354 130340 34356
rect 130284 34302 130286 34354
rect 130286 34302 130338 34354
rect 130338 34302 130340 34354
rect 130284 34300 130340 34302
rect 129164 34188 129220 34244
rect 128604 33404 128660 33460
rect 128716 33516 128772 33572
rect 128268 33068 128324 33124
rect 130060 33964 130116 34020
rect 130082 33738 130138 33740
rect 130082 33686 130084 33738
rect 130084 33686 130136 33738
rect 130136 33686 130138 33738
rect 130082 33684 130138 33686
rect 130186 33738 130242 33740
rect 130186 33686 130188 33738
rect 130188 33686 130240 33738
rect 130240 33686 130242 33738
rect 130186 33684 130242 33686
rect 130290 33738 130346 33740
rect 130290 33686 130292 33738
rect 130292 33686 130344 33738
rect 130344 33686 130346 33738
rect 130290 33684 130346 33686
rect 129276 33516 129332 33572
rect 129612 33234 129668 33236
rect 129612 33182 129614 33234
rect 129614 33182 129666 33234
rect 129666 33182 129668 33234
rect 129612 33180 129668 33182
rect 129052 33068 129108 33124
rect 130172 32956 130228 33012
rect 130082 32170 130138 32172
rect 130082 32118 130084 32170
rect 130084 32118 130136 32170
rect 130136 32118 130138 32170
rect 130082 32116 130138 32118
rect 130186 32170 130242 32172
rect 130186 32118 130188 32170
rect 130188 32118 130240 32170
rect 130240 32118 130242 32170
rect 130186 32116 130242 32118
rect 130290 32170 130346 32172
rect 130290 32118 130292 32170
rect 130292 32118 130344 32170
rect 130344 32118 130346 32170
rect 130290 32116 130346 32118
rect 128156 31948 128212 32004
rect 130082 30602 130138 30604
rect 130082 30550 130084 30602
rect 130084 30550 130136 30602
rect 130136 30550 130138 30602
rect 130082 30548 130138 30550
rect 130186 30602 130242 30604
rect 130186 30550 130188 30602
rect 130188 30550 130240 30602
rect 130240 30550 130242 30602
rect 130186 30548 130242 30550
rect 130290 30602 130346 30604
rect 130290 30550 130292 30602
rect 130292 30550 130344 30602
rect 130344 30550 130346 30602
rect 130290 30548 130346 30550
rect 130082 29034 130138 29036
rect 130082 28982 130084 29034
rect 130084 28982 130136 29034
rect 130136 28982 130138 29034
rect 130082 28980 130138 28982
rect 130186 29034 130242 29036
rect 130186 28982 130188 29034
rect 130188 28982 130240 29034
rect 130240 28982 130242 29034
rect 130186 28980 130242 28982
rect 130290 29034 130346 29036
rect 130290 28982 130292 29034
rect 130292 28982 130344 29034
rect 130344 28982 130346 29034
rect 130290 28980 130346 28982
rect 130082 27466 130138 27468
rect 130082 27414 130084 27466
rect 130084 27414 130136 27466
rect 130136 27414 130138 27466
rect 130082 27412 130138 27414
rect 130186 27466 130242 27468
rect 130186 27414 130188 27466
rect 130188 27414 130240 27466
rect 130240 27414 130242 27466
rect 130186 27412 130242 27414
rect 130290 27466 130346 27468
rect 130290 27414 130292 27466
rect 130292 27414 130344 27466
rect 130344 27414 130346 27466
rect 130290 27412 130346 27414
rect 128156 26796 128212 26852
rect 130082 25898 130138 25900
rect 130082 25846 130084 25898
rect 130084 25846 130136 25898
rect 130136 25846 130138 25898
rect 130082 25844 130138 25846
rect 130186 25898 130242 25900
rect 130186 25846 130188 25898
rect 130188 25846 130240 25898
rect 130240 25846 130242 25898
rect 130186 25844 130242 25846
rect 130290 25898 130346 25900
rect 130290 25846 130292 25898
rect 130292 25846 130344 25898
rect 130344 25846 130346 25898
rect 130290 25844 130346 25846
rect 130082 24330 130138 24332
rect 130082 24278 130084 24330
rect 130084 24278 130136 24330
rect 130136 24278 130138 24330
rect 130082 24276 130138 24278
rect 130186 24330 130242 24332
rect 130186 24278 130188 24330
rect 130188 24278 130240 24330
rect 130240 24278 130242 24330
rect 130186 24276 130242 24278
rect 130290 24330 130346 24332
rect 130290 24278 130292 24330
rect 130292 24278 130344 24330
rect 130344 24278 130346 24330
rect 130290 24276 130346 24278
rect 130082 22762 130138 22764
rect 130082 22710 130084 22762
rect 130084 22710 130136 22762
rect 130136 22710 130138 22762
rect 130082 22708 130138 22710
rect 130186 22762 130242 22764
rect 130186 22710 130188 22762
rect 130188 22710 130240 22762
rect 130240 22710 130242 22762
rect 130186 22708 130242 22710
rect 130290 22762 130346 22764
rect 130290 22710 130292 22762
rect 130292 22710 130344 22762
rect 130344 22710 130346 22762
rect 130290 22708 130346 22710
rect 130082 21194 130138 21196
rect 130082 21142 130084 21194
rect 130084 21142 130136 21194
rect 130136 21142 130138 21194
rect 130082 21140 130138 21142
rect 130186 21194 130242 21196
rect 130186 21142 130188 21194
rect 130188 21142 130240 21194
rect 130240 21142 130242 21194
rect 130186 21140 130242 21142
rect 130290 21194 130346 21196
rect 130290 21142 130292 21194
rect 130292 21142 130344 21194
rect 130344 21142 130346 21194
rect 130290 21140 130346 21142
rect 130082 19626 130138 19628
rect 130082 19574 130084 19626
rect 130084 19574 130136 19626
rect 130136 19574 130138 19626
rect 130082 19572 130138 19574
rect 130186 19626 130242 19628
rect 130186 19574 130188 19626
rect 130188 19574 130240 19626
rect 130240 19574 130242 19626
rect 130186 19572 130242 19574
rect 130290 19626 130346 19628
rect 130290 19574 130292 19626
rect 130292 19574 130344 19626
rect 130344 19574 130346 19626
rect 130290 19572 130346 19574
rect 130082 18058 130138 18060
rect 130082 18006 130084 18058
rect 130084 18006 130136 18058
rect 130136 18006 130138 18058
rect 130082 18004 130138 18006
rect 130186 18058 130242 18060
rect 130186 18006 130188 18058
rect 130188 18006 130240 18058
rect 130240 18006 130242 18058
rect 130186 18004 130242 18006
rect 130290 18058 130346 18060
rect 130290 18006 130292 18058
rect 130292 18006 130344 18058
rect 130344 18006 130346 18058
rect 130290 18004 130346 18006
rect 130082 16490 130138 16492
rect 130082 16438 130084 16490
rect 130084 16438 130136 16490
rect 130136 16438 130138 16490
rect 130082 16436 130138 16438
rect 130186 16490 130242 16492
rect 130186 16438 130188 16490
rect 130188 16438 130240 16490
rect 130240 16438 130242 16490
rect 130186 16436 130242 16438
rect 130290 16490 130346 16492
rect 130290 16438 130292 16490
rect 130292 16438 130344 16490
rect 130344 16438 130346 16490
rect 130290 16436 130346 16438
rect 130082 14922 130138 14924
rect 130082 14870 130084 14922
rect 130084 14870 130136 14922
rect 130136 14870 130138 14922
rect 130082 14868 130138 14870
rect 130186 14922 130242 14924
rect 130186 14870 130188 14922
rect 130188 14870 130240 14922
rect 130240 14870 130242 14922
rect 130186 14868 130242 14870
rect 130290 14922 130346 14924
rect 130290 14870 130292 14922
rect 130292 14870 130344 14922
rect 130344 14870 130346 14922
rect 130290 14868 130346 14870
rect 130082 13354 130138 13356
rect 130082 13302 130084 13354
rect 130084 13302 130136 13354
rect 130136 13302 130138 13354
rect 130082 13300 130138 13302
rect 130186 13354 130242 13356
rect 130186 13302 130188 13354
rect 130188 13302 130240 13354
rect 130240 13302 130242 13354
rect 130186 13300 130242 13302
rect 130290 13354 130346 13356
rect 130290 13302 130292 13354
rect 130292 13302 130344 13354
rect 130344 13302 130346 13354
rect 130290 13300 130346 13302
rect 130082 11786 130138 11788
rect 130082 11734 130084 11786
rect 130084 11734 130136 11786
rect 130136 11734 130138 11786
rect 130082 11732 130138 11734
rect 130186 11786 130242 11788
rect 130186 11734 130188 11786
rect 130188 11734 130240 11786
rect 130240 11734 130242 11786
rect 130186 11732 130242 11734
rect 130290 11786 130346 11788
rect 130290 11734 130292 11786
rect 130292 11734 130344 11786
rect 130344 11734 130346 11786
rect 130290 11732 130346 11734
rect 130082 10218 130138 10220
rect 130082 10166 130084 10218
rect 130084 10166 130136 10218
rect 130136 10166 130138 10218
rect 130082 10164 130138 10166
rect 130186 10218 130242 10220
rect 130186 10166 130188 10218
rect 130188 10166 130240 10218
rect 130240 10166 130242 10218
rect 130186 10164 130242 10166
rect 130290 10218 130346 10220
rect 130290 10166 130292 10218
rect 130292 10166 130344 10218
rect 130344 10166 130346 10218
rect 130290 10164 130346 10166
rect 130082 8650 130138 8652
rect 130082 8598 130084 8650
rect 130084 8598 130136 8650
rect 130136 8598 130138 8650
rect 130082 8596 130138 8598
rect 130186 8650 130242 8652
rect 130186 8598 130188 8650
rect 130188 8598 130240 8650
rect 130240 8598 130242 8650
rect 130186 8596 130242 8598
rect 130290 8650 130346 8652
rect 130290 8598 130292 8650
rect 130292 8598 130344 8650
rect 130344 8598 130346 8650
rect 130290 8596 130346 8598
rect 126812 8034 126868 8036
rect 126812 7982 126814 8034
rect 126814 7982 126866 8034
rect 126866 7982 126868 8034
rect 126812 7980 126868 7982
rect 127260 7868 127316 7924
rect 126812 7698 126868 7700
rect 126812 7646 126814 7698
rect 126814 7646 126866 7698
rect 126866 7646 126868 7698
rect 126812 7644 126868 7646
rect 126588 6412 126644 6468
rect 127260 7084 127316 7140
rect 127260 6130 127316 6132
rect 127260 6078 127262 6130
rect 127262 6078 127314 6130
rect 127314 6078 127316 6130
rect 127260 6076 127316 6078
rect 127484 6076 127540 6132
rect 126700 5516 126756 5572
rect 127372 5516 127428 5572
rect 127260 5180 127316 5236
rect 130082 7082 130138 7084
rect 130082 7030 130084 7082
rect 130084 7030 130136 7082
rect 130136 7030 130138 7082
rect 130082 7028 130138 7030
rect 130186 7082 130242 7084
rect 130186 7030 130188 7082
rect 130188 7030 130240 7082
rect 130240 7030 130242 7082
rect 130186 7028 130242 7030
rect 130290 7082 130346 7084
rect 130290 7030 130292 7082
rect 130292 7030 130344 7082
rect 130344 7030 130346 7082
rect 130290 7028 130346 7030
rect 128044 5964 128100 6020
rect 128380 6412 128436 6468
rect 127596 5740 127652 5796
rect 127932 5682 127988 5684
rect 127932 5630 127934 5682
rect 127934 5630 127986 5682
rect 127986 5630 127988 5682
rect 127932 5628 127988 5630
rect 128044 5516 128100 5572
rect 128044 4956 128100 5012
rect 128604 6300 128660 6356
rect 129388 6466 129444 6468
rect 129388 6414 129390 6466
rect 129390 6414 129442 6466
rect 129442 6414 129444 6466
rect 129388 6412 129444 6414
rect 129388 6130 129444 6132
rect 129388 6078 129390 6130
rect 129390 6078 129442 6130
rect 129442 6078 129444 6130
rect 129388 6076 129444 6078
rect 127484 4620 127540 4676
rect 127260 3778 127316 3780
rect 127260 3726 127262 3778
rect 127262 3726 127314 3778
rect 127314 3726 127316 3778
rect 127260 3724 127316 3726
rect 128156 4620 128212 4676
rect 128044 4562 128100 4564
rect 128044 4510 128046 4562
rect 128046 4510 128098 4562
rect 128098 4510 128100 4562
rect 128044 4508 128100 4510
rect 127484 4450 127540 4452
rect 127484 4398 127486 4450
rect 127486 4398 127538 4450
rect 127538 4398 127540 4450
rect 127484 4396 127540 4398
rect 129052 5516 129108 5572
rect 128380 4284 128436 4340
rect 128940 4338 128996 4340
rect 128940 4286 128942 4338
rect 128942 4286 128994 4338
rect 128994 4286 128996 4338
rect 128940 4284 128996 4286
rect 129276 3948 129332 4004
rect 129388 5068 129444 5124
rect 129500 4396 129556 4452
rect 129500 3724 129556 3780
rect 128044 3388 128100 3444
rect 128604 3442 128660 3444
rect 128604 3390 128606 3442
rect 128606 3390 128658 3442
rect 128658 3390 128660 3442
rect 128604 3388 128660 3390
rect 130082 5514 130138 5516
rect 130082 5462 130084 5514
rect 130084 5462 130136 5514
rect 130136 5462 130138 5514
rect 130082 5460 130138 5462
rect 130186 5514 130242 5516
rect 130186 5462 130188 5514
rect 130188 5462 130240 5514
rect 130240 5462 130242 5514
rect 130186 5460 130242 5462
rect 130290 5514 130346 5516
rect 130290 5462 130292 5514
rect 130292 5462 130344 5514
rect 130344 5462 130346 5514
rect 130290 5460 130346 5462
rect 130284 5068 130340 5124
rect 129948 4732 130004 4788
rect 130082 3946 130138 3948
rect 130082 3894 130084 3946
rect 130084 3894 130136 3946
rect 130136 3894 130138 3946
rect 130082 3892 130138 3894
rect 130186 3946 130242 3948
rect 130186 3894 130188 3946
rect 130188 3894 130240 3946
rect 130240 3894 130242 3946
rect 130186 3892 130242 3894
rect 130290 3946 130346 3948
rect 130290 3894 130292 3946
rect 130292 3894 130344 3946
rect 130344 3894 130346 3946
rect 130290 3892 130346 3894
rect 131068 34860 131124 34916
rect 131404 35532 131460 35588
rect 131628 35586 131684 35588
rect 131628 35534 131630 35586
rect 131630 35534 131682 35586
rect 131682 35534 131684 35586
rect 131628 35532 131684 35534
rect 131740 35420 131796 35476
rect 131292 34860 131348 34916
rect 131516 35196 131572 35252
rect 130844 34076 130900 34132
rect 131180 34242 131236 34244
rect 131180 34190 131182 34242
rect 131182 34190 131234 34242
rect 131234 34190 131236 34242
rect 131180 34188 131236 34190
rect 130620 32956 130676 33012
rect 130844 5964 130900 6020
rect 132076 35644 132132 35700
rect 132524 35756 132580 35812
rect 132076 35196 132132 35252
rect 131964 34914 132020 34916
rect 131964 34862 131966 34914
rect 131966 34862 132018 34914
rect 132018 34862 132020 34914
rect 131964 34860 132020 34862
rect 132188 6300 132244 6356
rect 131852 5292 131908 5348
rect 131964 5740 132020 5796
rect 130956 4620 131012 4676
rect 132076 5180 132132 5236
rect 133756 36876 133812 36932
rect 133644 35756 133700 35812
rect 132972 35644 133028 35700
rect 132748 34860 132804 34916
rect 132636 34636 132692 34692
rect 135212 38108 135268 38164
rect 134988 36258 135044 36260
rect 134988 36206 134990 36258
rect 134990 36206 135042 36258
rect 135042 36206 135044 36258
rect 134988 36204 135044 36206
rect 134764 35810 134820 35812
rect 134764 35758 134766 35810
rect 134766 35758 134818 35810
rect 134818 35758 134820 35810
rect 134764 35756 134820 35758
rect 134540 35644 134596 35700
rect 133868 35084 133924 35140
rect 133196 34914 133252 34916
rect 133196 34862 133198 34914
rect 133198 34862 133250 34914
rect 133250 34862 133252 34914
rect 133196 34860 133252 34862
rect 133756 34690 133812 34692
rect 133756 34638 133758 34690
rect 133758 34638 133810 34690
rect 133810 34638 133812 34690
rect 133756 34636 133812 34638
rect 132412 6076 132468 6132
rect 133532 33852 133588 33908
rect 132188 5516 132244 5572
rect 133196 5906 133252 5908
rect 133196 5854 133198 5906
rect 133198 5854 133250 5906
rect 133250 5854 133252 5906
rect 133196 5852 133252 5854
rect 132972 5628 133028 5684
rect 132300 5180 132356 5236
rect 131628 3724 131684 3780
rect 133420 5346 133476 5348
rect 133420 5294 133422 5346
rect 133422 5294 133474 5346
rect 133474 5294 133476 5346
rect 133420 5292 133476 5294
rect 132300 3724 132356 3780
rect 133084 5122 133140 5124
rect 133084 5070 133086 5122
rect 133086 5070 133138 5122
rect 133138 5070 133140 5122
rect 133084 5068 133140 5070
rect 133308 4844 133364 4900
rect 132972 4226 133028 4228
rect 132972 4174 132974 4226
rect 132974 4174 133026 4226
rect 133026 4174 133028 4226
rect 132972 4172 133028 4174
rect 134092 33852 134148 33908
rect 134764 34524 134820 34580
rect 135772 38108 135828 38164
rect 135436 35084 135492 35140
rect 135548 36316 135604 36372
rect 136332 36428 136388 36484
rect 136220 36370 136276 36372
rect 136220 36318 136222 36370
rect 136222 36318 136274 36370
rect 136274 36318 136276 36370
rect 136220 36316 136276 36318
rect 136556 36092 136612 36148
rect 136220 35980 136276 36036
rect 137116 35980 137172 36036
rect 135884 35698 135940 35700
rect 135884 35646 135886 35698
rect 135886 35646 135938 35698
rect 135938 35646 135940 35698
rect 135884 35644 135940 35646
rect 136892 35698 136948 35700
rect 136892 35646 136894 35698
rect 136894 35646 136946 35698
rect 136946 35646 136948 35698
rect 136892 35644 136948 35646
rect 135660 35532 135716 35588
rect 136332 35084 136388 35140
rect 134428 33852 134484 33908
rect 137116 34636 137172 34692
rect 135772 33180 135828 33236
rect 135996 33964 136052 34020
rect 135996 30156 136052 30212
rect 136780 8876 136836 8932
rect 135660 7868 135716 7924
rect 135772 7196 135828 7252
rect 137116 7980 137172 8036
rect 136780 6690 136836 6692
rect 136780 6638 136782 6690
rect 136782 6638 136834 6690
rect 136834 6638 136836 6690
rect 136780 6636 136836 6638
rect 135996 6578 136052 6580
rect 135996 6526 135998 6578
rect 135998 6526 136050 6578
rect 136050 6526 136052 6578
rect 135996 6524 136052 6526
rect 135772 6188 135828 6244
rect 134204 6130 134260 6132
rect 134204 6078 134206 6130
rect 134206 6078 134258 6130
rect 134258 6078 134260 6130
rect 134204 6076 134260 6078
rect 133756 5852 133812 5908
rect 134652 5628 134708 5684
rect 135212 5740 135268 5796
rect 133756 5180 133812 5236
rect 133980 5516 134036 5572
rect 134204 5180 134260 5236
rect 134764 5234 134820 5236
rect 134764 5182 134766 5234
rect 134766 5182 134818 5234
rect 134818 5182 134820 5234
rect 134764 5180 134820 5182
rect 135772 5010 135828 5012
rect 135772 4958 135774 5010
rect 135774 4958 135826 5010
rect 135826 4958 135828 5010
rect 135772 4956 135828 4958
rect 133308 4172 133364 4228
rect 132636 3612 132692 3668
rect 131068 3554 131124 3556
rect 131068 3502 131070 3554
rect 131070 3502 131122 3554
rect 131122 3502 131124 3554
rect 131068 3500 131124 3502
rect 133868 4172 133924 4228
rect 132076 3388 132132 3444
rect 132636 3442 132692 3444
rect 132636 3390 132638 3442
rect 132638 3390 132690 3442
rect 132690 3390 132692 3442
rect 132636 3388 132692 3390
rect 134428 4226 134484 4228
rect 134428 4174 134430 4226
rect 134430 4174 134482 4226
rect 134482 4174 134484 4226
rect 134428 4172 134484 4174
rect 137004 5404 137060 5460
rect 135996 4844 136052 4900
rect 137340 36204 137396 36260
rect 137788 36482 137844 36484
rect 137788 36430 137790 36482
rect 137790 36430 137842 36482
rect 137842 36430 137844 36482
rect 137788 36428 137844 36430
rect 137564 36092 137620 36148
rect 137900 35922 137956 35924
rect 137900 35870 137902 35922
rect 137902 35870 137954 35922
rect 137954 35870 137956 35922
rect 137900 35868 137956 35870
rect 139020 36652 139076 36708
rect 140588 38668 140644 38724
rect 138572 35980 138628 36036
rect 137452 35196 137508 35252
rect 138124 35196 138180 35252
rect 137452 34300 137508 34356
rect 139916 35868 139972 35924
rect 139356 35474 139412 35476
rect 139356 35422 139358 35474
rect 139358 35422 139410 35474
rect 139410 35422 139412 35474
rect 139356 35420 139412 35422
rect 139132 34636 139188 34692
rect 138908 33964 138964 34020
rect 138012 31836 138068 31892
rect 137564 7644 137620 7700
rect 139132 7698 139188 7700
rect 139132 7646 139134 7698
rect 139134 7646 139186 7698
rect 139186 7646 139188 7698
rect 139132 7644 139188 7646
rect 139804 35420 139860 35476
rect 140028 34300 140084 34356
rect 139692 7644 139748 7700
rect 139916 7756 139972 7812
rect 138124 6636 138180 6692
rect 137788 6578 137844 6580
rect 137788 6526 137790 6578
rect 137790 6526 137842 6578
rect 137842 6526 137844 6578
rect 137788 6524 137844 6526
rect 137340 6076 137396 6132
rect 137452 6188 137508 6244
rect 137228 5292 137284 5348
rect 137452 5068 137508 5124
rect 137900 5852 137956 5908
rect 137788 5404 137844 5460
rect 137788 5180 137844 5236
rect 138124 5852 138180 5908
rect 138460 6524 138516 6580
rect 138236 5180 138292 5236
rect 139356 6802 139412 6804
rect 139356 6750 139358 6802
rect 139358 6750 139410 6802
rect 139410 6750 139412 6802
rect 139356 6748 139412 6750
rect 138572 6130 138628 6132
rect 138572 6078 138574 6130
rect 138574 6078 138626 6130
rect 138626 6078 138628 6130
rect 138572 6076 138628 6078
rect 139132 6578 139188 6580
rect 139132 6526 139134 6578
rect 139134 6526 139186 6578
rect 139186 6526 139188 6578
rect 139132 6524 139188 6526
rect 138684 5516 138740 5572
rect 139020 5852 139076 5908
rect 138460 5404 138516 5460
rect 138796 5292 138852 5348
rect 138348 4562 138404 4564
rect 138348 4510 138350 4562
rect 138350 4510 138402 4562
rect 138402 4510 138404 4562
rect 138348 4508 138404 4510
rect 139580 5906 139636 5908
rect 139580 5854 139582 5906
rect 139582 5854 139634 5906
rect 139634 5854 139636 5906
rect 139580 5852 139636 5854
rect 139468 5234 139524 5236
rect 139468 5182 139470 5234
rect 139470 5182 139522 5234
rect 139522 5182 139524 5234
rect 139468 5180 139524 5182
rect 139804 5964 139860 6020
rect 139692 5068 139748 5124
rect 136108 3388 136164 3444
rect 136668 3442 136724 3444
rect 136668 3390 136670 3442
rect 136670 3390 136722 3442
rect 136722 3390 136724 3442
rect 136668 3388 136724 3390
rect 137452 3388 137508 3444
rect 140476 35980 140532 36036
rect 140812 36540 140868 36596
rect 140924 36988 140980 37044
rect 140364 34354 140420 34356
rect 140364 34302 140366 34354
rect 140366 34302 140418 34354
rect 140418 34302 140420 34354
rect 140364 34300 140420 34302
rect 141596 36652 141652 36708
rect 142156 35980 142212 36036
rect 142604 35868 142660 35924
rect 141260 35586 141316 35588
rect 141260 35534 141262 35586
rect 141262 35534 141314 35586
rect 141314 35534 141316 35586
rect 141260 35532 141316 35534
rect 141260 35308 141316 35364
rect 141036 34524 141092 34580
rect 140252 6748 140308 6804
rect 140812 6748 140868 6804
rect 140140 6018 140196 6020
rect 140140 5966 140142 6018
rect 140142 5966 140194 6018
rect 140194 5966 140196 6018
rect 140140 5964 140196 5966
rect 140700 6018 140756 6020
rect 140700 5966 140702 6018
rect 140702 5966 140754 6018
rect 140754 5966 140756 6018
rect 140700 5964 140756 5966
rect 141932 35532 141988 35588
rect 141484 34188 141540 34244
rect 141260 6524 141316 6580
rect 142156 34802 142212 34804
rect 142156 34750 142158 34802
rect 142158 34750 142210 34802
rect 142210 34750 142212 34802
rect 142156 34748 142212 34750
rect 142940 35308 142996 35364
rect 143612 36594 143668 36596
rect 143612 36542 143614 36594
rect 143614 36542 143666 36594
rect 143666 36542 143668 36594
rect 143612 36540 143668 36542
rect 144396 36540 144452 36596
rect 143724 35868 143780 35924
rect 145852 37548 145908 37604
rect 145404 36594 145460 36596
rect 145404 36542 145406 36594
rect 145406 36542 145458 36594
rect 145458 36542 145460 36594
rect 145404 36540 145460 36542
rect 145292 35868 145348 35924
rect 148492 36090 148548 36092
rect 148492 36038 148494 36090
rect 148494 36038 148546 36090
rect 148546 36038 148548 36090
rect 148492 36036 148548 36038
rect 148596 36090 148652 36092
rect 148596 36038 148598 36090
rect 148598 36038 148650 36090
rect 148650 36038 148652 36090
rect 148596 36036 148652 36038
rect 148700 36090 148756 36092
rect 148700 36038 148702 36090
rect 148702 36038 148754 36090
rect 148754 36038 148756 36090
rect 148700 36036 148756 36038
rect 146188 35868 146244 35924
rect 146636 35922 146692 35924
rect 146636 35870 146638 35922
rect 146638 35870 146690 35922
rect 146690 35870 146692 35922
rect 146636 35868 146692 35870
rect 145180 34972 145236 35028
rect 145516 35026 145572 35028
rect 145516 34974 145518 35026
rect 145518 34974 145570 35026
rect 145570 34974 145572 35026
rect 145516 34972 145572 34974
rect 143500 34860 143556 34916
rect 142940 34802 142996 34804
rect 142940 34750 142942 34802
rect 142942 34750 142994 34802
rect 142994 34750 142996 34802
rect 142940 34748 142996 34750
rect 143948 34914 144004 34916
rect 143948 34862 143950 34914
rect 143950 34862 144002 34914
rect 144002 34862 144004 34914
rect 143948 34860 144004 34862
rect 142268 34242 142324 34244
rect 142268 34190 142270 34242
rect 142270 34190 142322 34242
rect 142322 34190 142324 34242
rect 142268 34188 142324 34190
rect 141596 5180 141652 5236
rect 140924 4508 140980 4564
rect 148492 34522 148548 34524
rect 148492 34470 148494 34522
rect 148494 34470 148546 34522
rect 148546 34470 148548 34522
rect 148492 34468 148548 34470
rect 148596 34522 148652 34524
rect 148596 34470 148598 34522
rect 148598 34470 148650 34522
rect 148650 34470 148652 34522
rect 148596 34468 148652 34470
rect 148700 34522 148756 34524
rect 148700 34470 148702 34522
rect 148702 34470 148754 34522
rect 148754 34470 148756 34522
rect 148700 34468 148756 34470
rect 148492 32954 148548 32956
rect 148492 32902 148494 32954
rect 148494 32902 148546 32954
rect 148546 32902 148548 32954
rect 148492 32900 148548 32902
rect 148596 32954 148652 32956
rect 148596 32902 148598 32954
rect 148598 32902 148650 32954
rect 148650 32902 148652 32954
rect 148596 32900 148652 32902
rect 148700 32954 148756 32956
rect 148700 32902 148702 32954
rect 148702 32902 148754 32954
rect 148754 32902 148756 32954
rect 148700 32900 148756 32902
rect 143724 31724 143780 31780
rect 143948 6860 144004 6916
rect 138012 3388 138068 3444
rect 140140 3388 140196 3444
rect 141260 3442 141316 3444
rect 141260 3390 141262 3442
rect 141262 3390 141314 3442
rect 141314 3390 141316 3442
rect 141260 3388 141316 3390
rect 148492 31386 148548 31388
rect 148492 31334 148494 31386
rect 148494 31334 148546 31386
rect 148546 31334 148548 31386
rect 148492 31332 148548 31334
rect 148596 31386 148652 31388
rect 148596 31334 148598 31386
rect 148598 31334 148650 31386
rect 148650 31334 148652 31386
rect 148596 31332 148652 31334
rect 148700 31386 148756 31388
rect 148700 31334 148702 31386
rect 148702 31334 148754 31386
rect 148754 31334 148756 31386
rect 148700 31332 148756 31334
rect 148492 29818 148548 29820
rect 148492 29766 148494 29818
rect 148494 29766 148546 29818
rect 148546 29766 148548 29818
rect 148492 29764 148548 29766
rect 148596 29818 148652 29820
rect 148596 29766 148598 29818
rect 148598 29766 148650 29818
rect 148650 29766 148652 29818
rect 148596 29764 148652 29766
rect 148700 29818 148756 29820
rect 148700 29766 148702 29818
rect 148702 29766 148754 29818
rect 148754 29766 148756 29818
rect 148700 29764 148756 29766
rect 148492 28250 148548 28252
rect 148492 28198 148494 28250
rect 148494 28198 148546 28250
rect 148546 28198 148548 28250
rect 148492 28196 148548 28198
rect 148596 28250 148652 28252
rect 148596 28198 148598 28250
rect 148598 28198 148650 28250
rect 148650 28198 148652 28250
rect 148596 28196 148652 28198
rect 148700 28250 148756 28252
rect 148700 28198 148702 28250
rect 148702 28198 148754 28250
rect 148754 28198 148756 28250
rect 148700 28196 148756 28198
rect 148492 26682 148548 26684
rect 148492 26630 148494 26682
rect 148494 26630 148546 26682
rect 148546 26630 148548 26682
rect 148492 26628 148548 26630
rect 148596 26682 148652 26684
rect 148596 26630 148598 26682
rect 148598 26630 148650 26682
rect 148650 26630 148652 26682
rect 148596 26628 148652 26630
rect 148700 26682 148756 26684
rect 148700 26630 148702 26682
rect 148702 26630 148754 26682
rect 148754 26630 148756 26682
rect 148700 26628 148756 26630
rect 148492 25114 148548 25116
rect 148492 25062 148494 25114
rect 148494 25062 148546 25114
rect 148546 25062 148548 25114
rect 148492 25060 148548 25062
rect 148596 25114 148652 25116
rect 148596 25062 148598 25114
rect 148598 25062 148650 25114
rect 148650 25062 148652 25114
rect 148596 25060 148652 25062
rect 148700 25114 148756 25116
rect 148700 25062 148702 25114
rect 148702 25062 148754 25114
rect 148754 25062 148756 25114
rect 148700 25060 148756 25062
rect 148492 23546 148548 23548
rect 148492 23494 148494 23546
rect 148494 23494 148546 23546
rect 148546 23494 148548 23546
rect 148492 23492 148548 23494
rect 148596 23546 148652 23548
rect 148596 23494 148598 23546
rect 148598 23494 148650 23546
rect 148650 23494 148652 23546
rect 148596 23492 148652 23494
rect 148700 23546 148756 23548
rect 148700 23494 148702 23546
rect 148702 23494 148754 23546
rect 148754 23494 148756 23546
rect 148700 23492 148756 23494
rect 148492 21978 148548 21980
rect 148492 21926 148494 21978
rect 148494 21926 148546 21978
rect 148546 21926 148548 21978
rect 148492 21924 148548 21926
rect 148596 21978 148652 21980
rect 148596 21926 148598 21978
rect 148598 21926 148650 21978
rect 148650 21926 148652 21978
rect 148596 21924 148652 21926
rect 148700 21978 148756 21980
rect 148700 21926 148702 21978
rect 148702 21926 148754 21978
rect 148754 21926 148756 21978
rect 148700 21924 148756 21926
rect 148492 20410 148548 20412
rect 148492 20358 148494 20410
rect 148494 20358 148546 20410
rect 148546 20358 148548 20410
rect 148492 20356 148548 20358
rect 148596 20410 148652 20412
rect 148596 20358 148598 20410
rect 148598 20358 148650 20410
rect 148650 20358 148652 20410
rect 148596 20356 148652 20358
rect 148700 20410 148756 20412
rect 148700 20358 148702 20410
rect 148702 20358 148754 20410
rect 148754 20358 148756 20410
rect 148700 20356 148756 20358
rect 148492 18842 148548 18844
rect 148492 18790 148494 18842
rect 148494 18790 148546 18842
rect 148546 18790 148548 18842
rect 148492 18788 148548 18790
rect 148596 18842 148652 18844
rect 148596 18790 148598 18842
rect 148598 18790 148650 18842
rect 148650 18790 148652 18842
rect 148596 18788 148652 18790
rect 148700 18842 148756 18844
rect 148700 18790 148702 18842
rect 148702 18790 148754 18842
rect 148754 18790 148756 18842
rect 148700 18788 148756 18790
rect 148492 17274 148548 17276
rect 148492 17222 148494 17274
rect 148494 17222 148546 17274
rect 148546 17222 148548 17274
rect 148492 17220 148548 17222
rect 148596 17274 148652 17276
rect 148596 17222 148598 17274
rect 148598 17222 148650 17274
rect 148650 17222 148652 17274
rect 148596 17220 148652 17222
rect 148700 17274 148756 17276
rect 148700 17222 148702 17274
rect 148702 17222 148754 17274
rect 148754 17222 148756 17274
rect 148700 17220 148756 17222
rect 148492 15706 148548 15708
rect 148492 15654 148494 15706
rect 148494 15654 148546 15706
rect 148546 15654 148548 15706
rect 148492 15652 148548 15654
rect 148596 15706 148652 15708
rect 148596 15654 148598 15706
rect 148598 15654 148650 15706
rect 148650 15654 148652 15706
rect 148596 15652 148652 15654
rect 148700 15706 148756 15708
rect 148700 15654 148702 15706
rect 148702 15654 148754 15706
rect 148754 15654 148756 15706
rect 148700 15652 148756 15654
rect 148492 14138 148548 14140
rect 148492 14086 148494 14138
rect 148494 14086 148546 14138
rect 148546 14086 148548 14138
rect 148492 14084 148548 14086
rect 148596 14138 148652 14140
rect 148596 14086 148598 14138
rect 148598 14086 148650 14138
rect 148650 14086 148652 14138
rect 148596 14084 148652 14086
rect 148700 14138 148756 14140
rect 148700 14086 148702 14138
rect 148702 14086 148754 14138
rect 148754 14086 148756 14138
rect 148700 14084 148756 14086
rect 148492 12570 148548 12572
rect 148492 12518 148494 12570
rect 148494 12518 148546 12570
rect 148546 12518 148548 12570
rect 148492 12516 148548 12518
rect 148596 12570 148652 12572
rect 148596 12518 148598 12570
rect 148598 12518 148650 12570
rect 148650 12518 148652 12570
rect 148596 12516 148652 12518
rect 148700 12570 148756 12572
rect 148700 12518 148702 12570
rect 148702 12518 148754 12570
rect 148754 12518 148756 12570
rect 148700 12516 148756 12518
rect 148492 11002 148548 11004
rect 148492 10950 148494 11002
rect 148494 10950 148546 11002
rect 148546 10950 148548 11002
rect 148492 10948 148548 10950
rect 148596 11002 148652 11004
rect 148596 10950 148598 11002
rect 148598 10950 148650 11002
rect 148650 10950 148652 11002
rect 148596 10948 148652 10950
rect 148700 11002 148756 11004
rect 148700 10950 148702 11002
rect 148702 10950 148754 11002
rect 148754 10950 148756 11002
rect 148700 10948 148756 10950
rect 148492 9434 148548 9436
rect 148492 9382 148494 9434
rect 148494 9382 148546 9434
rect 148546 9382 148548 9434
rect 148492 9380 148548 9382
rect 148596 9434 148652 9436
rect 148596 9382 148598 9434
rect 148598 9382 148650 9434
rect 148650 9382 148652 9434
rect 148596 9380 148652 9382
rect 148700 9434 148756 9436
rect 148700 9382 148702 9434
rect 148702 9382 148754 9434
rect 148754 9382 148756 9434
rect 148700 9380 148756 9382
rect 148492 7866 148548 7868
rect 148492 7814 148494 7866
rect 148494 7814 148546 7866
rect 148546 7814 148548 7866
rect 148492 7812 148548 7814
rect 148596 7866 148652 7868
rect 148596 7814 148598 7866
rect 148598 7814 148650 7866
rect 148650 7814 148652 7866
rect 148596 7812 148652 7814
rect 148700 7866 148756 7868
rect 148700 7814 148702 7866
rect 148702 7814 148754 7866
rect 148754 7814 148756 7866
rect 148700 7812 148756 7814
rect 148492 6298 148548 6300
rect 148492 6246 148494 6298
rect 148494 6246 148546 6298
rect 148546 6246 148548 6298
rect 148492 6244 148548 6246
rect 148596 6298 148652 6300
rect 148596 6246 148598 6298
rect 148598 6246 148650 6298
rect 148650 6246 148652 6298
rect 148596 6244 148652 6246
rect 148700 6298 148756 6300
rect 148700 6246 148702 6298
rect 148702 6246 148754 6298
rect 148754 6246 148756 6298
rect 148700 6244 148756 6246
rect 148492 4730 148548 4732
rect 148492 4678 148494 4730
rect 148494 4678 148546 4730
rect 148546 4678 148548 4730
rect 148492 4676 148548 4678
rect 148596 4730 148652 4732
rect 148596 4678 148598 4730
rect 148598 4678 148650 4730
rect 148650 4678 148652 4730
rect 148596 4676 148652 4678
rect 148700 4730 148756 4732
rect 148700 4678 148702 4730
rect 148702 4678 148754 4730
rect 148754 4678 148756 4730
rect 148700 4676 148756 4678
rect 144172 3388 144228 3444
rect 145292 3442 145348 3444
rect 145292 3390 145294 3442
rect 145294 3390 145346 3442
rect 145346 3390 145348 3442
rect 145292 3388 145348 3390
rect 148492 3162 148548 3164
rect 148492 3110 148494 3162
rect 148494 3110 148546 3162
rect 148546 3110 148548 3162
rect 148492 3108 148548 3110
rect 148596 3162 148652 3164
rect 148596 3110 148598 3162
rect 148598 3110 148650 3162
rect 148650 3110 148652 3162
rect 148596 3108 148652 3110
rect 148700 3162 148756 3164
rect 148700 3110 148702 3162
rect 148702 3110 148754 3162
rect 148754 3110 148756 3162
rect 148700 3108 148756 3110
<< metal3 >>
rect 80322 38780 80332 38836
rect 80388 38780 111132 38836
rect 111188 38780 111198 38836
rect 72818 38668 72828 38724
rect 72884 38668 140588 38724
rect 140644 38668 140654 38724
rect 58930 38556 58940 38612
rect 58996 38556 123116 38612
rect 123172 38556 123182 38612
rect 23090 38444 23100 38500
rect 23156 38444 82012 38500
rect 82068 38444 82078 38500
rect 38994 38332 39004 38388
rect 39060 38332 88172 38388
rect 88228 38332 88238 38388
rect 56914 38220 56924 38276
rect 56980 38220 92316 38276
rect 92372 38220 92382 38276
rect 65650 38108 65660 38164
rect 65716 38108 135212 38164
rect 135268 38108 135772 38164
rect 135828 38108 135838 38164
rect 57138 37996 57148 38052
rect 57204 37996 103740 38052
rect 103796 37996 103806 38052
rect 61394 37884 61404 37940
rect 61460 37884 110236 37940
rect 110292 37884 110302 37940
rect 30146 37772 30156 37828
rect 30212 37772 68796 37828
rect 68852 37772 68862 37828
rect 69682 37772 69692 37828
rect 69748 37772 118748 37828
rect 118804 37772 118814 37828
rect 60722 37660 60732 37716
rect 60788 37660 113148 37716
rect 113204 37660 113214 37716
rect 26562 37548 26572 37604
rect 26628 37548 80556 37604
rect 80612 37548 80622 37604
rect 89058 37548 89068 37604
rect 89124 37548 145852 37604
rect 145908 37548 145918 37604
rect 64306 37436 64316 37492
rect 64372 37436 121548 37492
rect 121604 37436 121614 37492
rect 15810 37324 15820 37380
rect 15876 37324 59612 37380
rect 59668 37324 59678 37380
rect 62626 37324 62636 37380
rect 62692 37324 86940 37380
rect 86996 37324 87006 37380
rect 28354 37212 28364 37268
rect 28420 37212 49308 37268
rect 49364 37212 52892 37268
rect 52948 37212 52958 37268
rect 64642 37212 64652 37268
rect 64708 37212 130844 37268
rect 130900 37212 130910 37268
rect 8866 37100 8876 37156
rect 8932 37100 72492 37156
rect 72548 37100 73836 37156
rect 73892 37100 73902 37156
rect 87266 37100 87276 37156
rect 87332 37100 103516 37156
rect 103572 37100 104188 37156
rect 104244 37100 104254 37156
rect 33842 36988 33852 37044
rect 33908 36988 62524 37044
rect 62580 36988 62590 37044
rect 102162 36988 102172 37044
rect 102228 36988 140924 37044
rect 140980 36988 140990 37044
rect 45714 36876 45724 36932
rect 45780 36876 47628 36932
rect 47684 36876 47694 36932
rect 68226 36876 68236 36932
rect 68292 36876 68908 36932
rect 68964 36876 68974 36932
rect 70018 36876 70028 36932
rect 70084 36876 70588 36932
rect 70644 36876 70654 36932
rect 75058 36876 75068 36932
rect 75124 36876 89068 36932
rect 89124 36876 89134 36932
rect 97234 36876 97244 36932
rect 97300 36876 97468 36932
rect 131842 36876 131852 36932
rect 131908 36876 133756 36932
rect 133812 36876 133822 36932
rect 19612 36820 19622 36876
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19886 36820 19896 36876
rect 56432 36820 56442 36876
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56706 36820 56716 36876
rect 93252 36820 93262 36876
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93526 36820 93536 36876
rect 97412 36820 97468 36876
rect 130072 36820 130082 36876
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130346 36820 130356 36876
rect 25778 36764 25788 36820
rect 25844 36764 41804 36820
rect 41860 36764 41870 36820
rect 61282 36764 61292 36820
rect 61348 36764 74396 36820
rect 74452 36764 74620 36820
rect 74676 36764 74686 36820
rect 78082 36764 78092 36820
rect 78148 36764 80892 36820
rect 80948 36764 80958 36820
rect 83458 36764 83468 36820
rect 83524 36764 84812 36820
rect 84868 36764 84878 36820
rect 85250 36764 85260 36820
rect 85316 36764 86156 36820
rect 86212 36764 86222 36820
rect 97412 36764 121100 36820
rect 121156 36764 121166 36820
rect 30146 36652 30156 36708
rect 30212 36652 31724 36708
rect 31780 36652 31790 36708
rect 46722 36652 46732 36708
rect 46788 36652 47628 36708
rect 47684 36652 47694 36708
rect 52658 36652 52668 36708
rect 52724 36652 53900 36708
rect 53956 36652 101052 36708
rect 101108 36652 101118 36708
rect 110338 36652 110348 36708
rect 110404 36652 112252 36708
rect 112308 36652 112318 36708
rect 139010 36652 139020 36708
rect 139076 36652 141596 36708
rect 141652 36652 141662 36708
rect 16034 36540 16044 36596
rect 16100 36540 17164 36596
rect 17220 36540 17230 36596
rect 21634 36540 21644 36596
rect 21700 36540 22204 36596
rect 22260 36540 22270 36596
rect 27794 36540 27804 36596
rect 27860 36540 28812 36596
rect 28868 36540 28878 36596
rect 33506 36540 33516 36596
rect 33572 36540 35084 36596
rect 35140 36540 36092 36596
rect 36148 36540 36158 36596
rect 48514 36540 48524 36596
rect 48580 36540 49532 36596
rect 49588 36540 49598 36596
rect 51314 36540 51324 36596
rect 51380 36540 52108 36596
rect 52164 36540 52174 36596
rect 64530 36540 64540 36596
rect 64596 36540 66108 36596
rect 66164 36540 66174 36596
rect 66434 36540 66444 36596
rect 66500 36540 67900 36596
rect 67956 36540 67966 36596
rect 68786 36540 68796 36596
rect 68852 36540 91980 36596
rect 92036 36540 92046 36596
rect 94210 36540 94220 36596
rect 94276 36540 96572 36596
rect 96628 36540 96638 36596
rect 96898 36540 96908 36596
rect 96964 36540 98364 36596
rect 98420 36540 98430 36596
rect 100482 36540 100492 36596
rect 100548 36540 102396 36596
rect 102452 36540 102462 36596
rect 103170 36540 103180 36596
rect 103236 36540 104412 36596
rect 104468 36540 104478 36596
rect 112130 36540 112140 36596
rect 112196 36540 114044 36596
rect 114100 36540 114110 36596
rect 115714 36540 115724 36596
rect 115780 36540 116620 36596
rect 116676 36540 116686 36596
rect 122882 36540 122892 36596
rect 122948 36540 126028 36596
rect 126084 36540 126094 36596
rect 126466 36540 126476 36596
rect 126532 36540 127932 36596
rect 127988 36540 127998 36596
rect 128258 36540 128268 36596
rect 128324 36540 129724 36596
rect 129780 36540 129790 36596
rect 140802 36540 140812 36596
rect 140868 36540 143612 36596
rect 143668 36540 143678 36596
rect 144386 36540 144396 36596
rect 144452 36540 145404 36596
rect 145460 36540 145470 36596
rect 8978 36428 8988 36484
rect 9044 36428 9772 36484
rect 9828 36428 9838 36484
rect 28466 36428 28476 36484
rect 28532 36428 29596 36484
rect 29652 36428 29662 36484
rect 31826 36428 31836 36484
rect 31892 36428 32172 36484
rect 32228 36428 32238 36484
rect 38434 36428 38444 36484
rect 38500 36428 39116 36484
rect 39172 36428 39182 36484
rect 40226 36428 40236 36484
rect 40292 36428 40908 36484
rect 40964 36428 40974 36484
rect 43362 36428 43372 36484
rect 43428 36428 44156 36484
rect 44212 36428 57596 36484
rect 57652 36428 57662 36484
rect 58818 36428 58828 36484
rect 58884 36428 59164 36484
rect 59220 36428 61404 36484
rect 61460 36428 61470 36484
rect 64978 36428 64988 36484
rect 65044 36428 65548 36484
rect 65604 36428 65614 36484
rect 66770 36428 66780 36484
rect 66836 36428 67676 36484
rect 67732 36428 67742 36484
rect 86930 36428 86940 36484
rect 86996 36428 87948 36484
rect 88004 36428 88014 36484
rect 88946 36428 88956 36484
rect 89012 36428 92820 36484
rect 92978 36428 92988 36484
rect 93044 36428 103348 36484
rect 106194 36428 106204 36484
rect 106260 36428 108668 36484
rect 108724 36428 108734 36484
rect 109330 36428 109340 36484
rect 109396 36428 110124 36484
rect 110180 36428 110190 36484
rect 118066 36428 118076 36484
rect 118132 36428 119532 36484
rect 119588 36428 119598 36484
rect 136322 36428 136332 36484
rect 136388 36428 137788 36484
rect 137844 36428 137854 36484
rect 17490 36316 17500 36372
rect 17556 36316 18172 36372
rect 18228 36316 19516 36372
rect 19572 36316 20188 36372
rect 20244 36316 20254 36372
rect 43250 36316 43260 36372
rect 43316 36316 45724 36372
rect 45780 36316 45790 36372
rect 65314 36316 65324 36372
rect 65380 36316 65660 36372
rect 65716 36316 65726 36372
rect 67778 36316 67788 36372
rect 67844 36316 69692 36372
rect 69748 36316 69758 36372
rect 78754 36316 78764 36372
rect 78820 36316 79436 36372
rect 79492 36316 79502 36372
rect 90692 36316 91196 36372
rect 91252 36316 91262 36372
rect 90692 36260 90748 36316
rect 92764 36260 92820 36428
rect 94322 36316 94332 36372
rect 94388 36316 95900 36372
rect 95956 36316 95966 36372
rect 103292 36260 103348 36428
rect 106418 36316 106428 36372
rect 106484 36316 107212 36372
rect 107268 36316 122444 36372
rect 122500 36316 122510 36372
rect 129602 36316 129612 36372
rect 129668 36316 135548 36372
rect 135604 36316 136220 36372
rect 136276 36316 136286 36372
rect 137340 36260 137396 36428
rect 45266 36204 45276 36260
rect 45332 36204 47516 36260
rect 47572 36204 55468 36260
rect 58706 36204 58716 36260
rect 58772 36204 59500 36260
rect 59556 36204 59566 36260
rect 72594 36204 72604 36260
rect 72660 36204 78428 36260
rect 78484 36204 78494 36260
rect 89506 36204 89516 36260
rect 89572 36204 89740 36260
rect 89796 36204 90748 36260
rect 92754 36204 92764 36260
rect 92820 36204 103236 36260
rect 103292 36204 116844 36260
rect 116900 36204 116910 36260
rect 117618 36204 117628 36260
rect 117684 36204 123452 36260
rect 123508 36204 123518 36260
rect 128146 36204 128156 36260
rect 128212 36204 131292 36260
rect 131348 36204 134988 36260
rect 135044 36204 135054 36260
rect 137330 36204 137340 36260
rect 137396 36204 137406 36260
rect 55412 36148 55468 36204
rect 19730 36092 19740 36148
rect 19796 36092 24220 36148
rect 24276 36092 24286 36148
rect 51986 36092 51996 36148
rect 52052 36092 54572 36148
rect 54628 36092 54638 36148
rect 55412 36092 68572 36148
rect 68628 36092 68638 36148
rect 70802 36092 70812 36148
rect 70868 36092 72828 36148
rect 72884 36092 72894 36148
rect 73714 36092 73724 36148
rect 73780 36092 74508 36148
rect 74564 36092 74574 36148
rect 84812 36092 93100 36148
rect 93156 36092 93772 36148
rect 93828 36092 93838 36148
rect 38022 36036 38032 36092
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38296 36036 38306 36092
rect 74842 36036 74852 36092
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 75116 36036 75126 36092
rect 10882 35980 10892 36036
rect 10948 35980 11788 36036
rect 11844 35980 11854 36036
rect 31892 35980 37940 36036
rect 46050 35980 46060 36036
rect 46116 35980 73108 36036
rect 77522 35980 77532 36036
rect 77588 35980 80332 36036
rect 80388 35980 80398 36036
rect 31892 35924 31948 35980
rect 37884 35924 37940 35980
rect 73052 35924 73108 35980
rect 84812 35924 84868 36092
rect 103180 36036 103236 36204
rect 108658 36092 108668 36148
rect 108724 36092 109228 36148
rect 109284 36092 109294 36148
rect 136546 36092 136556 36148
rect 136612 36092 137564 36148
rect 137620 36092 137630 36148
rect 111662 36036 111672 36092
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111936 36036 111946 36092
rect 148482 36036 148492 36092
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148756 36036 148766 36092
rect 90626 35980 90636 36036
rect 90692 35980 91868 36036
rect 91924 35980 91934 36036
rect 92306 35980 92316 36036
rect 92372 35980 100604 36036
rect 100660 35980 100670 36036
rect 103180 35980 109228 36036
rect 136210 35980 136220 36036
rect 136276 35980 137116 36036
rect 137172 35980 138572 36036
rect 138628 35980 140476 36036
rect 140532 35980 142156 36036
rect 142212 35980 142222 36036
rect 6066 35868 6076 35924
rect 6132 35868 6972 35924
rect 7028 35868 31948 35924
rect 32172 35868 36316 35924
rect 36372 35868 36382 35924
rect 37884 35868 42588 35924
rect 42644 35868 42654 35924
rect 53778 35868 53788 35924
rect 53844 35868 54796 35924
rect 54852 35868 72996 35924
rect 73052 35868 84868 35924
rect 87612 35868 99820 35924
rect 99876 35868 99886 35924
rect 32172 35812 32228 35868
rect 72940 35812 72996 35868
rect 6402 35756 6412 35812
rect 6468 35756 7532 35812
rect 7588 35756 7598 35812
rect 13234 35756 13244 35812
rect 13300 35756 13804 35812
rect 13860 35756 13870 35812
rect 20402 35756 20412 35812
rect 20468 35756 32228 35812
rect 32386 35756 32396 35812
rect 32452 35756 34524 35812
rect 34580 35756 34590 35812
rect 39890 35756 39900 35812
rect 39956 35756 41132 35812
rect 41188 35756 41198 35812
rect 41794 35756 41804 35812
rect 41860 35756 43932 35812
rect 43988 35756 43998 35812
rect 46386 35756 46396 35812
rect 46452 35756 46956 35812
rect 47012 35756 47022 35812
rect 58594 35756 58604 35812
rect 58660 35756 59276 35812
rect 59332 35756 60172 35812
rect 60228 35756 60238 35812
rect 70466 35756 70476 35812
rect 70532 35756 70924 35812
rect 70980 35756 70990 35812
rect 72940 35756 83300 35812
rect 83458 35756 83468 35812
rect 83524 35756 87388 35812
rect 87444 35756 87454 35812
rect 83244 35700 83300 35756
rect 87612 35700 87668 35868
rect 89954 35756 89964 35812
rect 90020 35756 93548 35812
rect 93604 35756 93614 35812
rect 101042 35756 101052 35812
rect 101108 35756 101612 35812
rect 101668 35756 101678 35812
rect 102274 35756 102284 35812
rect 102340 35756 102844 35812
rect 102900 35756 102910 35812
rect 103730 35756 103740 35812
rect 103796 35756 106316 35812
rect 106372 35756 107548 35812
rect 107604 35756 107614 35812
rect 109172 35700 109228 35980
rect 111346 35868 111356 35924
rect 111412 35868 113372 35924
rect 113428 35868 113438 35924
rect 119858 35868 119868 35924
rect 119924 35868 121324 35924
rect 121380 35868 121390 35924
rect 122322 35868 122332 35924
rect 122388 35868 125244 35924
rect 125300 35868 125310 35924
rect 137890 35868 137900 35924
rect 137956 35868 139916 35924
rect 139972 35868 139982 35924
rect 142594 35868 142604 35924
rect 142660 35868 143724 35924
rect 143780 35868 143790 35924
rect 145282 35868 145292 35924
rect 145348 35868 146188 35924
rect 146244 35868 146636 35924
rect 146692 35868 146702 35924
rect 112242 35756 112252 35812
rect 112308 35756 114268 35812
rect 114324 35756 114334 35812
rect 116274 35756 116284 35812
rect 116340 35756 117740 35812
rect 117796 35756 117806 35812
rect 123106 35756 123116 35812
rect 123172 35756 124124 35812
rect 124180 35756 124460 35812
rect 124516 35756 124526 35812
rect 124674 35756 124684 35812
rect 124740 35756 126252 35812
rect 126308 35756 126318 35812
rect 130834 35756 130844 35812
rect 130900 35756 132524 35812
rect 132580 35756 132590 35812
rect 133634 35756 133644 35812
rect 133700 35756 134764 35812
rect 134820 35756 134830 35812
rect 12002 35644 12012 35700
rect 12068 35644 18956 35700
rect 19012 35644 19022 35700
rect 29362 35644 29372 35700
rect 29428 35644 32620 35700
rect 32676 35644 32686 35700
rect 54898 35644 54908 35700
rect 54964 35644 55244 35700
rect 55300 35644 55310 35700
rect 56690 35644 56700 35700
rect 56756 35644 57484 35700
rect 57540 35644 57550 35700
rect 66098 35644 66108 35700
rect 66164 35644 66668 35700
rect 66724 35644 66734 35700
rect 69906 35644 69916 35700
rect 69972 35644 78540 35700
rect 78596 35644 78606 35700
rect 78754 35644 78764 35700
rect 78820 35644 79100 35700
rect 79156 35644 79166 35700
rect 80546 35644 80556 35700
rect 80612 35644 81340 35700
rect 81396 35644 81406 35700
rect 83244 35644 87668 35700
rect 90178 35644 90188 35700
rect 90244 35644 92988 35700
rect 93044 35644 93054 35700
rect 94322 35644 94332 35700
rect 94388 35644 97244 35700
rect 97300 35644 97310 35700
rect 109172 35644 113092 35700
rect 113474 35644 113484 35700
rect 113540 35644 115500 35700
rect 115556 35644 115566 35700
rect 123666 35644 123676 35700
rect 123732 35644 125356 35700
rect 125412 35644 125422 35700
rect 127922 35644 127932 35700
rect 127988 35644 129052 35700
rect 129108 35644 130060 35700
rect 130116 35644 131292 35700
rect 131348 35644 131358 35700
rect 132066 35644 132076 35700
rect 132132 35644 132972 35700
rect 133028 35644 133038 35700
rect 134530 35644 134540 35700
rect 134596 35644 135884 35700
rect 135940 35644 136892 35700
rect 136948 35644 136958 35700
rect 8754 35532 8764 35588
rect 8820 35532 9660 35588
rect 9716 35532 20188 35588
rect 23426 35532 23436 35588
rect 23492 35532 24332 35588
rect 24388 35532 24398 35588
rect 29698 35532 29708 35588
rect 29764 35532 31500 35588
rect 31556 35532 31566 35588
rect 37538 35532 37548 35588
rect 37604 35532 38108 35588
rect 38164 35532 39340 35588
rect 39396 35532 39564 35588
rect 39620 35532 39630 35588
rect 45602 35532 45612 35588
rect 45668 35532 46172 35588
rect 46228 35532 46238 35588
rect 53778 35532 53788 35588
rect 53844 35532 54236 35588
rect 54292 35532 61292 35588
rect 61348 35532 61358 35588
rect 74274 35532 74284 35588
rect 74340 35532 74620 35588
rect 74676 35532 75852 35588
rect 75908 35532 75918 35588
rect 77186 35532 77196 35588
rect 77252 35532 79212 35588
rect 79268 35532 79278 35588
rect 80770 35532 80780 35588
rect 80836 35532 82012 35588
rect 82068 35532 82078 35588
rect 87042 35532 87052 35588
rect 87108 35532 87948 35588
rect 88004 35532 88014 35588
rect 106530 35532 106540 35588
rect 106596 35532 107324 35588
rect 107380 35532 107390 35588
rect 20132 35476 20188 35532
rect 113036 35476 113092 35644
rect 113922 35532 113932 35588
rect 113988 35532 114828 35588
rect 114884 35532 114894 35588
rect 117506 35532 117516 35588
rect 117572 35532 118412 35588
rect 118468 35532 118478 35588
rect 121986 35532 121996 35588
rect 122052 35532 122780 35588
rect 122836 35532 122846 35588
rect 124562 35532 124572 35588
rect 124628 35532 127372 35588
rect 127428 35532 131404 35588
rect 131460 35532 131470 35588
rect 131618 35532 131628 35588
rect 131684 35532 135660 35588
rect 135716 35532 135726 35588
rect 141250 35532 141260 35588
rect 141316 35532 141932 35588
rect 141988 35532 141998 35588
rect 18274 35420 18284 35476
rect 18340 35420 19404 35476
rect 19460 35420 19470 35476
rect 20132 35420 25676 35476
rect 25732 35420 25900 35476
rect 25956 35420 26236 35476
rect 26292 35420 26302 35476
rect 40786 35420 40796 35476
rect 40852 35420 44380 35476
rect 44436 35420 44446 35476
rect 52994 35420 53004 35476
rect 53060 35420 53676 35476
rect 53732 35420 53742 35476
rect 66546 35420 66556 35476
rect 66612 35420 67452 35476
rect 67508 35420 67518 35476
rect 75394 35420 75404 35476
rect 75460 35420 76748 35476
rect 76804 35420 76814 35476
rect 90402 35420 90412 35476
rect 90468 35420 90972 35476
rect 91028 35420 91038 35476
rect 105522 35420 105532 35476
rect 105588 35420 109228 35476
rect 109284 35420 109294 35476
rect 110338 35420 110348 35476
rect 110404 35420 112812 35476
rect 112868 35420 112878 35476
rect 113036 35420 115052 35476
rect 115108 35420 115118 35476
rect 119522 35420 119532 35476
rect 119588 35420 123564 35476
rect 123620 35420 123630 35476
rect 123890 35420 123900 35476
rect 123956 35420 125132 35476
rect 125188 35420 131740 35476
rect 131796 35420 131806 35476
rect 139346 35420 139356 35476
rect 139412 35420 139804 35476
rect 139860 35420 139870 35476
rect 20066 35308 20076 35364
rect 20132 35308 20748 35364
rect 20804 35308 20814 35364
rect 20972 35308 22092 35364
rect 22148 35308 22158 35364
rect 23986 35308 23996 35364
rect 24052 35308 51660 35364
rect 51716 35308 51726 35364
rect 73266 35308 73276 35364
rect 73332 35308 74732 35364
rect 74788 35308 74798 35364
rect 108322 35308 108332 35364
rect 108388 35308 127260 35364
rect 127316 35308 127326 35364
rect 141250 35308 141260 35364
rect 141316 35308 142940 35364
rect 142996 35308 143006 35364
rect 19612 35252 19622 35308
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19886 35252 19896 35308
rect 20132 35252 20188 35308
rect 20972 35252 21028 35308
rect 56432 35252 56442 35308
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56706 35252 56716 35308
rect 93252 35252 93262 35308
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93526 35252 93536 35308
rect 130072 35252 130082 35308
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130346 35252 130356 35308
rect 20132 35196 21028 35252
rect 23090 35196 23100 35252
rect 23156 35196 37772 35252
rect 37828 35196 37838 35252
rect 43652 35196 49196 35252
rect 49252 35196 49532 35252
rect 49588 35196 49598 35252
rect 61394 35196 61404 35252
rect 61460 35196 69580 35252
rect 69636 35196 70140 35252
rect 70196 35196 70206 35252
rect 71586 35196 71596 35252
rect 71652 35196 78204 35252
rect 78260 35196 78270 35252
rect 79874 35196 79884 35252
rect 79940 35196 82684 35252
rect 82740 35196 82750 35252
rect 93874 35196 93884 35252
rect 93940 35196 95564 35252
rect 95620 35196 95630 35252
rect 98802 35196 98812 35252
rect 98868 35196 99596 35252
rect 99652 35196 100044 35252
rect 100100 35196 100110 35252
rect 107314 35196 107324 35252
rect 107380 35196 111468 35252
rect 111524 35196 111534 35252
rect 131058 35196 131068 35252
rect 131124 35196 131516 35252
rect 131572 35196 132076 35252
rect 132132 35196 132142 35252
rect 137442 35196 137452 35252
rect 137508 35196 138124 35252
rect 138180 35196 138190 35252
rect 20132 35140 20188 35196
rect 43652 35140 43708 35196
rect 7858 35084 7868 35140
rect 7924 35084 8876 35140
rect 8932 35084 8942 35140
rect 9090 35084 9100 35140
rect 9156 35084 10108 35140
rect 10164 35084 10174 35140
rect 13580 35084 20188 35140
rect 30594 35084 30604 35140
rect 30660 35084 31388 35140
rect 31444 35084 43708 35140
rect 45042 35084 45052 35140
rect 45108 35084 45724 35140
rect 45780 35084 45790 35140
rect 49970 35084 49980 35140
rect 50036 35084 78092 35140
rect 78148 35084 78158 35140
rect 78418 35084 78428 35140
rect 78484 35084 85540 35140
rect 88050 35084 88060 35140
rect 88116 35084 88844 35140
rect 88900 35084 88910 35140
rect 89618 35084 89628 35140
rect 89684 35084 91868 35140
rect 91924 35084 91934 35140
rect 95106 35084 95116 35140
rect 95172 35084 96012 35140
rect 96068 35084 96078 35140
rect 106978 35084 106988 35140
rect 107044 35084 108780 35140
rect 108836 35084 108846 35140
rect 108994 35084 109004 35140
rect 109060 35084 109788 35140
rect 109844 35084 109854 35140
rect 113026 35084 113036 35140
rect 113092 35084 114380 35140
rect 114436 35084 114446 35140
rect 115490 35084 115500 35140
rect 115556 35084 117516 35140
rect 117572 35084 117852 35140
rect 117908 35084 117918 35140
rect 118626 35084 118636 35140
rect 118692 35084 119868 35140
rect 119924 35084 120428 35140
rect 120484 35084 120494 35140
rect 128034 35084 128044 35140
rect 128100 35084 133868 35140
rect 133924 35084 133934 35140
rect 135426 35084 135436 35140
rect 135492 35084 136332 35140
rect 136388 35084 136398 35140
rect 10322 34972 10332 35028
rect 10388 34972 11004 35028
rect 11060 34972 11070 35028
rect 13580 34916 13636 35084
rect 13804 34972 61292 35028
rect 61348 34972 61358 35028
rect 62850 34972 62860 35028
rect 62916 34972 63420 35028
rect 63476 34972 63486 35028
rect 66658 34972 66668 35028
rect 66724 34972 68516 35028
rect 68674 34972 68684 35028
rect 68740 34972 69132 35028
rect 69188 34972 69198 35028
rect 72034 34972 72044 35028
rect 72100 34972 72716 35028
rect 72772 34972 72782 35028
rect 76290 34972 76300 35028
rect 76356 34972 77980 35028
rect 78036 34972 78046 35028
rect 78306 34972 78316 35028
rect 78372 34972 78988 35028
rect 81666 34972 81676 35028
rect 81732 34972 82572 35028
rect 82628 34972 82638 35028
rect 6178 34860 6188 34916
rect 6244 34860 6972 34916
rect 7028 34860 8428 34916
rect 12898 34860 12908 34916
rect 12964 34860 13580 34916
rect 13636 34860 13646 34916
rect 8372 34804 8428 34860
rect 13804 34804 13860 34972
rect 68460 34916 68516 34972
rect 78932 34916 78988 34972
rect 14578 34860 14588 34916
rect 14644 34860 14812 34916
rect 14868 34860 15820 34916
rect 15876 34860 15886 34916
rect 19282 34860 19292 34916
rect 19348 34860 20300 34916
rect 20356 34860 20366 34916
rect 27916 34860 29372 34916
rect 29428 34860 29438 34916
rect 29922 34860 29932 34916
rect 29988 34860 31948 34916
rect 32834 34860 32844 34916
rect 32900 34860 33292 34916
rect 33348 34860 33358 34916
rect 37762 34860 37772 34916
rect 37828 34860 38332 34916
rect 38388 34860 38398 34916
rect 54562 34860 54572 34916
rect 54628 34860 55020 34916
rect 55076 34860 55086 34916
rect 56018 34860 56028 34916
rect 56084 34860 57372 34916
rect 57428 34860 57438 34916
rect 59602 34860 59612 34916
rect 59668 34860 62188 34916
rect 62244 34860 62254 34916
rect 67106 34860 67116 34916
rect 67172 34860 67340 34916
rect 67396 34860 67564 34916
rect 67620 34860 67630 34916
rect 68460 34860 74732 34916
rect 74788 34860 74798 34916
rect 75282 34860 75292 34916
rect 75348 34860 75628 34916
rect 75684 34860 75694 34916
rect 76178 34860 76188 34916
rect 76244 34860 77308 34916
rect 77364 34860 77374 34916
rect 78932 34860 85260 34916
rect 85316 34860 85326 34916
rect 27916 34804 27972 34860
rect 31892 34804 31948 34860
rect 85484 34804 85540 35084
rect 88722 34972 88732 35028
rect 88788 34972 90188 35028
rect 90244 34972 90254 35028
rect 92418 34972 92428 35028
rect 92484 34972 93996 35028
rect 94052 34972 94062 35028
rect 96114 34972 96124 35028
rect 96180 34972 97356 35028
rect 97412 34972 97422 35028
rect 104962 34972 104972 35028
rect 105028 34972 105868 35028
rect 105924 34972 105934 35028
rect 107314 34972 107324 35028
rect 107380 34972 145180 35028
rect 145236 34972 145516 35028
rect 145572 34972 145582 35028
rect 85698 34860 85708 34916
rect 85764 34860 96628 34916
rect 8372 34748 11116 34804
rect 11172 34748 13860 34804
rect 19506 34748 19516 34804
rect 19572 34748 27972 34804
rect 28130 34748 28140 34804
rect 28196 34748 28700 34804
rect 28756 34748 28766 34804
rect 31892 34748 56476 34804
rect 56532 34748 56542 34804
rect 63858 34748 63868 34804
rect 63924 34748 74396 34804
rect 74452 34748 75404 34804
rect 75460 34748 75470 34804
rect 85484 34748 90748 34804
rect 90692 34692 90748 34748
rect 96572 34692 96628 34860
rect 97412 34860 120988 34916
rect 122098 34860 122108 34916
rect 122164 34860 122668 34916
rect 122724 34860 122734 34916
rect 124002 34860 124012 34916
rect 124068 34860 124796 34916
rect 124852 34860 125244 34916
rect 125300 34860 125310 34916
rect 125570 34860 125580 34916
rect 125636 34860 126588 34916
rect 126644 34860 127036 34916
rect 127092 34860 127102 34916
rect 127474 34860 127484 34916
rect 127540 34860 128828 34916
rect 128884 34860 129388 34916
rect 129444 34860 129454 34916
rect 129938 34860 129948 34916
rect 130004 34860 131068 34916
rect 131124 34860 131134 34916
rect 131282 34860 131292 34916
rect 131348 34860 131964 34916
rect 132020 34860 132030 34916
rect 132738 34860 132748 34916
rect 132804 34860 133196 34916
rect 133252 34860 133262 34916
rect 143490 34860 143500 34916
rect 143556 34860 143948 34916
rect 144004 34860 144014 34916
rect 97412 34692 97468 34860
rect 120932 34804 120988 34860
rect 103282 34748 103292 34804
rect 103348 34748 106988 34804
rect 107044 34748 107054 34804
rect 107202 34748 107212 34804
rect 107268 34748 107278 34804
rect 114370 34748 114380 34804
rect 114436 34748 115836 34804
rect 115892 34748 115902 34804
rect 120932 34748 142156 34804
rect 142212 34748 142940 34804
rect 142996 34748 143006 34804
rect 15474 34636 15484 34692
rect 15540 34636 29036 34692
rect 29092 34636 30156 34692
rect 30212 34636 30222 34692
rect 37762 34636 37772 34692
rect 37828 34636 46844 34692
rect 46900 34636 46910 34692
rect 48066 34636 48076 34692
rect 48132 34636 50316 34692
rect 50372 34636 50382 34692
rect 74722 34636 74732 34692
rect 74788 34636 76636 34692
rect 76692 34636 78764 34692
rect 78820 34636 78830 34692
rect 79426 34636 79436 34692
rect 79492 34636 80668 34692
rect 80724 34636 85708 34692
rect 85764 34636 85774 34692
rect 90692 34636 93324 34692
rect 93380 34636 96236 34692
rect 96292 34636 96302 34692
rect 96572 34636 97468 34692
rect 99922 34636 99932 34692
rect 99988 34636 101612 34692
rect 101668 34636 102956 34692
rect 103012 34636 103022 34692
rect 107212 34580 107268 34748
rect 22866 34524 22876 34580
rect 22932 34524 22942 34580
rect 54002 34524 54012 34580
rect 54068 34524 73164 34580
rect 73220 34524 73836 34580
rect 73892 34524 73902 34580
rect 75394 34524 75404 34580
rect 75460 34524 87388 34580
rect 87444 34524 87948 34580
rect 88004 34524 89292 34580
rect 89348 34524 89358 34580
rect 92418 34524 92428 34580
rect 92484 34524 93436 34580
rect 93492 34524 107268 34580
rect 107324 34636 108556 34692
rect 108612 34636 110796 34692
rect 110852 34636 110862 34692
rect 111244 34636 111580 34692
rect 111636 34636 111646 34692
rect 113474 34636 113484 34692
rect 113540 34636 115948 34692
rect 116004 34636 116014 34692
rect 121874 34636 121884 34692
rect 121940 34636 122108 34692
rect 122164 34636 127708 34692
rect 127764 34636 127774 34692
rect 132626 34636 132636 34692
rect 132692 34636 133756 34692
rect 133812 34636 133822 34692
rect 137106 34636 137116 34692
rect 137172 34636 139132 34692
rect 139188 34636 139198 34692
rect 22876 34468 22932 34524
rect 38022 34468 38032 34524
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38296 34468 38306 34524
rect 74842 34468 74852 34524
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 75116 34468 75126 34524
rect 107324 34468 107380 34636
rect 111244 34580 111300 34636
rect 111234 34524 111244 34580
rect 111300 34524 111310 34580
rect 111662 34468 111672 34524
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111936 34468 111946 34524
rect 132692 34468 132748 34636
rect 134754 34524 134764 34580
rect 134820 34524 141036 34580
rect 141092 34524 141102 34580
rect 148482 34468 148492 34524
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148756 34468 148766 34524
rect 8530 34412 8540 34468
rect 8596 34412 8876 34468
rect 8932 34412 9660 34468
rect 9716 34412 23324 34468
rect 23380 34412 23390 34468
rect 42578 34412 42588 34468
rect 42644 34412 52220 34468
rect 52276 34412 52286 34468
rect 56018 34412 56028 34468
rect 56084 34412 65436 34468
rect 65492 34412 65772 34468
rect 65828 34412 65838 34468
rect 84018 34412 84028 34468
rect 84084 34412 84588 34468
rect 84644 34412 97468 34468
rect 105522 34412 105532 34468
rect 105588 34412 107380 34468
rect 109218 34412 109228 34468
rect 109284 34412 109452 34468
rect 109508 34412 109900 34468
rect 109956 34412 109966 34468
rect 118066 34412 118076 34468
rect 118132 34412 132748 34468
rect 97412 34356 97468 34412
rect 10994 34300 11004 34356
rect 11060 34300 20076 34356
rect 20132 34300 20142 34356
rect 25442 34300 25452 34356
rect 25508 34300 26012 34356
rect 26068 34300 26078 34356
rect 28690 34300 28700 34356
rect 28756 34300 47068 34356
rect 47124 34300 47292 34356
rect 47348 34300 47740 34356
rect 47796 34300 47806 34356
rect 48850 34300 48860 34356
rect 48916 34300 49644 34356
rect 49700 34300 49710 34356
rect 50978 34300 50988 34356
rect 51044 34300 60116 34356
rect 62626 34300 62636 34356
rect 62692 34300 63084 34356
rect 63140 34300 63868 34356
rect 63924 34300 63934 34356
rect 73938 34300 73948 34356
rect 74004 34300 75964 34356
rect 76020 34300 76030 34356
rect 77410 34300 77420 34356
rect 77476 34300 78204 34356
rect 78260 34300 78270 34356
rect 78754 34300 78764 34356
rect 78820 34300 78988 34356
rect 79044 34300 79436 34356
rect 79492 34300 79502 34356
rect 91522 34300 91532 34356
rect 91588 34300 92652 34356
rect 92708 34300 92718 34356
rect 97412 34300 123004 34356
rect 123060 34300 123340 34356
rect 123396 34300 123406 34356
rect 130274 34300 130284 34356
rect 130340 34300 137452 34356
rect 137508 34300 137518 34356
rect 140018 34300 140028 34356
rect 140084 34300 140364 34356
rect 140420 34300 140430 34356
rect 60060 34244 60116 34300
rect 8754 34188 8764 34244
rect 8820 34188 17500 34244
rect 17556 34188 17836 34244
rect 17892 34188 17902 34244
rect 20402 34188 20412 34244
rect 20468 34188 25004 34244
rect 25060 34188 25070 34244
rect 46050 34188 46060 34244
rect 46116 34188 48524 34244
rect 48580 34188 48590 34244
rect 51650 34188 51660 34244
rect 51716 34188 53116 34244
rect 53172 34188 53182 34244
rect 53442 34188 53452 34244
rect 53508 34188 56028 34244
rect 56084 34188 56094 34244
rect 60060 34188 64764 34244
rect 64820 34188 64830 34244
rect 74162 34188 74172 34244
rect 74228 34188 80444 34244
rect 80500 34188 80510 34244
rect 82338 34188 82348 34244
rect 82404 34188 83132 34244
rect 83188 34188 83198 34244
rect 86034 34188 86044 34244
rect 86100 34188 102172 34244
rect 102228 34188 102238 34244
rect 105634 34188 105644 34244
rect 105700 34188 106428 34244
rect 106484 34188 106494 34244
rect 109172 34188 114044 34244
rect 114100 34188 114110 34244
rect 129154 34188 129164 34244
rect 129220 34188 131180 34244
rect 131236 34188 131246 34244
rect 141474 34188 141484 34244
rect 141540 34188 142268 34244
rect 142324 34188 142334 34244
rect 109172 34132 109228 34188
rect 24882 34076 24892 34132
rect 24948 34076 25564 34132
rect 25620 34076 37548 34132
rect 37604 34076 37614 34132
rect 44706 34076 44716 34132
rect 44772 34076 47180 34132
rect 47236 34076 48188 34132
rect 48244 34076 60060 34132
rect 60116 34076 60126 34132
rect 60610 34076 60620 34132
rect 60676 34076 61180 34132
rect 61236 34076 62300 34132
rect 62356 34076 62366 34132
rect 66322 34076 66332 34132
rect 66388 34076 67004 34132
rect 67060 34076 67070 34132
rect 78194 34076 78204 34132
rect 78260 34076 109228 34132
rect 123778 34076 123788 34132
rect 123844 34076 125580 34132
rect 125636 34076 130844 34132
rect 130900 34076 130910 34132
rect 13010 33964 13020 34020
rect 13076 33964 13468 34020
rect 13524 33964 34524 34020
rect 34580 33964 35084 34020
rect 35140 33964 35150 34020
rect 43586 33964 43596 34020
rect 43652 33964 44492 34020
rect 44548 33964 45276 34020
rect 45332 33964 45342 34020
rect 46946 33964 46956 34020
rect 47012 33964 47404 34020
rect 47460 33964 48412 34020
rect 48468 33964 48478 34020
rect 51202 33964 51212 34020
rect 51268 33964 52332 34020
rect 52388 33964 52398 34020
rect 56130 33964 56140 34020
rect 56196 33964 56476 34020
rect 56532 33964 59052 34020
rect 59108 33964 59118 34020
rect 59826 33964 59836 34020
rect 59892 33964 60172 34020
rect 60228 33964 60238 34020
rect 72146 33964 72156 34020
rect 72212 33964 76860 34020
rect 76916 33964 77196 34020
rect 77252 33964 77262 34020
rect 90290 33964 90300 34020
rect 90356 33964 90636 34020
rect 90692 33964 90702 34020
rect 123554 33964 123564 34020
rect 123620 33964 124348 34020
rect 124404 33964 124414 34020
rect 126466 33964 126476 34020
rect 126532 33964 126924 34020
rect 126980 33964 130060 34020
rect 130116 33964 130126 34020
rect 135986 33964 135996 34020
rect 136052 33964 138908 34020
rect 138964 33964 138974 34020
rect 21298 33852 21308 33908
rect 21364 33852 21756 33908
rect 21812 33852 40684 33908
rect 40740 33852 41916 33908
rect 41972 33852 41982 33908
rect 52098 33852 52108 33908
rect 52164 33852 56028 33908
rect 56084 33852 56094 33908
rect 56252 33852 56588 33908
rect 56644 33852 56654 33908
rect 78932 33852 95452 33908
rect 95508 33852 95518 33908
rect 108770 33852 108780 33908
rect 108836 33852 125020 33908
rect 125076 33852 125086 33908
rect 126812 33852 133532 33908
rect 133588 33852 134092 33908
rect 134148 33852 134428 33908
rect 134484 33852 134494 33908
rect 22418 33740 22428 33796
rect 22484 33740 37436 33796
rect 37492 33740 38556 33796
rect 38612 33740 39116 33796
rect 39172 33740 39182 33796
rect 19612 33684 19622 33740
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19886 33684 19896 33740
rect 56252 33684 56308 33852
rect 78932 33796 78988 33852
rect 126812 33796 126868 33852
rect 68562 33740 68572 33796
rect 68628 33740 78988 33796
rect 100706 33740 100716 33796
rect 100772 33740 104300 33796
rect 104356 33740 104366 33796
rect 113922 33740 113932 33796
rect 113988 33740 114380 33796
rect 114436 33740 118076 33796
rect 118132 33740 118142 33796
rect 119298 33740 119308 33796
rect 119364 33740 126868 33796
rect 56432 33684 56442 33740
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56706 33684 56716 33740
rect 93252 33684 93262 33740
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93526 33684 93536 33740
rect 130072 33684 130082 33740
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130346 33684 130356 33740
rect 20066 33628 20076 33684
rect 20132 33628 20636 33684
rect 20692 33628 21756 33684
rect 21812 33628 21822 33684
rect 34178 33628 34188 33684
rect 34244 33628 56252 33684
rect 56308 33628 56318 33684
rect 61394 33628 61404 33684
rect 61460 33628 63532 33684
rect 63588 33628 63598 33684
rect 89394 33628 89404 33684
rect 89460 33628 90524 33684
rect 90580 33628 90590 33684
rect 102498 33628 102508 33684
rect 102564 33628 106092 33684
rect 106148 33628 106158 33684
rect 18610 33516 18620 33572
rect 18676 33516 19852 33572
rect 19908 33516 19918 33572
rect 27122 33516 27132 33572
rect 27188 33516 50652 33572
rect 50708 33516 51212 33572
rect 51268 33516 51278 33572
rect 55794 33516 55804 33572
rect 55860 33516 83692 33572
rect 83748 33516 83758 33572
rect 88498 33516 88508 33572
rect 88564 33516 105756 33572
rect 105812 33516 106204 33572
rect 106260 33516 108332 33572
rect 108388 33516 109452 33572
rect 109508 33516 109518 33572
rect 111010 33516 111020 33572
rect 111076 33516 112252 33572
rect 112308 33516 112318 33572
rect 126466 33516 126476 33572
rect 126532 33516 127372 33572
rect 127428 33516 128716 33572
rect 128772 33516 129276 33572
rect 129332 33516 129342 33572
rect 18386 33404 18396 33460
rect 18452 33404 19292 33460
rect 19348 33404 19358 33460
rect 30034 33404 30044 33460
rect 30100 33404 30604 33460
rect 30660 33404 31052 33460
rect 31108 33404 44716 33460
rect 44772 33404 44782 33460
rect 45826 33404 45836 33460
rect 45892 33404 46284 33460
rect 46340 33404 46350 33460
rect 53330 33404 53340 33460
rect 53396 33404 54012 33460
rect 54068 33404 54078 33460
rect 60274 33404 60284 33460
rect 60340 33404 60732 33460
rect 60788 33404 60798 33460
rect 61730 33404 61740 33460
rect 61796 33404 61964 33460
rect 62020 33404 62030 33460
rect 63410 33404 63420 33460
rect 63476 33404 65100 33460
rect 65156 33404 67228 33460
rect 72706 33404 72716 33460
rect 72772 33404 92092 33460
rect 92148 33404 92158 33460
rect 110002 33404 110012 33460
rect 110068 33404 110796 33460
rect 110852 33404 128604 33460
rect 128660 33404 128670 33460
rect 67172 33348 67228 33404
rect 31154 33292 31164 33348
rect 31220 33292 51548 33348
rect 51604 33292 51614 33348
rect 52434 33292 52444 33348
rect 52500 33292 52780 33348
rect 52836 33292 54460 33348
rect 54516 33292 61292 33348
rect 61348 33292 62748 33348
rect 62804 33292 63308 33348
rect 63364 33292 63756 33348
rect 63812 33292 63822 33348
rect 67172 33292 102508 33348
rect 102564 33292 102574 33348
rect 110114 33292 110124 33348
rect 110180 33292 126812 33348
rect 126868 33292 126878 33348
rect 17042 33180 17052 33236
rect 17108 33180 37772 33236
rect 37828 33180 38332 33236
rect 38388 33180 38668 33236
rect 38724 33180 38734 33236
rect 48514 33180 48524 33236
rect 48580 33180 89516 33236
rect 89572 33180 89582 33236
rect 96002 33180 96012 33236
rect 96068 33180 119644 33236
rect 119700 33180 119710 33236
rect 129602 33180 129612 33236
rect 129668 33180 135772 33236
rect 135828 33180 135838 33236
rect 19842 33068 19852 33124
rect 19908 33068 28364 33124
rect 28420 33068 28430 33124
rect 37986 33068 37996 33124
rect 38052 33068 43148 33124
rect 43204 33068 43214 33124
rect 62066 33068 62076 33124
rect 62132 33068 62412 33124
rect 62468 33068 62478 33124
rect 102610 33068 102620 33124
rect 102676 33068 106876 33124
rect 106932 33068 107996 33124
rect 108052 33068 108062 33124
rect 110898 33068 110908 33124
rect 110964 33068 128268 33124
rect 128324 33068 129052 33124
rect 129108 33068 129118 33124
rect 118178 32956 118188 33012
rect 118244 32956 130172 33012
rect 130228 32956 130620 33012
rect 130676 32956 130686 33012
rect 38022 32900 38032 32956
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38296 32900 38306 32956
rect 74842 32900 74852 32956
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 75116 32900 75126 32956
rect 111662 32900 111672 32956
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111936 32900 111946 32956
rect 148482 32900 148492 32956
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148756 32900 148766 32956
rect 38546 32844 38556 32900
rect 38612 32844 65884 32900
rect 65940 32844 65950 32900
rect 18274 32732 18284 32788
rect 18340 32732 58716 32788
rect 58772 32732 58782 32788
rect 61618 32732 61628 32788
rect 61684 32732 62972 32788
rect 63028 32732 63038 32788
rect 63186 32732 63196 32788
rect 63252 32732 64204 32788
rect 64260 32732 100716 32788
rect 100772 32732 100782 32788
rect 101602 32732 101612 32788
rect 101668 32732 111020 32788
rect 111076 32732 111086 32788
rect 43026 32620 43036 32676
rect 43092 32620 76076 32676
rect 76132 32620 76142 32676
rect 79762 32620 79772 32676
rect 79828 32620 105196 32676
rect 105252 32620 105262 32676
rect 36754 32508 36764 32564
rect 36820 32508 52108 32564
rect 52164 32508 52174 32564
rect 67442 32508 67452 32564
rect 67508 32508 107548 32564
rect 107604 32508 107614 32564
rect 20290 32396 20300 32452
rect 20356 32396 60284 32452
rect 60340 32396 61852 32452
rect 61908 32396 61918 32452
rect 40338 32284 40348 32340
rect 40404 32284 72156 32340
rect 72212 32284 72222 32340
rect 19612 32116 19622 32172
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19886 32116 19896 32172
rect 56432 32116 56442 32172
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56706 32116 56716 32172
rect 93252 32116 93262 32172
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93526 32116 93536 32172
rect 130072 32116 130082 32172
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130346 32116 130356 32172
rect 62626 31948 62636 32004
rect 62692 31948 128156 32004
rect 128212 31948 128222 32004
rect 33058 31836 33068 31892
rect 33124 31836 62076 31892
rect 62132 31836 62142 31892
rect 69682 31836 69692 31892
rect 69748 31836 138012 31892
rect 138068 31836 138078 31892
rect 76738 31724 76748 31780
rect 76804 31724 143724 31780
rect 143780 31724 143790 31780
rect 66434 31612 66444 31668
rect 66500 31612 125916 31668
rect 125972 31612 125982 31668
rect 57698 31500 57708 31556
rect 57764 31500 109116 31556
rect 109172 31500 109182 31556
rect 38022 31332 38032 31388
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38296 31332 38306 31388
rect 74842 31332 74852 31388
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 75116 31332 75126 31388
rect 111662 31332 111672 31388
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111936 31332 111946 31388
rect 148482 31332 148492 31388
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148756 31332 148766 31388
rect 19282 31164 19292 31220
rect 19348 31164 25116 31220
rect 25172 31164 25182 31220
rect 56018 31164 56028 31220
rect 56084 31164 96348 31220
rect 96404 31164 96414 31220
rect 14242 31052 14252 31108
rect 14308 31052 53340 31108
rect 53396 31052 53406 31108
rect 54338 31052 54348 31108
rect 54404 31052 103740 31108
rect 103796 31052 103806 31108
rect 24994 30940 25004 30996
rect 25060 30940 81452 30996
rect 81508 30940 81518 30996
rect 64754 30828 64764 30884
rect 64820 30828 105084 30884
rect 105140 30828 105150 30884
rect 19612 30548 19622 30604
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19886 30548 19896 30604
rect 56432 30548 56442 30604
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56706 30548 56716 30604
rect 93252 30548 93262 30604
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93526 30548 93536 30604
rect 130072 30548 130082 30604
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130346 30548 130356 30604
rect 51986 30156 51996 30212
rect 52052 30156 58156 30212
rect 58212 30156 58222 30212
rect 68002 30156 68012 30212
rect 68068 30156 135996 30212
rect 136052 30156 136062 30212
rect 58930 30044 58940 30100
rect 58996 30044 123564 30100
rect 123620 30044 123630 30100
rect 55346 29932 55356 29988
rect 55412 29932 105532 29988
rect 105588 29932 105598 29988
rect 38022 29764 38032 29820
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38296 29764 38306 29820
rect 74842 29764 74852 29820
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 75116 29764 75126 29820
rect 111662 29764 111672 29820
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111936 29764 111946 29820
rect 148482 29764 148492 29820
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148756 29764 148766 29820
rect 52434 29596 52444 29652
rect 52500 29596 98364 29652
rect 98420 29596 98430 29652
rect 57474 29484 57484 29540
rect 57540 29484 102060 29540
rect 102116 29484 102126 29540
rect 16482 29372 16492 29428
rect 16548 29372 26908 29428
rect 26964 29372 26974 29428
rect 36306 29260 36316 29316
rect 36372 29260 83916 29316
rect 83972 29260 83982 29316
rect 34850 29148 34860 29204
rect 34916 29148 84364 29204
rect 84420 29148 84430 29204
rect 19612 28980 19622 29036
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19886 28980 19896 29036
rect 56432 28980 56442 29036
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56706 28980 56716 29036
rect 93252 28980 93262 29036
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93526 28980 93536 29036
rect 130072 28980 130082 29036
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130346 28980 130356 29036
rect 44482 28812 44492 28868
rect 44548 28812 91196 28868
rect 91252 28812 91262 28868
rect 69010 28476 69020 28532
rect 69076 28476 126140 28532
rect 126196 28476 126206 28532
rect 41122 28364 41132 28420
rect 41188 28364 95116 28420
rect 95172 28364 95182 28420
rect 38022 28196 38032 28252
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38296 28196 38306 28252
rect 74842 28196 74852 28252
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 75116 28196 75126 28252
rect 111662 28196 111672 28252
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111936 28196 111946 28252
rect 148482 28196 148492 28252
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148756 28196 148766 28252
rect 49858 28028 49868 28084
rect 49924 28028 101164 28084
rect 101220 28028 101230 28084
rect 62962 27916 62972 27972
rect 63028 27916 113596 27972
rect 113652 27916 113662 27972
rect 59938 27804 59948 27860
rect 60004 27804 90860 27860
rect 90916 27804 90926 27860
rect 96562 27692 96572 27748
rect 96628 27692 120316 27748
rect 120372 27692 120382 27748
rect 28354 27580 28364 27636
rect 28420 27580 79212 27636
rect 79268 27580 79278 27636
rect 19612 27412 19622 27468
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19886 27412 19896 27468
rect 56432 27412 56442 27468
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56706 27412 56716 27468
rect 93252 27412 93262 27468
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93526 27412 93536 27468
rect 130072 27412 130082 27468
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130346 27412 130356 27468
rect 39442 27244 39452 27300
rect 39508 27244 93884 27300
rect 93940 27244 93950 27300
rect 43586 27132 43596 27188
rect 43652 27132 97132 27188
rect 97188 27132 97198 27188
rect 45266 26908 45276 26964
rect 45332 26908 47068 26964
rect 47124 26908 47134 26964
rect 60274 26796 60284 26852
rect 60340 26796 128156 26852
rect 128212 26796 128222 26852
rect 38022 26628 38032 26684
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38296 26628 38306 26684
rect 74842 26628 74852 26684
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 75116 26628 75126 26684
rect 111662 26628 111672 26684
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111936 26628 111946 26684
rect 148482 26628 148492 26684
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148756 26628 148766 26684
rect 26898 26460 26908 26516
rect 26964 26460 27804 26516
rect 27860 26460 83804 26516
rect 83860 26460 83870 26516
rect 32610 26348 32620 26404
rect 32676 26348 86380 26404
rect 86436 26348 86446 26404
rect 50306 26236 50316 26292
rect 50372 26236 98028 26292
rect 98084 26236 98094 26292
rect 44594 26124 44604 26180
rect 44660 26124 89628 26180
rect 89684 26124 89694 26180
rect 91522 26124 91532 26180
rect 91588 26124 116284 26180
rect 116340 26124 116350 26180
rect 49522 26012 49532 26068
rect 49588 26012 51660 26068
rect 51716 26012 51726 26068
rect 83122 26012 83132 26068
rect 83188 26012 111468 26068
rect 111524 26012 111534 26068
rect 19612 25844 19622 25900
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19886 25844 19896 25900
rect 56432 25844 56442 25900
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56706 25844 56716 25900
rect 93252 25844 93262 25900
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93526 25844 93536 25900
rect 130072 25844 130082 25900
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130346 25844 130356 25900
rect 24322 25676 24332 25732
rect 24388 25676 82796 25732
rect 82852 25676 82862 25732
rect 25106 25564 25116 25620
rect 25172 25564 90300 25620
rect 90356 25564 90366 25620
rect 67890 25452 67900 25508
rect 67956 25452 109676 25508
rect 109732 25452 109742 25508
rect 38022 25060 38032 25116
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38296 25060 38306 25116
rect 74842 25060 74852 25116
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 75116 25060 75126 25116
rect 111662 25060 111672 25116
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111936 25060 111946 25116
rect 148482 25060 148492 25116
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148756 25060 148766 25116
rect 75506 24668 75516 24724
rect 75572 24668 103292 24724
rect 103348 24668 103358 24724
rect 73042 24556 73052 24612
rect 73108 24556 106652 24612
rect 106708 24556 106718 24612
rect 48402 24444 48412 24500
rect 48468 24444 81452 24500
rect 81508 24444 81518 24500
rect 19612 24276 19622 24332
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19886 24276 19896 24332
rect 56432 24276 56442 24332
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56706 24276 56716 24332
rect 93252 24276 93262 24332
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93526 24276 93536 24332
rect 130072 24276 130082 24332
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130346 24276 130356 24332
rect 38022 23492 38032 23548
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38296 23492 38306 23548
rect 74842 23492 74852 23548
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 75116 23492 75126 23548
rect 111662 23492 111672 23548
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111936 23492 111946 23548
rect 148482 23492 148492 23548
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148756 23492 148766 23548
rect 39890 22876 39900 22932
rect 39956 22876 68796 22932
rect 68852 22876 68862 22932
rect 19612 22708 19622 22764
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19886 22708 19896 22764
rect 56432 22708 56442 22764
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56706 22708 56716 22764
rect 93252 22708 93262 22764
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93526 22708 93536 22764
rect 130072 22708 130082 22764
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130346 22708 130356 22764
rect 38022 21924 38032 21980
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38296 21924 38306 21980
rect 74842 21924 74852 21980
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 75116 21924 75126 21980
rect 111662 21924 111672 21980
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111936 21924 111946 21980
rect 148482 21924 148492 21980
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148756 21924 148766 21980
rect 19612 21140 19622 21196
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19886 21140 19896 21196
rect 56432 21140 56442 21196
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56706 21140 56716 21196
rect 93252 21140 93262 21196
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93526 21140 93536 21196
rect 130072 21140 130082 21196
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130346 21140 130356 21196
rect 41234 20972 41244 21028
rect 41300 20972 69804 21028
rect 69860 20972 69870 21028
rect 71362 20972 71372 21028
rect 71428 20972 86604 21028
rect 86660 20972 86670 21028
rect 38022 20356 38032 20412
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38296 20356 38306 20412
rect 74842 20356 74852 20412
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 75116 20356 75126 20412
rect 111662 20356 111672 20412
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111936 20356 111946 20412
rect 148482 20356 148492 20412
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148756 20356 148766 20412
rect 19612 19572 19622 19628
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19886 19572 19896 19628
rect 56432 19572 56442 19628
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56706 19572 56716 19628
rect 93252 19572 93262 19628
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93526 19572 93536 19628
rect 130072 19572 130082 19628
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130346 19572 130356 19628
rect 42914 19404 42924 19460
rect 42980 19404 74172 19460
rect 74228 19404 74238 19460
rect 55234 19292 55244 19348
rect 55300 19292 98140 19348
rect 98196 19292 98206 19348
rect 38022 18788 38032 18844
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38296 18788 38306 18844
rect 74842 18788 74852 18844
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 75116 18788 75126 18844
rect 111662 18788 111672 18844
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111936 18788 111946 18844
rect 148482 18788 148492 18844
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148756 18788 148766 18844
rect 19612 18004 19622 18060
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19886 18004 19896 18060
rect 56432 18004 56442 18060
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56706 18004 56716 18060
rect 93252 18004 93262 18060
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93526 18004 93536 18060
rect 130072 18004 130082 18060
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130346 18004 130356 18060
rect 68898 17724 68908 17780
rect 68964 17724 104412 17780
rect 104468 17724 104478 17780
rect 46050 17612 46060 17668
rect 46116 17612 85820 17668
rect 85876 17612 85886 17668
rect 104178 17612 104188 17668
rect 104244 17612 121996 17668
rect 122052 17612 122062 17668
rect 38022 17220 38032 17276
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38296 17220 38306 17276
rect 74842 17220 74852 17276
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 75116 17220 75126 17276
rect 111662 17220 111672 17276
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111936 17220 111946 17276
rect 148482 17220 148492 17276
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148756 17220 148766 17276
rect 19612 16436 19622 16492
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19886 16436 19896 16492
rect 56432 16436 56442 16492
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56706 16436 56716 16492
rect 93252 16436 93262 16492
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93526 16436 93536 16492
rect 130072 16436 130082 16492
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130346 16436 130356 16492
rect 38022 15652 38032 15708
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38296 15652 38306 15708
rect 74842 15652 74852 15708
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 75116 15652 75126 15708
rect 111662 15652 111672 15708
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111936 15652 111946 15708
rect 148482 15652 148492 15708
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148756 15652 148766 15708
rect 67330 15372 67340 15428
rect 67396 15372 68796 15428
rect 68852 15372 68862 15428
rect 19612 14868 19622 14924
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19886 14868 19896 14924
rect 56432 14868 56442 14924
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56706 14868 56716 14924
rect 93252 14868 93262 14924
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93526 14868 93536 14924
rect 130072 14868 130082 14924
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130346 14868 130356 14924
rect 52994 14252 53004 14308
rect 53060 14252 59052 14308
rect 59108 14252 59118 14308
rect 60274 14252 60284 14308
rect 60340 14252 80108 14308
rect 80164 14252 80174 14308
rect 38022 14084 38032 14140
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38296 14084 38306 14140
rect 74842 14084 74852 14140
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 75116 14084 75126 14140
rect 111662 14084 111672 14140
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111936 14084 111946 14140
rect 148482 14084 148492 14140
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148756 14084 148766 14140
rect 19612 13300 19622 13356
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19886 13300 19896 13356
rect 56432 13300 56442 13356
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56706 13300 56716 13356
rect 93252 13300 93262 13356
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93526 13300 93536 13356
rect 130072 13300 130082 13356
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130346 13300 130356 13356
rect 57810 12684 57820 12740
rect 57876 12684 78204 12740
rect 78260 12684 78270 12740
rect 81442 12684 81452 12740
rect 81508 12684 113148 12740
rect 113204 12684 113214 12740
rect 113362 12572 113372 12628
rect 113428 12572 118524 12628
rect 118580 12572 118590 12628
rect 38022 12516 38032 12572
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38296 12516 38306 12572
rect 74842 12516 74852 12572
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 75116 12516 75126 12572
rect 111662 12516 111672 12572
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111936 12516 111946 12572
rect 148482 12516 148492 12572
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148756 12516 148766 12572
rect 98130 11788 98140 11844
rect 98196 11788 104188 11844
rect 104244 11788 104254 11844
rect 19612 11732 19622 11788
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19886 11732 19896 11788
rect 56432 11732 56442 11788
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56706 11732 56716 11788
rect 93252 11732 93262 11788
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93526 11732 93536 11788
rect 130072 11732 130082 11788
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130346 11732 130356 11788
rect 85810 11676 85820 11732
rect 85876 11676 91532 11732
rect 91588 11676 91598 11732
rect 36082 11564 36092 11620
rect 36148 11564 59052 11620
rect 59108 11564 60284 11620
rect 60340 11564 60350 11620
rect 48626 11228 48636 11284
rect 48692 11228 89068 11284
rect 89124 11228 89134 11284
rect 75730 11116 75740 11172
rect 75796 11116 120764 11172
rect 120820 11116 120830 11172
rect 38022 10948 38032 11004
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38296 10948 38306 11004
rect 74842 10948 74852 11004
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 75116 10948 75126 11004
rect 111662 10948 111672 11004
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111936 10948 111946 11004
rect 148482 10948 148492 11004
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148756 10948 148766 11004
rect 19612 10164 19622 10220
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19886 10164 19896 10220
rect 56432 10164 56442 10220
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56706 10164 56716 10220
rect 93252 10164 93262 10220
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93526 10164 93536 10220
rect 130072 10164 130082 10220
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130346 10164 130356 10220
rect 38022 9380 38032 9436
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38296 9380 38306 9436
rect 74842 9380 74852 9436
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 75116 9380 75126 9436
rect 111662 9380 111672 9436
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111936 9380 111946 9436
rect 148482 9380 148492 9436
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148756 9380 148766 9436
rect 18162 9324 18172 9380
rect 18228 9324 33516 9380
rect 33572 9324 33582 9380
rect 14578 9212 14588 9268
rect 14644 9212 26460 9268
rect 26516 9212 26526 9268
rect 32386 9212 32396 9268
rect 32452 9212 59612 9268
rect 59668 9212 59678 9268
rect 103282 8876 103292 8932
rect 103348 8876 123116 8932
rect 123172 8876 124124 8932
rect 124180 8876 124190 8932
rect 124338 8876 124348 8932
rect 124404 8876 124908 8932
rect 124964 8876 125468 8932
rect 125524 8876 136780 8932
rect 136836 8876 136846 8932
rect 19612 8596 19622 8652
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19886 8596 19896 8652
rect 56432 8596 56442 8652
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56706 8596 56716 8652
rect 93252 8596 93262 8652
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93526 8596 93536 8652
rect 130072 8596 130082 8652
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130346 8596 130356 8652
rect 62178 8428 62188 8484
rect 62244 8428 64540 8484
rect 64596 8428 64606 8484
rect 123554 8428 123564 8484
rect 123620 8428 124124 8484
rect 124180 8428 124190 8484
rect 65762 8316 65772 8372
rect 65828 8316 68348 8372
rect 68404 8316 68414 8372
rect 120754 8316 120764 8372
rect 120820 8316 121884 8372
rect 121940 8316 122780 8372
rect 122836 8316 122846 8372
rect 124786 8316 124796 8372
rect 124852 8316 125916 8372
rect 125972 8316 125982 8372
rect 63634 8204 63644 8260
rect 63700 8204 64540 8260
rect 64596 8204 67004 8260
rect 67060 8204 67070 8260
rect 87938 8204 87948 8260
rect 88004 8204 89404 8260
rect 89460 8204 89470 8260
rect 89852 8204 90748 8260
rect 90804 8204 90814 8260
rect 94770 8204 94780 8260
rect 94836 8204 96124 8260
rect 96180 8204 96190 8260
rect 105746 8204 105756 8260
rect 105812 8204 106652 8260
rect 106708 8204 107100 8260
rect 107156 8204 107166 8260
rect 123778 8204 123788 8260
rect 123844 8204 125244 8260
rect 125300 8204 125310 8260
rect 89852 8148 89908 8204
rect 58146 8092 58156 8148
rect 58212 8092 63980 8148
rect 64036 8092 65436 8148
rect 65492 8092 66556 8148
rect 66612 8092 66622 8148
rect 82898 8092 82908 8148
rect 82964 8092 88508 8148
rect 88564 8092 89852 8148
rect 89908 8092 89918 8148
rect 90066 8092 90076 8148
rect 90132 8092 93604 8148
rect 93762 8092 93772 8148
rect 93828 8092 94892 8148
rect 94948 8092 95564 8148
rect 95620 8092 105532 8148
rect 105588 8092 105980 8148
rect 106036 8092 106046 8148
rect 123442 8092 123452 8148
rect 123508 8092 124348 8148
rect 124404 8092 125972 8148
rect 93548 8036 93604 8092
rect 125916 8036 125972 8092
rect 28018 7980 28028 8036
rect 28084 7980 28924 8036
rect 28980 7980 28990 8036
rect 65986 7980 65996 8036
rect 66052 7980 85484 8036
rect 85540 7980 86044 8036
rect 86100 7980 92540 8036
rect 92596 7980 93100 8036
rect 93156 7980 93166 8036
rect 93548 7980 95340 8036
rect 95396 7980 96684 8036
rect 96740 7980 98028 8036
rect 98084 7980 98094 8036
rect 102946 7980 102956 8036
rect 103012 7980 103964 8036
rect 104020 7980 106316 8036
rect 106372 7980 106382 8036
rect 123106 7980 123116 8036
rect 123172 7980 125020 8036
rect 125076 7980 125086 8036
rect 125906 7980 125916 8036
rect 125972 7980 125982 8036
rect 126802 7980 126812 8036
rect 126868 7980 137116 8036
rect 137172 7980 137182 8036
rect 126812 7924 126868 7980
rect 123330 7868 123340 7924
rect 123396 7868 126868 7924
rect 127250 7868 127260 7924
rect 127316 7868 135660 7924
rect 135716 7868 135726 7924
rect 38022 7812 38032 7868
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38296 7812 38306 7868
rect 74842 7812 74852 7868
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 75116 7812 75126 7868
rect 111662 7812 111672 7868
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111936 7812 111946 7868
rect 148482 7812 148492 7868
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148756 7812 148766 7868
rect 125906 7756 125916 7812
rect 125972 7756 139916 7812
rect 139972 7756 139982 7812
rect 66434 7644 66444 7700
rect 66500 7644 67228 7700
rect 67284 7644 67294 7700
rect 87714 7644 87724 7700
rect 87780 7644 89180 7700
rect 89236 7644 89246 7700
rect 95106 7644 95116 7700
rect 95172 7644 96012 7700
rect 96068 7644 96078 7700
rect 105970 7644 105980 7700
rect 106036 7644 107100 7700
rect 107156 7644 107166 7700
rect 125794 7644 125804 7700
rect 125860 7644 126812 7700
rect 126868 7644 126878 7700
rect 137554 7644 137564 7700
rect 137620 7644 139132 7700
rect 139188 7644 139692 7700
rect 139748 7644 139758 7700
rect 7858 7532 7868 7588
rect 7924 7532 15708 7588
rect 15764 7532 15774 7588
rect 26562 7532 26572 7588
rect 26628 7532 27244 7588
rect 27300 7532 27310 7588
rect 57698 7532 57708 7588
rect 57764 7532 59164 7588
rect 59220 7532 59230 7588
rect 62850 7532 62860 7588
rect 62916 7532 64204 7588
rect 64260 7532 66892 7588
rect 66948 7532 66958 7588
rect 87042 7532 87052 7588
rect 87108 7532 87836 7588
rect 87892 7532 88284 7588
rect 88340 7532 88350 7588
rect 104066 7532 104076 7588
rect 104132 7532 105420 7588
rect 105476 7532 105486 7588
rect 115378 7532 115388 7588
rect 115444 7532 116620 7588
rect 116676 7532 118300 7588
rect 118356 7532 118366 7588
rect 26674 7420 26684 7476
rect 26740 7420 28028 7476
rect 28084 7420 28094 7476
rect 28578 7420 28588 7476
rect 28644 7420 30380 7476
rect 30436 7420 30446 7476
rect 59490 7420 59500 7476
rect 59556 7420 60956 7476
rect 61012 7420 61022 7476
rect 62066 7420 62076 7476
rect 62132 7420 63420 7476
rect 63476 7420 63868 7476
rect 63924 7420 65548 7476
rect 65604 7420 65614 7476
rect 77074 7420 77084 7476
rect 77140 7420 78428 7476
rect 78484 7420 78494 7476
rect 86258 7420 86268 7476
rect 86324 7420 94444 7476
rect 94500 7420 96460 7476
rect 96516 7420 98924 7476
rect 98980 7420 98990 7476
rect 105746 7420 105756 7476
rect 105812 7420 106764 7476
rect 106820 7420 107548 7476
rect 107604 7420 107614 7476
rect 116386 7420 116396 7476
rect 116452 7420 117740 7476
rect 117796 7420 117806 7476
rect 19282 7308 19292 7364
rect 19348 7308 20300 7364
rect 20356 7308 26908 7364
rect 26964 7308 28364 7364
rect 28420 7308 28812 7364
rect 28868 7308 29932 7364
rect 29988 7308 29998 7364
rect 44146 7308 44156 7364
rect 44212 7308 45164 7364
rect 45220 7308 46172 7364
rect 46228 7308 47180 7364
rect 47236 7308 47246 7364
rect 51650 7308 51660 7364
rect 51716 7308 56252 7364
rect 56308 7308 56318 7364
rect 88386 7308 88396 7364
rect 88452 7308 89628 7364
rect 89684 7308 89694 7364
rect 103058 7308 103068 7364
rect 103124 7308 103516 7364
rect 103572 7308 106316 7364
rect 106372 7308 106382 7364
rect 116946 7308 116956 7364
rect 117012 7308 118188 7364
rect 118244 7308 118254 7364
rect 47180 7252 47236 7308
rect 27122 7196 27132 7252
rect 27188 7196 28252 7252
rect 28308 7196 28318 7252
rect 47180 7196 52556 7252
rect 52612 7196 53452 7252
rect 53508 7196 54572 7252
rect 54628 7196 54638 7252
rect 61618 7196 61628 7252
rect 61684 7196 63532 7252
rect 63588 7196 66108 7252
rect 66164 7196 66174 7252
rect 115042 7196 115052 7252
rect 115108 7196 116060 7252
rect 116116 7196 116126 7252
rect 126354 7196 126364 7252
rect 126420 7196 135772 7252
rect 135828 7196 135838 7252
rect 76402 7084 76412 7140
rect 76468 7084 76860 7140
rect 76916 7084 77980 7140
rect 78036 7084 86492 7140
rect 86548 7084 86558 7140
rect 123330 7084 123340 7140
rect 123396 7084 127260 7140
rect 127316 7084 127326 7140
rect 19612 7028 19622 7084
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19886 7028 19896 7084
rect 56432 7028 56442 7084
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56706 7028 56716 7084
rect 93252 7028 93262 7084
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93526 7028 93536 7084
rect 130072 7028 130082 7084
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130346 7028 130356 7084
rect 19618 6860 19628 6916
rect 19684 6860 19964 6916
rect 20020 6860 20524 6916
rect 20580 6860 20590 6916
rect 43362 6860 43372 6916
rect 43428 6860 44940 6916
rect 44996 6860 45006 6916
rect 45938 6860 45948 6916
rect 46004 6860 47852 6916
rect 47908 6860 47918 6916
rect 126130 6860 126140 6916
rect 126196 6860 143948 6916
rect 144004 6860 144014 6916
rect 75618 6748 75628 6804
rect 75684 6748 77756 6804
rect 77812 6748 78540 6804
rect 78596 6748 78606 6804
rect 114258 6748 114268 6804
rect 114324 6748 117516 6804
rect 117572 6748 117582 6804
rect 139346 6748 139356 6804
rect 139412 6748 140252 6804
rect 140308 6748 140812 6804
rect 140868 6748 140878 6804
rect 18274 6636 18284 6692
rect 18340 6636 27692 6692
rect 27748 6636 27758 6692
rect 44594 6636 44604 6692
rect 44660 6636 45612 6692
rect 45668 6636 45678 6692
rect 64642 6636 64652 6692
rect 64708 6636 66332 6692
rect 66388 6636 67676 6692
rect 67732 6636 68124 6692
rect 68180 6636 68190 6692
rect 68562 6636 68572 6692
rect 68628 6636 69356 6692
rect 69412 6636 69422 6692
rect 87042 6636 87052 6692
rect 87108 6636 95452 6692
rect 95508 6636 95676 6692
rect 95732 6636 102508 6692
rect 102564 6636 102574 6692
rect 104402 6636 104412 6692
rect 104468 6636 105980 6692
rect 106036 6636 106046 6692
rect 122658 6636 122668 6692
rect 122724 6636 124908 6692
rect 124964 6636 126252 6692
rect 126308 6636 126318 6692
rect 136770 6636 136780 6692
rect 136836 6636 138124 6692
rect 138180 6636 138190 6692
rect 27906 6524 27916 6580
rect 27972 6524 29596 6580
rect 29652 6524 38892 6580
rect 38948 6524 39452 6580
rect 39508 6524 39518 6580
rect 59938 6524 59948 6580
rect 60004 6524 61852 6580
rect 61908 6524 61918 6580
rect 104738 6524 104748 6580
rect 104804 6524 106092 6580
rect 106148 6524 106158 6580
rect 135986 6524 135996 6580
rect 136052 6524 137788 6580
rect 137844 6524 137854 6580
rect 138450 6524 138460 6580
rect 138516 6524 139132 6580
rect 139188 6524 141260 6580
rect 141316 6524 141326 6580
rect 14578 6412 14588 6468
rect 14644 6412 15484 6468
rect 15540 6412 18732 6468
rect 18788 6412 18798 6468
rect 27346 6412 27356 6468
rect 27412 6412 28252 6468
rect 28308 6412 28318 6468
rect 50530 6412 50540 6468
rect 50596 6412 50988 6468
rect 51044 6412 51054 6468
rect 60274 6412 60284 6468
rect 60340 6412 61292 6468
rect 61348 6412 62412 6468
rect 62468 6412 62478 6468
rect 76290 6412 76300 6468
rect 76356 6412 79100 6468
rect 79156 6412 80892 6468
rect 80948 6412 80958 6468
rect 95330 6412 95340 6468
rect 95396 6412 95788 6468
rect 95844 6412 95854 6468
rect 105746 6412 105756 6468
rect 105812 6412 107100 6468
rect 107156 6412 107166 6468
rect 113698 6412 113708 6468
rect 113764 6412 114716 6468
rect 114772 6412 114782 6468
rect 123778 6412 123788 6468
rect 123844 6412 126588 6468
rect 126644 6412 126654 6468
rect 128370 6412 128380 6468
rect 128436 6412 129388 6468
rect 129444 6412 129454 6468
rect 51314 6300 51324 6356
rect 51380 6300 52668 6356
rect 52724 6300 54012 6356
rect 54068 6300 65996 6356
rect 66052 6300 66062 6356
rect 117170 6300 117180 6356
rect 117236 6300 128604 6356
rect 128660 6300 132188 6356
rect 132244 6300 132254 6356
rect 38022 6244 38032 6300
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38296 6244 38306 6300
rect 74842 6244 74852 6300
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 75116 6244 75126 6300
rect 111662 6244 111672 6300
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111936 6244 111946 6300
rect 148482 6244 148492 6300
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148756 6244 148766 6300
rect 29362 6188 29372 6244
rect 29428 6188 31388 6244
rect 31444 6188 31454 6244
rect 114212 6188 131908 6244
rect 135762 6188 135772 6244
rect 135828 6188 137452 6244
rect 137508 6188 137518 6244
rect 114212 6132 114268 6188
rect 16146 6076 16156 6132
rect 16212 6076 17612 6132
rect 17668 6076 17678 6132
rect 26012 6076 39788 6132
rect 39844 6076 39854 6132
rect 55234 6076 55244 6132
rect 55300 6076 55692 6132
rect 55748 6076 55758 6132
rect 63074 6076 63084 6132
rect 63140 6076 63980 6132
rect 64036 6076 64046 6132
rect 66098 6076 66108 6132
rect 66164 6076 67564 6132
rect 67620 6076 67630 6132
rect 84578 6076 84588 6132
rect 84644 6076 95564 6132
rect 95620 6076 95630 6132
rect 103730 6076 103740 6132
rect 103796 6076 104412 6132
rect 104468 6076 104478 6132
rect 108210 6076 108220 6132
rect 108276 6076 109228 6132
rect 109284 6076 109294 6132
rect 110786 6076 110796 6132
rect 110852 6076 114268 6132
rect 125570 6076 125580 6132
rect 125636 6076 127260 6132
rect 127316 6076 127326 6132
rect 127474 6076 127484 6132
rect 127540 6076 129388 6132
rect 129444 6076 129454 6132
rect 17714 5964 17724 6020
rect 17780 5964 19628 6020
rect 19684 5964 19694 6020
rect 15922 5852 15932 5908
rect 15988 5852 17836 5908
rect 17892 5852 17902 5908
rect 18162 5852 18172 5908
rect 18228 5852 18844 5908
rect 18900 5852 21532 5908
rect 21588 5852 21598 5908
rect 26012 5796 26068 6076
rect 131852 6020 131908 6188
rect 132402 6076 132412 6132
rect 132468 6076 134204 6132
rect 134260 6076 134270 6132
rect 137330 6076 137340 6132
rect 137396 6076 138572 6132
rect 138628 6076 138638 6132
rect 27682 5964 27692 6020
rect 27748 5964 31724 6020
rect 31780 5964 31948 6020
rect 52882 5964 52892 6020
rect 52948 5964 53116 6020
rect 53172 5964 60732 6020
rect 60788 5964 61740 6020
rect 61796 5964 61806 6020
rect 76514 5964 76524 6020
rect 76580 5964 79884 6020
rect 79940 5964 79950 6020
rect 108322 5964 108332 6020
rect 108388 5964 109340 6020
rect 109396 5964 110236 6020
rect 110292 5964 114940 6020
rect 114996 5964 115006 6020
rect 128034 5964 128044 6020
rect 128100 5964 130844 6020
rect 130900 5964 130910 6020
rect 131852 5964 139804 6020
rect 139860 5964 140140 6020
rect 140196 5964 140700 6020
rect 140756 5964 140766 6020
rect 31892 5908 31948 5964
rect 31892 5852 43820 5908
rect 43876 5852 47628 5908
rect 47684 5852 55356 5908
rect 55412 5852 57148 5908
rect 57204 5852 57820 5908
rect 57876 5852 59836 5908
rect 59892 5852 60284 5908
rect 60340 5852 60350 5908
rect 77634 5852 77644 5908
rect 77700 5852 78764 5908
rect 78820 5852 78830 5908
rect 79426 5852 79436 5908
rect 79492 5852 80444 5908
rect 80500 5852 80510 5908
rect 102498 5852 102508 5908
rect 102564 5852 104524 5908
rect 104580 5852 105308 5908
rect 105364 5852 106652 5908
rect 106708 5852 112364 5908
rect 112420 5852 113260 5908
rect 113316 5852 120204 5908
rect 120260 5852 121996 5908
rect 122052 5852 122444 5908
rect 122500 5852 122510 5908
rect 125234 5852 125244 5908
rect 125300 5852 133028 5908
rect 133186 5852 133196 5908
rect 133252 5852 133756 5908
rect 133812 5852 133822 5908
rect 137732 5852 137900 5908
rect 137956 5852 137966 5908
rect 138114 5852 138124 5908
rect 138180 5852 139020 5908
rect 139076 5852 139580 5908
rect 139636 5852 139646 5908
rect 132972 5796 133028 5852
rect 137732 5796 137788 5852
rect 16706 5740 16716 5796
rect 16772 5740 17500 5796
rect 17556 5740 26068 5796
rect 47730 5740 47740 5796
rect 47796 5740 58268 5796
rect 58324 5740 59388 5796
rect 59444 5740 63308 5796
rect 63364 5740 63374 5796
rect 110908 5740 111580 5796
rect 111636 5740 115388 5796
rect 115444 5740 115454 5796
rect 127586 5740 127596 5796
rect 127652 5740 131964 5796
rect 132020 5740 132030 5796
rect 132972 5740 135212 5796
rect 135268 5740 137788 5796
rect 110908 5684 110964 5740
rect 39442 5628 39452 5684
rect 39508 5628 50540 5684
rect 50596 5628 50606 5684
rect 55682 5628 55692 5684
rect 55748 5628 58884 5684
rect 70130 5628 70140 5684
rect 70196 5628 75740 5684
rect 75796 5628 75806 5684
rect 89618 5628 89628 5684
rect 89684 5628 96572 5684
rect 96628 5628 97244 5684
rect 97300 5628 98364 5684
rect 98420 5628 98924 5684
rect 98980 5628 102732 5684
rect 102788 5628 103180 5684
rect 103236 5628 103628 5684
rect 103684 5628 104300 5684
rect 104356 5628 104366 5684
rect 110226 5628 110236 5684
rect 110292 5628 110908 5684
rect 110964 5628 110974 5684
rect 125794 5628 125804 5684
rect 125860 5628 127932 5684
rect 127988 5628 127998 5684
rect 132962 5628 132972 5684
rect 133028 5628 134652 5684
rect 134708 5628 134718 5684
rect 58828 5572 58884 5628
rect 45938 5516 45948 5572
rect 46004 5516 46508 5572
rect 46564 5516 47292 5572
rect 47348 5516 47358 5572
rect 58818 5516 58828 5572
rect 58884 5516 58894 5572
rect 126690 5516 126700 5572
rect 126756 5516 127372 5572
rect 127428 5516 128044 5572
rect 128100 5516 129052 5572
rect 129108 5516 129118 5572
rect 132178 5516 132188 5572
rect 132244 5516 133980 5572
rect 134036 5516 134046 5572
rect 134194 5516 134204 5572
rect 134260 5516 138684 5572
rect 138740 5516 138750 5572
rect 19612 5460 19622 5516
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19886 5460 19896 5516
rect 56432 5460 56442 5516
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56706 5460 56716 5516
rect 93252 5460 93262 5516
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93526 5460 93536 5516
rect 130072 5460 130082 5516
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130346 5460 130356 5516
rect 20290 5404 20300 5460
rect 20356 5404 27916 5460
rect 27972 5404 27982 5460
rect 57922 5404 57932 5460
rect 57988 5404 60508 5460
rect 60564 5404 60574 5460
rect 66098 5404 66108 5460
rect 66164 5404 67676 5460
rect 67732 5404 67742 5460
rect 69132 5404 78988 5460
rect 69132 5348 69188 5404
rect 78932 5348 78988 5404
rect 131516 5404 137004 5460
rect 137060 5404 137070 5460
rect 137778 5404 137788 5460
rect 137844 5404 138460 5460
rect 138516 5404 138526 5460
rect 131516 5348 131572 5404
rect 19058 5292 19068 5348
rect 19124 5292 20748 5348
rect 20804 5292 20814 5348
rect 29698 5292 29708 5348
rect 29764 5292 30604 5348
rect 30660 5292 30670 5348
rect 39778 5292 39788 5348
rect 39844 5292 69188 5348
rect 69346 5292 69356 5348
rect 69412 5292 75572 5348
rect 78932 5292 111020 5348
rect 111076 5292 111086 5348
rect 118514 5292 118524 5348
rect 118580 5292 119532 5348
rect 119588 5292 119598 5348
rect 121202 5292 121212 5348
rect 121268 5292 123900 5348
rect 123956 5292 131572 5348
rect 131842 5292 131852 5348
rect 131908 5292 133420 5348
rect 133476 5292 133486 5348
rect 137218 5292 137228 5348
rect 137284 5292 138796 5348
rect 138852 5292 138862 5348
rect 75516 5236 75572 5292
rect 8866 5180 8876 5236
rect 8932 5180 15036 5236
rect 15092 5180 15102 5236
rect 26562 5180 26572 5236
rect 26628 5180 28588 5236
rect 28644 5180 28654 5236
rect 44146 5180 44156 5236
rect 44212 5180 46396 5236
rect 46452 5180 46462 5236
rect 46610 5180 46620 5236
rect 46676 5180 47180 5236
rect 47236 5180 47246 5236
rect 53666 5180 53676 5236
rect 53732 5180 54460 5236
rect 54516 5180 54526 5236
rect 54674 5180 54684 5236
rect 54740 5180 55692 5236
rect 55748 5180 55758 5236
rect 58258 5180 58268 5236
rect 58324 5180 59276 5236
rect 59332 5180 59342 5236
rect 62524 5180 63980 5236
rect 64036 5180 68908 5236
rect 68964 5180 69692 5236
rect 69748 5180 69758 5236
rect 75506 5180 75516 5236
rect 75572 5180 77420 5236
rect 77476 5180 78988 5236
rect 79044 5180 86828 5236
rect 86884 5180 86894 5236
rect 107538 5180 107548 5236
rect 107604 5180 109228 5236
rect 109284 5180 109294 5236
rect 109554 5180 109564 5236
rect 109620 5180 111356 5236
rect 111412 5180 111422 5236
rect 114930 5180 114940 5236
rect 114996 5180 115500 5236
rect 115556 5180 116284 5236
rect 116340 5180 116956 5236
rect 117012 5180 117852 5236
rect 117908 5180 117918 5236
rect 124338 5180 124348 5236
rect 124404 5180 126028 5236
rect 127250 5180 127260 5236
rect 127316 5180 132076 5236
rect 132132 5180 132142 5236
rect 132290 5180 132300 5236
rect 132356 5180 133364 5236
rect 133746 5180 133756 5236
rect 133812 5180 134204 5236
rect 134260 5180 134764 5236
rect 134820 5180 137788 5236
rect 137844 5180 137854 5236
rect 138226 5180 138236 5236
rect 138292 5180 139468 5236
rect 139524 5180 141596 5236
rect 141652 5180 141662 5236
rect 62524 5124 62580 5180
rect 125972 5124 126028 5180
rect 133308 5124 133364 5180
rect 7746 5068 7756 5124
rect 7812 5068 9884 5124
rect 9940 5068 11676 5124
rect 11732 5068 13748 5124
rect 17266 5068 17276 5124
rect 17332 5068 21532 5124
rect 21588 5068 25116 5124
rect 25172 5068 28700 5124
rect 28756 5068 41020 5124
rect 41076 5068 45388 5124
rect 45444 5068 62580 5124
rect 62850 5068 62860 5124
rect 62916 5068 63868 5124
rect 63924 5068 67116 5124
rect 67172 5068 70700 5124
rect 70756 5068 70766 5124
rect 75282 5068 75292 5124
rect 75348 5068 77756 5124
rect 77812 5068 77822 5124
rect 78418 5068 78428 5124
rect 78484 5068 80444 5124
rect 80500 5068 85932 5124
rect 85988 5068 86380 5124
rect 86436 5068 93884 5124
rect 93940 5068 94556 5124
rect 94612 5068 102620 5124
rect 102676 5068 103964 5124
rect 104020 5068 105308 5124
rect 105364 5068 106764 5124
rect 106820 5068 114380 5124
rect 114436 5068 114446 5124
rect 115602 5068 115612 5124
rect 115668 5068 116172 5124
rect 116228 5068 116238 5124
rect 121314 5068 121324 5124
rect 121380 5068 124908 5124
rect 124964 5068 125244 5124
rect 125300 5068 125310 5124
rect 125972 5068 129388 5124
rect 129444 5068 129454 5124
rect 130274 5068 130284 5124
rect 130340 5068 133084 5124
rect 133140 5068 133150 5124
rect 133308 5068 134204 5124
rect 134260 5068 134270 5124
rect 137442 5068 137452 5124
rect 137508 5068 139692 5124
rect 139748 5068 139758 5124
rect 13692 5012 13748 5068
rect 17276 5012 17332 5068
rect 12114 4956 12124 5012
rect 12180 4956 12684 5012
rect 12740 4956 12750 5012
rect 13682 4956 13692 5012
rect 13748 4956 17332 5012
rect 57474 4956 57484 5012
rect 57540 4956 58156 5012
rect 58212 4956 59276 5012
rect 59332 4956 59342 5012
rect 60610 4956 60620 5012
rect 60676 4956 62188 5012
rect 62244 4956 62254 5012
rect 69794 4956 69804 5012
rect 69860 4956 73052 5012
rect 73108 4956 73118 5012
rect 81330 4956 81340 5012
rect 81396 4956 85596 5012
rect 85652 4956 89404 5012
rect 89460 4956 89964 5012
rect 90020 4956 90412 5012
rect 90468 4956 90748 5012
rect 114818 4956 114828 5012
rect 114884 4956 117740 5012
rect 117796 4956 117806 5012
rect 120194 4956 120204 5012
rect 120260 4956 120876 5012
rect 120932 4956 120942 5012
rect 128034 4956 128044 5012
rect 128100 4956 135772 5012
rect 135828 4956 135838 5012
rect 60620 4900 60676 4956
rect 11330 4844 11340 4900
rect 11396 4844 14252 4900
rect 14308 4844 14318 4900
rect 20132 4844 20300 4900
rect 20356 4844 20366 4900
rect 29586 4844 29596 4900
rect 29652 4844 30156 4900
rect 30212 4844 30222 4900
rect 40226 4844 40236 4900
rect 40292 4844 44044 4900
rect 44100 4844 44716 4900
rect 44772 4844 44782 4900
rect 59042 4844 59052 4900
rect 59108 4844 60676 4900
rect 90692 4900 90748 4956
rect 90692 4844 90860 4900
rect 90916 4844 90926 4900
rect 133298 4844 133308 4900
rect 133364 4844 135996 4900
rect 136052 4844 136062 4900
rect 20132 4788 20188 4844
rect 5842 4732 5852 4788
rect 5908 4732 6188 4788
rect 6244 4732 8428 4788
rect 13346 4732 13356 4788
rect 13412 4732 16940 4788
rect 16996 4732 20188 4788
rect 59602 4732 59612 4788
rect 59668 4732 71372 4788
rect 71428 4732 71438 4788
rect 125458 4732 125468 4788
rect 125524 4732 129948 4788
rect 130004 4732 130014 4788
rect 8372 4676 8428 4732
rect 38022 4676 38032 4732
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38296 4676 38306 4732
rect 74842 4676 74852 4732
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 75116 4676 75126 4732
rect 111662 4676 111672 4732
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111936 4676 111946 4732
rect 148482 4676 148492 4732
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148756 4676 148766 4732
rect 8372 4620 16268 4676
rect 16324 4620 16334 4676
rect 127474 4620 127484 4676
rect 127540 4620 128156 4676
rect 128212 4620 130956 4676
rect 131012 4620 131022 4676
rect 15362 4508 15372 4564
rect 15428 4508 18732 4564
rect 18788 4508 18798 4564
rect 20132 4508 27132 4564
rect 27188 4508 29148 4564
rect 29204 4508 29214 4564
rect 48178 4508 48188 4564
rect 48244 4508 55244 4564
rect 55300 4508 55310 4564
rect 56802 4508 56812 4564
rect 56868 4508 58492 4564
rect 58548 4508 58558 4564
rect 70242 4508 70252 4564
rect 70308 4508 84476 4564
rect 84532 4508 85260 4564
rect 85316 4508 88508 4564
rect 88564 4508 89292 4564
rect 89348 4508 89358 4564
rect 108434 4508 108444 4564
rect 108500 4508 110908 4564
rect 110964 4508 112812 4564
rect 112868 4508 112878 4564
rect 123778 4508 123788 4564
rect 123844 4508 128044 4564
rect 128100 4508 128110 4564
rect 138338 4508 138348 4564
rect 138404 4508 140924 4564
rect 140980 4508 140990 4564
rect 20132 4452 20188 4508
rect 7746 4396 7756 4452
rect 7812 4396 10220 4452
rect 10276 4396 10286 4452
rect 12338 4396 12348 4452
rect 12404 4396 12684 4452
rect 12740 4396 12908 4452
rect 12964 4396 16156 4452
rect 16212 4396 16828 4452
rect 16884 4396 20188 4452
rect 20402 4396 20412 4452
rect 20468 4396 27468 4452
rect 27524 4396 28140 4452
rect 28196 4396 29596 4452
rect 29652 4396 29662 4452
rect 79874 4396 79884 4452
rect 79940 4396 80444 4452
rect 80500 4396 81340 4452
rect 81396 4396 81406 4452
rect 110450 4396 110460 4452
rect 110516 4396 111356 4452
rect 111412 4396 116732 4452
rect 116788 4396 116798 4452
rect 127474 4396 127484 4452
rect 127540 4396 129500 4452
rect 129556 4396 129566 4452
rect 6962 4284 6972 4340
rect 7028 4284 8988 4340
rect 9044 4284 9054 4340
rect 16258 4284 16268 4340
rect 16324 4284 17612 4340
rect 17668 4284 17948 4340
rect 18004 4284 18014 4340
rect 20514 4284 20524 4340
rect 20580 4284 22092 4340
rect 22148 4284 22540 4340
rect 22596 4284 22606 4340
rect 45042 4284 45052 4340
rect 45108 4284 53452 4340
rect 53508 4284 54012 4340
rect 54068 4284 54078 4340
rect 66882 4284 66892 4340
rect 66948 4284 68348 4340
rect 68404 4284 68414 4340
rect 70690 4284 70700 4340
rect 70756 4284 72604 4340
rect 72660 4284 74844 4340
rect 74900 4284 79100 4340
rect 79156 4284 79166 4340
rect 105746 4284 105756 4340
rect 105812 4284 107212 4340
rect 107268 4284 107278 4340
rect 114370 4284 114380 4340
rect 114436 4284 118524 4340
rect 118580 4284 120876 4340
rect 120932 4284 121548 4340
rect 121604 4284 122220 4340
rect 122276 4284 122892 4340
rect 122948 4284 128380 4340
rect 128436 4284 128940 4340
rect 128996 4284 129006 4340
rect 14466 4172 14476 4228
rect 14532 4172 15148 4228
rect 15204 4172 15214 4228
rect 16930 4172 16940 4228
rect 16996 4172 18172 4228
rect 18228 4172 18238 4228
rect 20290 4172 20300 4228
rect 20356 4172 20636 4228
rect 20692 4172 20702 4228
rect 24994 4172 25004 4228
rect 25060 4172 25900 4228
rect 25956 4172 25966 4228
rect 36306 4172 36316 4228
rect 36372 4172 37212 4228
rect 37268 4172 45948 4228
rect 46004 4172 46014 4228
rect 46162 4172 46172 4228
rect 46228 4172 47180 4228
rect 47236 4172 47246 4228
rect 51426 4172 51436 4228
rect 51492 4172 51884 4228
rect 51940 4172 51950 4228
rect 66546 4172 66556 4228
rect 66612 4172 70252 4228
rect 70308 4172 70318 4228
rect 107874 4172 107884 4228
rect 107940 4172 109452 4228
rect 109508 4172 109518 4228
rect 126354 4172 126364 4228
rect 126420 4172 132972 4228
rect 133028 4172 133308 4228
rect 133364 4172 133374 4228
rect 133858 4172 133868 4228
rect 133924 4172 134428 4228
rect 134484 4172 134494 4228
rect 14914 4060 14924 4116
rect 14980 4060 16492 4116
rect 16548 4060 16558 4116
rect 25666 4060 25676 4116
rect 25732 4060 27244 4116
rect 27300 4060 27310 4116
rect 29138 4060 29148 4116
rect 29204 4060 56364 4116
rect 56420 4060 56430 4116
rect 113362 4060 113372 4116
rect 113428 4060 114828 4116
rect 114884 4060 114894 4116
rect 117058 3948 117068 4004
rect 117124 3948 118300 4004
rect 118356 3948 119308 4004
rect 119364 3948 129276 4004
rect 129332 3948 129342 4004
rect 19612 3892 19622 3948
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19886 3892 19896 3948
rect 56432 3892 56442 3948
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56706 3892 56716 3948
rect 93252 3892 93262 3948
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93526 3892 93536 3948
rect 130072 3892 130082 3948
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130346 3892 130356 3948
rect 8530 3836 8540 3892
rect 8596 3836 8988 3892
rect 9044 3836 9772 3892
rect 9828 3836 17612 3892
rect 17668 3836 17678 3892
rect 102732 3836 108780 3892
rect 108836 3836 110124 3892
rect 110180 3836 110190 3892
rect 102732 3780 102788 3836
rect 10434 3724 10444 3780
rect 10500 3724 12236 3780
rect 12292 3724 12302 3780
rect 55122 3724 55132 3780
rect 55188 3724 57596 3780
rect 57652 3724 57662 3780
rect 58716 3724 63532 3780
rect 63588 3724 63598 3780
rect 78932 3724 89852 3780
rect 89908 3724 89918 3780
rect 101266 3724 101276 3780
rect 101332 3724 102732 3780
rect 102788 3724 102798 3780
rect 107426 3724 107436 3780
rect 107492 3724 108108 3780
rect 108164 3724 108174 3780
rect 125682 3724 125692 3780
rect 125748 3724 127260 3780
rect 127316 3724 127326 3780
rect 129490 3724 129500 3780
rect 129556 3724 131628 3780
rect 131684 3724 132300 3780
rect 132356 3724 132366 3780
rect 58716 3668 58772 3724
rect 78932 3668 78988 3724
rect 8306 3612 8316 3668
rect 8372 3612 8764 3668
rect 8820 3612 9996 3668
rect 10052 3612 10062 3668
rect 20132 3612 20412 3668
rect 20468 3612 20478 3668
rect 54002 3612 54012 3668
rect 54068 3612 58772 3668
rect 58930 3612 58940 3668
rect 58996 3612 60844 3668
rect 60900 3612 60910 3668
rect 63644 3612 66556 3668
rect 66612 3612 66622 3668
rect 75618 3612 75628 3668
rect 75684 3612 77532 3668
rect 77588 3612 78988 3668
rect 85362 3612 85372 3668
rect 85428 3612 86268 3668
rect 86324 3612 86334 3668
rect 93202 3612 93212 3668
rect 93268 3612 94668 3668
rect 94724 3612 103068 3668
rect 103124 3612 103134 3668
rect 115714 3612 115724 3668
rect 115780 3612 117180 3668
rect 117236 3612 117246 3668
rect 121426 3612 121436 3668
rect 121492 3612 123340 3668
rect 123396 3612 132636 3668
rect 132692 3612 132702 3668
rect 5842 3500 5852 3556
rect 5908 3500 7308 3556
rect 7364 3500 8428 3556
rect 8484 3500 8494 3556
rect 20132 3444 20188 3612
rect 63644 3556 63700 3612
rect 40674 3500 40684 3556
rect 40740 3500 41244 3556
rect 41300 3500 41310 3556
rect 44146 3500 44156 3556
rect 44212 3500 45052 3556
rect 45108 3500 45118 3556
rect 51986 3500 51996 3556
rect 52052 3500 52332 3556
rect 52388 3500 52780 3556
rect 52836 3500 52846 3556
rect 53778 3500 53788 3556
rect 53844 3500 55916 3556
rect 55972 3500 59836 3556
rect 59892 3500 62412 3556
rect 62468 3500 62478 3556
rect 62738 3500 62748 3556
rect 62804 3500 63644 3556
rect 63700 3500 63710 3556
rect 64978 3500 64988 3556
rect 65044 3500 67564 3556
rect 67620 3500 70588 3556
rect 70644 3500 70654 3556
rect 71698 3500 71708 3556
rect 71764 3500 73612 3556
rect 73668 3500 76300 3556
rect 76356 3500 76366 3556
rect 81442 3500 81452 3556
rect 81508 3500 82908 3556
rect 82964 3500 82974 3556
rect 97234 3500 97244 3556
rect 97300 3500 98700 3556
rect 98756 3500 102956 3556
rect 103012 3500 103022 3556
rect 105298 3500 105308 3556
rect 105364 3500 109004 3556
rect 109060 3500 109070 3556
rect 109218 3500 109228 3556
rect 109284 3500 110684 3556
rect 110740 3500 110750 3556
rect 125346 3500 125356 3556
rect 125412 3500 126140 3556
rect 126196 3500 131068 3556
rect 131124 3500 131134 3556
rect 6290 3388 6300 3444
rect 6356 3388 6524 3444
rect 6580 3388 7084 3444
rect 7140 3388 7150 3444
rect 9762 3388 9772 3444
rect 9828 3388 10108 3444
rect 10164 3388 10332 3444
rect 10388 3388 10398 3444
rect 11106 3388 11116 3444
rect 11172 3388 11676 3444
rect 11732 3388 11742 3444
rect 13794 3388 13804 3444
rect 13860 3388 14364 3444
rect 14420 3388 14430 3444
rect 15922 3388 15932 3444
rect 15988 3388 18844 3444
rect 18900 3388 20188 3444
rect 24546 3388 24556 3444
rect 24612 3388 25676 3444
rect 25732 3388 25742 3444
rect 28578 3388 28588 3444
rect 28644 3388 29596 3444
rect 29652 3388 29662 3444
rect 29922 3388 29932 3444
rect 29988 3388 30492 3444
rect 30548 3388 30558 3444
rect 31266 3388 31276 3444
rect 31332 3388 31836 3444
rect 31892 3388 31902 3444
rect 32610 3388 32620 3444
rect 32676 3388 32956 3444
rect 33012 3388 33180 3444
rect 33236 3388 33246 3444
rect 51202 3388 51212 3444
rect 51268 3388 53340 3444
rect 53396 3388 54124 3444
rect 54180 3388 54190 3444
rect 55458 3388 55468 3444
rect 55524 3388 57036 3444
rect 57092 3388 57102 3444
rect 59602 3388 59612 3444
rect 59668 3388 60956 3444
rect 61012 3388 61022 3444
rect 63522 3388 63532 3444
rect 63588 3388 64876 3444
rect 64932 3388 64942 3444
rect 67666 3388 67676 3444
rect 67732 3388 68796 3444
rect 68852 3388 68862 3444
rect 71586 3388 71596 3444
rect 71652 3388 72716 3444
rect 72772 3388 72782 3444
rect 72930 3388 72940 3444
rect 72996 3388 74508 3444
rect 74564 3388 74956 3444
rect 75012 3388 75022 3444
rect 75618 3388 75628 3444
rect 75684 3388 76636 3444
rect 76692 3388 76702 3444
rect 76962 3388 76972 3444
rect 77028 3388 78428 3444
rect 78484 3388 79324 3444
rect 79380 3388 79390 3444
rect 79650 3388 79660 3444
rect 79716 3388 80556 3444
rect 80612 3388 80622 3444
rect 80994 3388 81004 3444
rect 81060 3388 81788 3444
rect 81844 3388 82012 3444
rect 82068 3388 82078 3444
rect 83682 3388 83692 3444
rect 83748 3388 84476 3444
rect 84532 3388 84542 3444
rect 85026 3388 85036 3444
rect 85092 3388 86268 3444
rect 86324 3388 86716 3444
rect 86772 3388 86782 3444
rect 87714 3388 87724 3444
rect 87780 3388 88396 3444
rect 88452 3388 88462 3444
rect 89170 3388 89180 3444
rect 89236 3388 90188 3444
rect 90244 3388 90636 3444
rect 90692 3388 90702 3444
rect 91746 3388 91756 3444
rect 91812 3388 92316 3444
rect 92372 3388 92382 3444
rect 93090 3388 93100 3444
rect 93156 3388 93772 3444
rect 93828 3388 93838 3444
rect 95778 3388 95788 3444
rect 95844 3388 96348 3444
rect 96404 3388 96414 3444
rect 97122 3388 97132 3444
rect 97188 3388 97580 3444
rect 97636 3388 97804 3444
rect 97860 3388 97870 3444
rect 99810 3388 99820 3444
rect 99876 3388 100380 3444
rect 100436 3388 100446 3444
rect 101154 3388 101164 3444
rect 101220 3388 101612 3444
rect 101668 3388 101836 3444
rect 101892 3388 101902 3444
rect 103842 3388 103852 3444
rect 103908 3388 104412 3444
rect 104468 3388 104478 3444
rect 105186 3388 105196 3444
rect 105252 3388 106204 3444
rect 106260 3388 106652 3444
rect 106708 3388 106718 3444
rect 109890 3388 109900 3444
rect 109956 3388 111468 3444
rect 111524 3388 111534 3444
rect 115938 3388 115948 3444
rect 116004 3388 116508 3444
rect 116564 3388 116574 3444
rect 119970 3388 119980 3444
rect 120036 3388 120540 3444
rect 120596 3388 120606 3444
rect 121314 3388 121324 3444
rect 121380 3388 121772 3444
rect 121828 3388 121996 3444
rect 122052 3388 122062 3444
rect 124002 3388 124012 3444
rect 124068 3388 124572 3444
rect 124628 3388 124638 3444
rect 128034 3388 128044 3444
rect 128100 3388 128604 3444
rect 128660 3388 128670 3444
rect 132066 3388 132076 3444
rect 132132 3388 132636 3444
rect 132692 3388 132702 3444
rect 136098 3388 136108 3444
rect 136164 3388 136668 3444
rect 136724 3388 136734 3444
rect 137442 3388 137452 3444
rect 137508 3388 138012 3444
rect 138068 3388 138078 3444
rect 140130 3388 140140 3444
rect 140196 3388 141260 3444
rect 141316 3388 141326 3444
rect 144162 3388 144172 3444
rect 144228 3388 145292 3444
rect 145348 3388 145358 3444
rect 6626 3276 6636 3332
rect 6692 3276 8652 3332
rect 8708 3276 8718 3332
rect 8866 3276 8876 3332
rect 8932 3276 11340 3332
rect 11396 3276 11406 3332
rect 15026 3276 15036 3332
rect 15092 3276 16716 3332
rect 16772 3276 16782 3332
rect 26226 3276 26236 3332
rect 26292 3276 29260 3332
rect 29316 3276 29326 3332
rect 39554 3276 39564 3332
rect 39620 3276 41020 3332
rect 41076 3276 41086 3332
rect 45938 3276 45948 3332
rect 46004 3276 49532 3332
rect 49588 3276 49598 3332
rect 89058 3276 89068 3332
rect 89124 3276 89852 3332
rect 89908 3276 89918 3332
rect 95554 3276 95564 3332
rect 95620 3276 102172 3332
rect 102228 3276 102238 3332
rect 11218 3164 11228 3220
rect 11284 3164 23772 3220
rect 23828 3164 23838 3220
rect 25106 3164 25116 3220
rect 25172 3164 32284 3220
rect 32340 3164 32350 3220
rect 43138 3164 43148 3220
rect 43204 3164 58604 3220
rect 58660 3164 58670 3220
rect 78194 3164 78204 3220
rect 78260 3164 83132 3220
rect 83188 3164 83198 3220
rect 94098 3164 94108 3220
rect 94164 3164 96460 3220
rect 96516 3164 96526 3220
rect 38022 3108 38032 3164
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38296 3108 38306 3164
rect 74842 3108 74852 3164
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 75116 3108 75126 3164
rect 111662 3108 111672 3164
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111936 3108 111946 3164
rect 148482 3108 148492 3164
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148756 3108 148766 3164
rect 7522 2940 7532 2996
rect 7588 2940 53788 2996
rect 53844 2940 53854 2996
rect 56914 2940 56924 2996
rect 56980 2940 59500 2996
rect 59556 2940 117068 2996
rect 117124 2940 117134 2996
rect 74162 2828 74172 2884
rect 74228 2828 101500 2884
rect 101556 2828 101566 2884
rect 58594 2716 58604 2772
rect 58660 2716 99932 2772
rect 99988 2716 99998 2772
rect 58370 2604 58380 2660
rect 58436 2604 94108 2660
rect 94164 2604 94174 2660
rect 89842 2492 89852 2548
rect 89908 2492 113260 2548
rect 113316 2492 113326 2548
rect 6402 28 6412 84
rect 6468 28 68572 84
rect 68628 28 68638 84
<< via3 >>
rect 19622 36820 19678 36876
rect 19726 36820 19782 36876
rect 19830 36820 19886 36876
rect 56442 36820 56498 36876
rect 56546 36820 56602 36876
rect 56650 36820 56706 36876
rect 93262 36820 93318 36876
rect 93366 36820 93422 36876
rect 93470 36820 93526 36876
rect 130082 36820 130138 36876
rect 130186 36820 130242 36876
rect 130290 36820 130346 36876
rect 38032 36036 38088 36092
rect 38136 36036 38192 36092
rect 38240 36036 38296 36092
rect 74852 36036 74908 36092
rect 74956 36036 75012 36092
rect 75060 36036 75116 36092
rect 111672 36036 111728 36092
rect 111776 36036 111832 36092
rect 111880 36036 111936 36092
rect 148492 36036 148548 36092
rect 148596 36036 148652 36092
rect 148700 36036 148756 36092
rect 78764 35644 78820 35700
rect 19622 35252 19678 35308
rect 19726 35252 19782 35308
rect 19830 35252 19886 35308
rect 56442 35252 56498 35308
rect 56546 35252 56602 35308
rect 56650 35252 56706 35308
rect 93262 35252 93318 35308
rect 93366 35252 93422 35308
rect 93470 35252 93526 35308
rect 130082 35252 130138 35308
rect 130186 35252 130242 35308
rect 130290 35252 130346 35308
rect 37772 35196 37828 35252
rect 61404 35196 61460 35252
rect 78204 35196 78260 35252
rect 61292 34972 61348 35028
rect 78316 34972 78372 35028
rect 107324 34972 107380 35028
rect 85708 34860 85764 34916
rect 107212 34748 107268 34804
rect 37772 34636 37828 34692
rect 78764 34636 78820 34692
rect 85708 34636 85764 34692
rect 38032 34468 38088 34524
rect 38136 34468 38192 34524
rect 38240 34468 38296 34524
rect 74852 34468 74908 34524
rect 74956 34468 75012 34524
rect 75060 34468 75116 34524
rect 111672 34468 111728 34524
rect 111776 34468 111832 34524
rect 111880 34468 111936 34524
rect 148492 34468 148548 34524
rect 148596 34468 148652 34524
rect 148700 34468 148756 34524
rect 56028 34412 56084 34468
rect 52108 33852 52164 33908
rect 56028 33852 56084 33908
rect 19622 33684 19678 33740
rect 19726 33684 19782 33740
rect 19830 33684 19886 33740
rect 56442 33684 56498 33740
rect 56546 33684 56602 33740
rect 56650 33684 56706 33740
rect 93262 33684 93318 33740
rect 93366 33684 93422 33740
rect 93470 33684 93526 33740
rect 130082 33684 130138 33740
rect 130186 33684 130242 33740
rect 130290 33684 130346 33740
rect 38032 32900 38088 32956
rect 38136 32900 38192 32956
rect 38240 32900 38296 32956
rect 74852 32900 74908 32956
rect 74956 32900 75012 32956
rect 75060 32900 75116 32956
rect 111672 32900 111728 32956
rect 111776 32900 111832 32956
rect 111880 32900 111936 32956
rect 148492 32900 148548 32956
rect 148596 32900 148652 32956
rect 148700 32900 148756 32956
rect 52108 32508 52164 32564
rect 19622 32116 19678 32172
rect 19726 32116 19782 32172
rect 19830 32116 19886 32172
rect 56442 32116 56498 32172
rect 56546 32116 56602 32172
rect 56650 32116 56706 32172
rect 93262 32116 93318 32172
rect 93366 32116 93422 32172
rect 93470 32116 93526 32172
rect 130082 32116 130138 32172
rect 130186 32116 130242 32172
rect 130290 32116 130346 32172
rect 38032 31332 38088 31388
rect 38136 31332 38192 31388
rect 38240 31332 38296 31388
rect 74852 31332 74908 31388
rect 74956 31332 75012 31388
rect 75060 31332 75116 31388
rect 111672 31332 111728 31388
rect 111776 31332 111832 31388
rect 111880 31332 111936 31388
rect 148492 31332 148548 31388
rect 148596 31332 148652 31388
rect 148700 31332 148756 31388
rect 19622 30548 19678 30604
rect 19726 30548 19782 30604
rect 19830 30548 19886 30604
rect 56442 30548 56498 30604
rect 56546 30548 56602 30604
rect 56650 30548 56706 30604
rect 93262 30548 93318 30604
rect 93366 30548 93422 30604
rect 93470 30548 93526 30604
rect 130082 30548 130138 30604
rect 130186 30548 130242 30604
rect 130290 30548 130346 30604
rect 38032 29764 38088 29820
rect 38136 29764 38192 29820
rect 38240 29764 38296 29820
rect 74852 29764 74908 29820
rect 74956 29764 75012 29820
rect 75060 29764 75116 29820
rect 111672 29764 111728 29820
rect 111776 29764 111832 29820
rect 111880 29764 111936 29820
rect 148492 29764 148548 29820
rect 148596 29764 148652 29820
rect 148700 29764 148756 29820
rect 19622 28980 19678 29036
rect 19726 28980 19782 29036
rect 19830 28980 19886 29036
rect 56442 28980 56498 29036
rect 56546 28980 56602 29036
rect 56650 28980 56706 29036
rect 93262 28980 93318 29036
rect 93366 28980 93422 29036
rect 93470 28980 93526 29036
rect 130082 28980 130138 29036
rect 130186 28980 130242 29036
rect 130290 28980 130346 29036
rect 38032 28196 38088 28252
rect 38136 28196 38192 28252
rect 38240 28196 38296 28252
rect 74852 28196 74908 28252
rect 74956 28196 75012 28252
rect 75060 28196 75116 28252
rect 111672 28196 111728 28252
rect 111776 28196 111832 28252
rect 111880 28196 111936 28252
rect 148492 28196 148548 28252
rect 148596 28196 148652 28252
rect 148700 28196 148756 28252
rect 19622 27412 19678 27468
rect 19726 27412 19782 27468
rect 19830 27412 19886 27468
rect 56442 27412 56498 27468
rect 56546 27412 56602 27468
rect 56650 27412 56706 27468
rect 93262 27412 93318 27468
rect 93366 27412 93422 27468
rect 93470 27412 93526 27468
rect 130082 27412 130138 27468
rect 130186 27412 130242 27468
rect 130290 27412 130346 27468
rect 38032 26628 38088 26684
rect 38136 26628 38192 26684
rect 38240 26628 38296 26684
rect 74852 26628 74908 26684
rect 74956 26628 75012 26684
rect 75060 26628 75116 26684
rect 111672 26628 111728 26684
rect 111776 26628 111832 26684
rect 111880 26628 111936 26684
rect 148492 26628 148548 26684
rect 148596 26628 148652 26684
rect 148700 26628 148756 26684
rect 19622 25844 19678 25900
rect 19726 25844 19782 25900
rect 19830 25844 19886 25900
rect 56442 25844 56498 25900
rect 56546 25844 56602 25900
rect 56650 25844 56706 25900
rect 93262 25844 93318 25900
rect 93366 25844 93422 25900
rect 93470 25844 93526 25900
rect 130082 25844 130138 25900
rect 130186 25844 130242 25900
rect 130290 25844 130346 25900
rect 38032 25060 38088 25116
rect 38136 25060 38192 25116
rect 38240 25060 38296 25116
rect 74852 25060 74908 25116
rect 74956 25060 75012 25116
rect 75060 25060 75116 25116
rect 111672 25060 111728 25116
rect 111776 25060 111832 25116
rect 111880 25060 111936 25116
rect 148492 25060 148548 25116
rect 148596 25060 148652 25116
rect 148700 25060 148756 25116
rect 19622 24276 19678 24332
rect 19726 24276 19782 24332
rect 19830 24276 19886 24332
rect 56442 24276 56498 24332
rect 56546 24276 56602 24332
rect 56650 24276 56706 24332
rect 93262 24276 93318 24332
rect 93366 24276 93422 24332
rect 93470 24276 93526 24332
rect 130082 24276 130138 24332
rect 130186 24276 130242 24332
rect 130290 24276 130346 24332
rect 38032 23492 38088 23548
rect 38136 23492 38192 23548
rect 38240 23492 38296 23548
rect 74852 23492 74908 23548
rect 74956 23492 75012 23548
rect 75060 23492 75116 23548
rect 111672 23492 111728 23548
rect 111776 23492 111832 23548
rect 111880 23492 111936 23548
rect 148492 23492 148548 23548
rect 148596 23492 148652 23548
rect 148700 23492 148756 23548
rect 19622 22708 19678 22764
rect 19726 22708 19782 22764
rect 19830 22708 19886 22764
rect 56442 22708 56498 22764
rect 56546 22708 56602 22764
rect 56650 22708 56706 22764
rect 93262 22708 93318 22764
rect 93366 22708 93422 22764
rect 93470 22708 93526 22764
rect 130082 22708 130138 22764
rect 130186 22708 130242 22764
rect 130290 22708 130346 22764
rect 38032 21924 38088 21980
rect 38136 21924 38192 21980
rect 38240 21924 38296 21980
rect 74852 21924 74908 21980
rect 74956 21924 75012 21980
rect 75060 21924 75116 21980
rect 111672 21924 111728 21980
rect 111776 21924 111832 21980
rect 111880 21924 111936 21980
rect 148492 21924 148548 21980
rect 148596 21924 148652 21980
rect 148700 21924 148756 21980
rect 19622 21140 19678 21196
rect 19726 21140 19782 21196
rect 19830 21140 19886 21196
rect 56442 21140 56498 21196
rect 56546 21140 56602 21196
rect 56650 21140 56706 21196
rect 93262 21140 93318 21196
rect 93366 21140 93422 21196
rect 93470 21140 93526 21196
rect 130082 21140 130138 21196
rect 130186 21140 130242 21196
rect 130290 21140 130346 21196
rect 38032 20356 38088 20412
rect 38136 20356 38192 20412
rect 38240 20356 38296 20412
rect 74852 20356 74908 20412
rect 74956 20356 75012 20412
rect 75060 20356 75116 20412
rect 111672 20356 111728 20412
rect 111776 20356 111832 20412
rect 111880 20356 111936 20412
rect 148492 20356 148548 20412
rect 148596 20356 148652 20412
rect 148700 20356 148756 20412
rect 19622 19572 19678 19628
rect 19726 19572 19782 19628
rect 19830 19572 19886 19628
rect 56442 19572 56498 19628
rect 56546 19572 56602 19628
rect 56650 19572 56706 19628
rect 93262 19572 93318 19628
rect 93366 19572 93422 19628
rect 93470 19572 93526 19628
rect 130082 19572 130138 19628
rect 130186 19572 130242 19628
rect 130290 19572 130346 19628
rect 38032 18788 38088 18844
rect 38136 18788 38192 18844
rect 38240 18788 38296 18844
rect 74852 18788 74908 18844
rect 74956 18788 75012 18844
rect 75060 18788 75116 18844
rect 111672 18788 111728 18844
rect 111776 18788 111832 18844
rect 111880 18788 111936 18844
rect 148492 18788 148548 18844
rect 148596 18788 148652 18844
rect 148700 18788 148756 18844
rect 19622 18004 19678 18060
rect 19726 18004 19782 18060
rect 19830 18004 19886 18060
rect 56442 18004 56498 18060
rect 56546 18004 56602 18060
rect 56650 18004 56706 18060
rect 93262 18004 93318 18060
rect 93366 18004 93422 18060
rect 93470 18004 93526 18060
rect 130082 18004 130138 18060
rect 130186 18004 130242 18060
rect 130290 18004 130346 18060
rect 38032 17220 38088 17276
rect 38136 17220 38192 17276
rect 38240 17220 38296 17276
rect 74852 17220 74908 17276
rect 74956 17220 75012 17276
rect 75060 17220 75116 17276
rect 111672 17220 111728 17276
rect 111776 17220 111832 17276
rect 111880 17220 111936 17276
rect 148492 17220 148548 17276
rect 148596 17220 148652 17276
rect 148700 17220 148756 17276
rect 19622 16436 19678 16492
rect 19726 16436 19782 16492
rect 19830 16436 19886 16492
rect 56442 16436 56498 16492
rect 56546 16436 56602 16492
rect 56650 16436 56706 16492
rect 93262 16436 93318 16492
rect 93366 16436 93422 16492
rect 93470 16436 93526 16492
rect 130082 16436 130138 16492
rect 130186 16436 130242 16492
rect 130290 16436 130346 16492
rect 38032 15652 38088 15708
rect 38136 15652 38192 15708
rect 38240 15652 38296 15708
rect 74852 15652 74908 15708
rect 74956 15652 75012 15708
rect 75060 15652 75116 15708
rect 111672 15652 111728 15708
rect 111776 15652 111832 15708
rect 111880 15652 111936 15708
rect 148492 15652 148548 15708
rect 148596 15652 148652 15708
rect 148700 15652 148756 15708
rect 19622 14868 19678 14924
rect 19726 14868 19782 14924
rect 19830 14868 19886 14924
rect 56442 14868 56498 14924
rect 56546 14868 56602 14924
rect 56650 14868 56706 14924
rect 93262 14868 93318 14924
rect 93366 14868 93422 14924
rect 93470 14868 93526 14924
rect 130082 14868 130138 14924
rect 130186 14868 130242 14924
rect 130290 14868 130346 14924
rect 38032 14084 38088 14140
rect 38136 14084 38192 14140
rect 38240 14084 38296 14140
rect 74852 14084 74908 14140
rect 74956 14084 75012 14140
rect 75060 14084 75116 14140
rect 111672 14084 111728 14140
rect 111776 14084 111832 14140
rect 111880 14084 111936 14140
rect 148492 14084 148548 14140
rect 148596 14084 148652 14140
rect 148700 14084 148756 14140
rect 19622 13300 19678 13356
rect 19726 13300 19782 13356
rect 19830 13300 19886 13356
rect 56442 13300 56498 13356
rect 56546 13300 56602 13356
rect 56650 13300 56706 13356
rect 93262 13300 93318 13356
rect 93366 13300 93422 13356
rect 93470 13300 93526 13356
rect 130082 13300 130138 13356
rect 130186 13300 130242 13356
rect 130290 13300 130346 13356
rect 38032 12516 38088 12572
rect 38136 12516 38192 12572
rect 38240 12516 38296 12572
rect 74852 12516 74908 12572
rect 74956 12516 75012 12572
rect 75060 12516 75116 12572
rect 111672 12516 111728 12572
rect 111776 12516 111832 12572
rect 111880 12516 111936 12572
rect 148492 12516 148548 12572
rect 148596 12516 148652 12572
rect 148700 12516 148756 12572
rect 19622 11732 19678 11788
rect 19726 11732 19782 11788
rect 19830 11732 19886 11788
rect 56442 11732 56498 11788
rect 56546 11732 56602 11788
rect 56650 11732 56706 11788
rect 93262 11732 93318 11788
rect 93366 11732 93422 11788
rect 93470 11732 93526 11788
rect 130082 11732 130138 11788
rect 130186 11732 130242 11788
rect 130290 11732 130346 11788
rect 38032 10948 38088 11004
rect 38136 10948 38192 11004
rect 38240 10948 38296 11004
rect 74852 10948 74908 11004
rect 74956 10948 75012 11004
rect 75060 10948 75116 11004
rect 111672 10948 111728 11004
rect 111776 10948 111832 11004
rect 111880 10948 111936 11004
rect 148492 10948 148548 11004
rect 148596 10948 148652 11004
rect 148700 10948 148756 11004
rect 19622 10164 19678 10220
rect 19726 10164 19782 10220
rect 19830 10164 19886 10220
rect 56442 10164 56498 10220
rect 56546 10164 56602 10220
rect 56650 10164 56706 10220
rect 93262 10164 93318 10220
rect 93366 10164 93422 10220
rect 93470 10164 93526 10220
rect 130082 10164 130138 10220
rect 130186 10164 130242 10220
rect 130290 10164 130346 10220
rect 38032 9380 38088 9436
rect 38136 9380 38192 9436
rect 38240 9380 38296 9436
rect 74852 9380 74908 9436
rect 74956 9380 75012 9436
rect 75060 9380 75116 9436
rect 111672 9380 111728 9436
rect 111776 9380 111832 9436
rect 111880 9380 111936 9436
rect 148492 9380 148548 9436
rect 148596 9380 148652 9436
rect 148700 9380 148756 9436
rect 19622 8596 19678 8652
rect 19726 8596 19782 8652
rect 19830 8596 19886 8652
rect 56442 8596 56498 8652
rect 56546 8596 56602 8652
rect 56650 8596 56706 8652
rect 93262 8596 93318 8652
rect 93366 8596 93422 8652
rect 93470 8596 93526 8652
rect 130082 8596 130138 8652
rect 130186 8596 130242 8652
rect 130290 8596 130346 8652
rect 38032 7812 38088 7868
rect 38136 7812 38192 7868
rect 38240 7812 38296 7868
rect 74852 7812 74908 7868
rect 74956 7812 75012 7868
rect 75060 7812 75116 7868
rect 111672 7812 111728 7868
rect 111776 7812 111832 7868
rect 111880 7812 111936 7868
rect 148492 7812 148548 7868
rect 148596 7812 148652 7868
rect 148700 7812 148756 7868
rect 19622 7028 19678 7084
rect 19726 7028 19782 7084
rect 19830 7028 19886 7084
rect 56442 7028 56498 7084
rect 56546 7028 56602 7084
rect 56650 7028 56706 7084
rect 93262 7028 93318 7084
rect 93366 7028 93422 7084
rect 93470 7028 93526 7084
rect 130082 7028 130138 7084
rect 130186 7028 130242 7084
rect 130290 7028 130346 7084
rect 38032 6244 38088 6300
rect 38136 6244 38192 6300
rect 38240 6244 38296 6300
rect 74852 6244 74908 6300
rect 74956 6244 75012 6300
rect 75060 6244 75116 6300
rect 111672 6244 111728 6300
rect 111776 6244 111832 6300
rect 111880 6244 111936 6300
rect 148492 6244 148548 6300
rect 148596 6244 148652 6300
rect 148700 6244 148756 6300
rect 134204 5516 134260 5572
rect 19622 5460 19678 5516
rect 19726 5460 19782 5516
rect 19830 5460 19886 5516
rect 56442 5460 56498 5516
rect 56546 5460 56602 5516
rect 56650 5460 56706 5516
rect 93262 5460 93318 5516
rect 93366 5460 93422 5516
rect 93470 5460 93526 5516
rect 130082 5460 130138 5516
rect 130186 5460 130242 5516
rect 130290 5460 130346 5516
rect 134204 5068 134260 5124
rect 38032 4676 38088 4732
rect 38136 4676 38192 4732
rect 38240 4676 38296 4732
rect 74852 4676 74908 4732
rect 74956 4676 75012 4732
rect 75060 4676 75116 4732
rect 111672 4676 111728 4732
rect 111776 4676 111832 4732
rect 111880 4676 111936 4732
rect 148492 4676 148548 4732
rect 148596 4676 148652 4732
rect 148700 4676 148756 4732
rect 19622 3892 19678 3948
rect 19726 3892 19782 3948
rect 19830 3892 19886 3948
rect 56442 3892 56498 3948
rect 56546 3892 56602 3948
rect 56650 3892 56706 3948
rect 93262 3892 93318 3948
rect 93366 3892 93422 3948
rect 93470 3892 93526 3948
rect 130082 3892 130138 3948
rect 130186 3892 130242 3948
rect 130290 3892 130346 3948
rect 38032 3108 38088 3164
rect 38136 3108 38192 3164
rect 38240 3108 38296 3164
rect 74852 3108 74908 3164
rect 74956 3108 75012 3164
rect 75060 3108 75116 3164
rect 111672 3108 111728 3164
rect 111776 3108 111832 3164
rect 111880 3108 111936 3164
rect 148492 3108 148548 3164
rect 148596 3108 148652 3164
rect 148700 3108 148756 3164
<< metal4 >>
rect 19594 36876 19914 36908
rect 19594 36820 19622 36876
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19886 36820 19914 36876
rect 19594 35308 19914 36820
rect 19594 35252 19622 35308
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19886 35252 19914 35308
rect 38004 36092 38324 36908
rect 38004 36036 38032 36092
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38296 36036 38324 36092
rect 19594 33740 19914 35252
rect 37772 35252 37828 35262
rect 37772 34692 37828 35196
rect 37772 34626 37828 34636
rect 19594 33684 19622 33740
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19886 33684 19914 33740
rect 19594 32172 19914 33684
rect 19594 32116 19622 32172
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19886 32116 19914 32172
rect 19594 30604 19914 32116
rect 19594 30548 19622 30604
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19886 30548 19914 30604
rect 19594 29036 19914 30548
rect 19594 28980 19622 29036
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19886 28980 19914 29036
rect 19594 27468 19914 28980
rect 19594 27412 19622 27468
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19886 27412 19914 27468
rect 19594 25900 19914 27412
rect 19594 25844 19622 25900
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19886 25844 19914 25900
rect 19594 24332 19914 25844
rect 19594 24276 19622 24332
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19886 24276 19914 24332
rect 19594 22764 19914 24276
rect 19594 22708 19622 22764
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19886 22708 19914 22764
rect 19594 21196 19914 22708
rect 19594 21140 19622 21196
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19886 21140 19914 21196
rect 19594 19628 19914 21140
rect 19594 19572 19622 19628
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19886 19572 19914 19628
rect 19594 18060 19914 19572
rect 19594 18004 19622 18060
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19886 18004 19914 18060
rect 19594 16492 19914 18004
rect 19594 16436 19622 16492
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19886 16436 19914 16492
rect 19594 14924 19914 16436
rect 19594 14868 19622 14924
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19886 14868 19914 14924
rect 19594 13356 19914 14868
rect 19594 13300 19622 13356
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19886 13300 19914 13356
rect 19594 11788 19914 13300
rect 19594 11732 19622 11788
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19886 11732 19914 11788
rect 19594 10220 19914 11732
rect 19594 10164 19622 10220
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19886 10164 19914 10220
rect 19594 8652 19914 10164
rect 19594 8596 19622 8652
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19886 8596 19914 8652
rect 19594 7084 19914 8596
rect 19594 7028 19622 7084
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19886 7028 19914 7084
rect 19594 5516 19914 7028
rect 19594 5460 19622 5516
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19886 5460 19914 5516
rect 19594 3948 19914 5460
rect 19594 3892 19622 3948
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19886 3892 19914 3948
rect 19594 3076 19914 3892
rect 38004 34524 38324 36036
rect 38004 34468 38032 34524
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38296 34468 38324 34524
rect 56414 36876 56734 36908
rect 56414 36820 56442 36876
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56706 36820 56734 36876
rect 56414 35308 56734 36820
rect 56414 35252 56442 35308
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56706 35252 56734 35308
rect 74824 36092 75144 36908
rect 74824 36036 74852 36092
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 75116 36036 75144 36092
rect 38004 32956 38324 34468
rect 56028 34468 56084 34478
rect 38004 32900 38032 32956
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38296 32900 38324 32956
rect 38004 31388 38324 32900
rect 52108 33908 52164 33918
rect 52108 32564 52164 33852
rect 56028 33908 56084 34412
rect 56028 33842 56084 33852
rect 52108 32498 52164 32508
rect 56414 33740 56734 35252
rect 61404 35252 61460 35262
rect 61292 35028 61348 35038
rect 61404 35028 61460 35196
rect 61348 34972 61460 35028
rect 61292 34962 61348 34972
rect 56414 33684 56442 33740
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56706 33684 56734 33740
rect 38004 31332 38032 31388
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38296 31332 38324 31388
rect 38004 29820 38324 31332
rect 38004 29764 38032 29820
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38296 29764 38324 29820
rect 38004 28252 38324 29764
rect 38004 28196 38032 28252
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38296 28196 38324 28252
rect 38004 26684 38324 28196
rect 38004 26628 38032 26684
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38296 26628 38324 26684
rect 38004 25116 38324 26628
rect 38004 25060 38032 25116
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38296 25060 38324 25116
rect 38004 23548 38324 25060
rect 38004 23492 38032 23548
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38296 23492 38324 23548
rect 38004 21980 38324 23492
rect 38004 21924 38032 21980
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38296 21924 38324 21980
rect 38004 20412 38324 21924
rect 38004 20356 38032 20412
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38296 20356 38324 20412
rect 38004 18844 38324 20356
rect 38004 18788 38032 18844
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38296 18788 38324 18844
rect 38004 17276 38324 18788
rect 38004 17220 38032 17276
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38296 17220 38324 17276
rect 38004 15708 38324 17220
rect 38004 15652 38032 15708
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38296 15652 38324 15708
rect 38004 14140 38324 15652
rect 38004 14084 38032 14140
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38296 14084 38324 14140
rect 38004 12572 38324 14084
rect 38004 12516 38032 12572
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38296 12516 38324 12572
rect 38004 11004 38324 12516
rect 38004 10948 38032 11004
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38296 10948 38324 11004
rect 38004 9436 38324 10948
rect 38004 9380 38032 9436
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38296 9380 38324 9436
rect 38004 7868 38324 9380
rect 38004 7812 38032 7868
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38296 7812 38324 7868
rect 38004 6300 38324 7812
rect 38004 6244 38032 6300
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38296 6244 38324 6300
rect 38004 4732 38324 6244
rect 38004 4676 38032 4732
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38296 4676 38324 4732
rect 38004 3164 38324 4676
rect 38004 3108 38032 3164
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38296 3108 38324 3164
rect 38004 3076 38324 3108
rect 56414 32172 56734 33684
rect 56414 32116 56442 32172
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56706 32116 56734 32172
rect 56414 30604 56734 32116
rect 56414 30548 56442 30604
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56706 30548 56734 30604
rect 56414 29036 56734 30548
rect 56414 28980 56442 29036
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56706 28980 56734 29036
rect 56414 27468 56734 28980
rect 56414 27412 56442 27468
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56706 27412 56734 27468
rect 56414 25900 56734 27412
rect 56414 25844 56442 25900
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56706 25844 56734 25900
rect 56414 24332 56734 25844
rect 56414 24276 56442 24332
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56706 24276 56734 24332
rect 56414 22764 56734 24276
rect 56414 22708 56442 22764
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56706 22708 56734 22764
rect 56414 21196 56734 22708
rect 56414 21140 56442 21196
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56706 21140 56734 21196
rect 56414 19628 56734 21140
rect 56414 19572 56442 19628
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56706 19572 56734 19628
rect 56414 18060 56734 19572
rect 56414 18004 56442 18060
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56706 18004 56734 18060
rect 56414 16492 56734 18004
rect 56414 16436 56442 16492
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56706 16436 56734 16492
rect 56414 14924 56734 16436
rect 56414 14868 56442 14924
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56706 14868 56734 14924
rect 56414 13356 56734 14868
rect 56414 13300 56442 13356
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56706 13300 56734 13356
rect 56414 11788 56734 13300
rect 56414 11732 56442 11788
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56706 11732 56734 11788
rect 56414 10220 56734 11732
rect 56414 10164 56442 10220
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56706 10164 56734 10220
rect 56414 8652 56734 10164
rect 56414 8596 56442 8652
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56706 8596 56734 8652
rect 56414 7084 56734 8596
rect 56414 7028 56442 7084
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56706 7028 56734 7084
rect 56414 5516 56734 7028
rect 56414 5460 56442 5516
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56706 5460 56734 5516
rect 56414 3948 56734 5460
rect 56414 3892 56442 3948
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56706 3892 56734 3948
rect 56414 3076 56734 3892
rect 74824 34524 75144 36036
rect 93234 36876 93554 36908
rect 93234 36820 93262 36876
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93526 36820 93554 36876
rect 78764 35700 78820 35710
rect 78204 35252 78260 35262
rect 78260 35196 78372 35252
rect 78204 35186 78260 35196
rect 78316 35028 78372 35196
rect 78316 34962 78372 34972
rect 78764 34692 78820 35644
rect 93234 35308 93554 36820
rect 93234 35252 93262 35308
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93526 35252 93554 35308
rect 78764 34626 78820 34636
rect 85708 34916 85764 34926
rect 85708 34692 85764 34860
rect 85708 34626 85764 34636
rect 74824 34468 74852 34524
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 75116 34468 75144 34524
rect 74824 32956 75144 34468
rect 74824 32900 74852 32956
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 75116 32900 75144 32956
rect 74824 31388 75144 32900
rect 74824 31332 74852 31388
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 75116 31332 75144 31388
rect 74824 29820 75144 31332
rect 74824 29764 74852 29820
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 75116 29764 75144 29820
rect 74824 28252 75144 29764
rect 74824 28196 74852 28252
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 75116 28196 75144 28252
rect 74824 26684 75144 28196
rect 74824 26628 74852 26684
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 75116 26628 75144 26684
rect 74824 25116 75144 26628
rect 74824 25060 74852 25116
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 75116 25060 75144 25116
rect 74824 23548 75144 25060
rect 74824 23492 74852 23548
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 75116 23492 75144 23548
rect 74824 21980 75144 23492
rect 74824 21924 74852 21980
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 75116 21924 75144 21980
rect 74824 20412 75144 21924
rect 74824 20356 74852 20412
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 75116 20356 75144 20412
rect 74824 18844 75144 20356
rect 74824 18788 74852 18844
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 75116 18788 75144 18844
rect 74824 17276 75144 18788
rect 74824 17220 74852 17276
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 75116 17220 75144 17276
rect 74824 15708 75144 17220
rect 74824 15652 74852 15708
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 75116 15652 75144 15708
rect 74824 14140 75144 15652
rect 74824 14084 74852 14140
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 75116 14084 75144 14140
rect 74824 12572 75144 14084
rect 74824 12516 74852 12572
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 75116 12516 75144 12572
rect 74824 11004 75144 12516
rect 74824 10948 74852 11004
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 75116 10948 75144 11004
rect 74824 9436 75144 10948
rect 74824 9380 74852 9436
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 75116 9380 75144 9436
rect 74824 7868 75144 9380
rect 74824 7812 74852 7868
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 75116 7812 75144 7868
rect 74824 6300 75144 7812
rect 74824 6244 74852 6300
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 75116 6244 75144 6300
rect 74824 4732 75144 6244
rect 74824 4676 74852 4732
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 75116 4676 75144 4732
rect 74824 3164 75144 4676
rect 74824 3108 74852 3164
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 75116 3108 75144 3164
rect 74824 3076 75144 3108
rect 93234 33740 93554 35252
rect 111644 36092 111964 36908
rect 111644 36036 111672 36092
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111936 36036 111964 36092
rect 107324 35028 107380 35038
rect 107212 34972 107324 35028
rect 107212 34804 107268 34972
rect 107324 34962 107380 34972
rect 107212 34738 107268 34748
rect 93234 33684 93262 33740
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93526 33684 93554 33740
rect 93234 32172 93554 33684
rect 93234 32116 93262 32172
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93526 32116 93554 32172
rect 93234 30604 93554 32116
rect 93234 30548 93262 30604
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93526 30548 93554 30604
rect 93234 29036 93554 30548
rect 93234 28980 93262 29036
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93526 28980 93554 29036
rect 93234 27468 93554 28980
rect 93234 27412 93262 27468
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93526 27412 93554 27468
rect 93234 25900 93554 27412
rect 93234 25844 93262 25900
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93526 25844 93554 25900
rect 93234 24332 93554 25844
rect 93234 24276 93262 24332
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93526 24276 93554 24332
rect 93234 22764 93554 24276
rect 93234 22708 93262 22764
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93526 22708 93554 22764
rect 93234 21196 93554 22708
rect 93234 21140 93262 21196
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93526 21140 93554 21196
rect 93234 19628 93554 21140
rect 93234 19572 93262 19628
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93526 19572 93554 19628
rect 93234 18060 93554 19572
rect 93234 18004 93262 18060
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93526 18004 93554 18060
rect 93234 16492 93554 18004
rect 93234 16436 93262 16492
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93526 16436 93554 16492
rect 93234 14924 93554 16436
rect 93234 14868 93262 14924
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93526 14868 93554 14924
rect 93234 13356 93554 14868
rect 93234 13300 93262 13356
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93526 13300 93554 13356
rect 93234 11788 93554 13300
rect 93234 11732 93262 11788
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93526 11732 93554 11788
rect 93234 10220 93554 11732
rect 93234 10164 93262 10220
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93526 10164 93554 10220
rect 93234 8652 93554 10164
rect 93234 8596 93262 8652
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93526 8596 93554 8652
rect 93234 7084 93554 8596
rect 93234 7028 93262 7084
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93526 7028 93554 7084
rect 93234 5516 93554 7028
rect 93234 5460 93262 5516
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93526 5460 93554 5516
rect 93234 3948 93554 5460
rect 93234 3892 93262 3948
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93526 3892 93554 3948
rect 93234 3076 93554 3892
rect 111644 34524 111964 36036
rect 111644 34468 111672 34524
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111936 34468 111964 34524
rect 111644 32956 111964 34468
rect 111644 32900 111672 32956
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111936 32900 111964 32956
rect 111644 31388 111964 32900
rect 111644 31332 111672 31388
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111936 31332 111964 31388
rect 111644 29820 111964 31332
rect 111644 29764 111672 29820
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111936 29764 111964 29820
rect 111644 28252 111964 29764
rect 111644 28196 111672 28252
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111936 28196 111964 28252
rect 111644 26684 111964 28196
rect 111644 26628 111672 26684
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111936 26628 111964 26684
rect 111644 25116 111964 26628
rect 111644 25060 111672 25116
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111936 25060 111964 25116
rect 111644 23548 111964 25060
rect 111644 23492 111672 23548
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111936 23492 111964 23548
rect 111644 21980 111964 23492
rect 111644 21924 111672 21980
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111936 21924 111964 21980
rect 111644 20412 111964 21924
rect 111644 20356 111672 20412
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111936 20356 111964 20412
rect 111644 18844 111964 20356
rect 111644 18788 111672 18844
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111936 18788 111964 18844
rect 111644 17276 111964 18788
rect 111644 17220 111672 17276
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111936 17220 111964 17276
rect 111644 15708 111964 17220
rect 111644 15652 111672 15708
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111936 15652 111964 15708
rect 111644 14140 111964 15652
rect 111644 14084 111672 14140
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111936 14084 111964 14140
rect 111644 12572 111964 14084
rect 111644 12516 111672 12572
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111936 12516 111964 12572
rect 111644 11004 111964 12516
rect 111644 10948 111672 11004
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111936 10948 111964 11004
rect 111644 9436 111964 10948
rect 111644 9380 111672 9436
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111936 9380 111964 9436
rect 111644 7868 111964 9380
rect 111644 7812 111672 7868
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111936 7812 111964 7868
rect 111644 6300 111964 7812
rect 111644 6244 111672 6300
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111936 6244 111964 6300
rect 111644 4732 111964 6244
rect 111644 4676 111672 4732
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111936 4676 111964 4732
rect 111644 3164 111964 4676
rect 111644 3108 111672 3164
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111936 3108 111964 3164
rect 111644 3076 111964 3108
rect 130054 36876 130374 36908
rect 130054 36820 130082 36876
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130346 36820 130374 36876
rect 130054 35308 130374 36820
rect 130054 35252 130082 35308
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130346 35252 130374 35308
rect 130054 33740 130374 35252
rect 130054 33684 130082 33740
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130346 33684 130374 33740
rect 130054 32172 130374 33684
rect 130054 32116 130082 32172
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130346 32116 130374 32172
rect 130054 30604 130374 32116
rect 130054 30548 130082 30604
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130346 30548 130374 30604
rect 130054 29036 130374 30548
rect 130054 28980 130082 29036
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130346 28980 130374 29036
rect 130054 27468 130374 28980
rect 130054 27412 130082 27468
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130346 27412 130374 27468
rect 130054 25900 130374 27412
rect 130054 25844 130082 25900
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130346 25844 130374 25900
rect 130054 24332 130374 25844
rect 130054 24276 130082 24332
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130346 24276 130374 24332
rect 130054 22764 130374 24276
rect 130054 22708 130082 22764
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130346 22708 130374 22764
rect 130054 21196 130374 22708
rect 130054 21140 130082 21196
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130346 21140 130374 21196
rect 130054 19628 130374 21140
rect 130054 19572 130082 19628
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130346 19572 130374 19628
rect 130054 18060 130374 19572
rect 130054 18004 130082 18060
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130346 18004 130374 18060
rect 130054 16492 130374 18004
rect 130054 16436 130082 16492
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130346 16436 130374 16492
rect 130054 14924 130374 16436
rect 130054 14868 130082 14924
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130346 14868 130374 14924
rect 130054 13356 130374 14868
rect 130054 13300 130082 13356
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130346 13300 130374 13356
rect 130054 11788 130374 13300
rect 130054 11732 130082 11788
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130346 11732 130374 11788
rect 130054 10220 130374 11732
rect 130054 10164 130082 10220
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130346 10164 130374 10220
rect 130054 8652 130374 10164
rect 130054 8596 130082 8652
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130346 8596 130374 8652
rect 130054 7084 130374 8596
rect 130054 7028 130082 7084
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130346 7028 130374 7084
rect 130054 5516 130374 7028
rect 148464 36092 148784 36908
rect 148464 36036 148492 36092
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148756 36036 148784 36092
rect 148464 34524 148784 36036
rect 148464 34468 148492 34524
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148756 34468 148784 34524
rect 148464 32956 148784 34468
rect 148464 32900 148492 32956
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148756 32900 148784 32956
rect 148464 31388 148784 32900
rect 148464 31332 148492 31388
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148756 31332 148784 31388
rect 148464 29820 148784 31332
rect 148464 29764 148492 29820
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148756 29764 148784 29820
rect 148464 28252 148784 29764
rect 148464 28196 148492 28252
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148756 28196 148784 28252
rect 148464 26684 148784 28196
rect 148464 26628 148492 26684
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148756 26628 148784 26684
rect 148464 25116 148784 26628
rect 148464 25060 148492 25116
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148756 25060 148784 25116
rect 148464 23548 148784 25060
rect 148464 23492 148492 23548
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148756 23492 148784 23548
rect 148464 21980 148784 23492
rect 148464 21924 148492 21980
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148756 21924 148784 21980
rect 148464 20412 148784 21924
rect 148464 20356 148492 20412
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148756 20356 148784 20412
rect 148464 18844 148784 20356
rect 148464 18788 148492 18844
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148756 18788 148784 18844
rect 148464 17276 148784 18788
rect 148464 17220 148492 17276
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148756 17220 148784 17276
rect 148464 15708 148784 17220
rect 148464 15652 148492 15708
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148756 15652 148784 15708
rect 148464 14140 148784 15652
rect 148464 14084 148492 14140
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148756 14084 148784 14140
rect 148464 12572 148784 14084
rect 148464 12516 148492 12572
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148756 12516 148784 12572
rect 148464 11004 148784 12516
rect 148464 10948 148492 11004
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148756 10948 148784 11004
rect 148464 9436 148784 10948
rect 148464 9380 148492 9436
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148756 9380 148784 9436
rect 148464 7868 148784 9380
rect 148464 7812 148492 7868
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148756 7812 148784 7868
rect 148464 6300 148784 7812
rect 148464 6244 148492 6300
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148756 6244 148784 6300
rect 130054 5460 130082 5516
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130346 5460 130374 5516
rect 130054 3948 130374 5460
rect 134204 5572 134260 5582
rect 134204 5124 134260 5516
rect 134204 5058 134260 5068
rect 130054 3892 130082 3948
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130346 3892 130374 3948
rect 130054 3076 130374 3892
rect 148464 4732 148784 6244
rect 148464 4676 148492 4732
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148756 4676 148784 4732
rect 148464 3164 148784 4676
rect 148464 3108 148492 3164
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148756 3108 148784 3164
rect 148464 3076 148784 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__I dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 60592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__I1
timestamp 1666464484
transform -1 0 75264 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__S
timestamp 1666464484
transform -1 0 73920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__I
timestamp 1666464484
transform 1 0 38864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__I
timestamp 1666464484
transform 1 0 139776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I0
timestamp 1666464484
transform 1 0 125888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I1
timestamp 1666464484
transform 1 0 123088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__S
timestamp 1666464484
transform 1 0 125440 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__I1
timestamp 1666464484
transform -1 0 76832 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__S
timestamp 1666464484
transform -1 0 74368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I0
timestamp 1666464484
transform -1 0 126000 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I1
timestamp 1666464484
transform -1 0 121968 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__S
timestamp 1666464484
transform 1 0 124096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__I
timestamp 1666464484
transform 1 0 60144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1666464484
transform 1 0 131936 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__I0
timestamp 1666464484
transform -1 0 140000 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__S
timestamp 1666464484
transform 1 0 142128 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I0
timestamp 1666464484
transform 1 0 135744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I1
timestamp 1666464484
transform -1 0 139552 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__S
timestamp 1666464484
transform -1 0 139104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I0
timestamp 1666464484
transform -1 0 138096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__S
timestamp 1666464484
transform 1 0 139104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I0
timestamp 1666464484
transform 1 0 136192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I1
timestamp 1666464484
transform -1 0 139216 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__S
timestamp 1666464484
transform 1 0 138096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I0
timestamp 1666464484
transform -1 0 138992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__S
timestamp 1666464484
transform -1 0 139440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1666464484
transform 1 0 140784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__I0
timestamp 1666464484
transform -1 0 138768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__I1
timestamp 1666464484
transform 1 0 140784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__S
timestamp 1666464484
transform 1 0 141232 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I0
timestamp 1666464484
transform -1 0 135296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__S
timestamp 1666464484
transform -1 0 135744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__I0
timestamp 1666464484
transform 1 0 135184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__I1
timestamp 1666464484
transform 1 0 138768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__S
timestamp 1666464484
transform 1 0 138432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__I
timestamp 1666464484
transform 1 0 130032 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__I0
timestamp 1666464484
transform 1 0 132496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__I0
timestamp 1666464484
transform 1 0 134624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__I1
timestamp 1666464484
transform 1 0 134176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__S
timestamp 1666464484
transform 1 0 133728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__I0
timestamp 1666464484
transform 1 0 134960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I0
timestamp 1666464484
transform 1 0 132160 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I1
timestamp 1666464484
transform -1 0 131936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__S
timestamp 1666464484
transform 1 0 134736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__I0
timestamp 1666464484
transform -1 0 124320 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__I1
timestamp 1666464484
transform 1 0 125104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__I
timestamp 1666464484
transform -1 0 110880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__I1
timestamp 1666464484
transform -1 0 119616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__S
timestamp 1666464484
transform 1 0 118272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I0
timestamp 1666464484
transform -1 0 123648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I1
timestamp 1666464484
transform 1 0 125552 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__I0
timestamp 1666464484
transform 1 0 118160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__I1
timestamp 1666464484
transform 1 0 117712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__S
timestamp 1666464484
transform 1 0 115360 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I
timestamp 1666464484
transform 1 0 60592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__I
timestamp 1666464484
transform 1 0 87360 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__I0
timestamp 1666464484
transform -1 0 109200 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__I1
timestamp 1666464484
transform -1 0 110880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__S
timestamp 1666464484
transform 1 0 109424 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I1
timestamp 1666464484
transform 1 0 110880 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__S
timestamp 1666464484
transform 1 0 110656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__I0
timestamp 1666464484
transform 1 0 110768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__I1
timestamp 1666464484
transform -1 0 110208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__S
timestamp 1666464484
transform -1 0 108304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__I0
timestamp 1666464484
transform -1 0 109984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__I1
timestamp 1666464484
transform 1 0 111328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__S
timestamp 1666464484
transform 1 0 110880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__I0
timestamp 1666464484
transform 1 0 107520 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__I1
timestamp 1666464484
transform -1 0 108864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__S
timestamp 1666464484
transform 1 0 105728 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__I
timestamp 1666464484
transform -1 0 50624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__I
timestamp 1666464484
transform 1 0 92512 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__I0
timestamp 1666464484
transform -1 0 104048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__I1
timestamp 1666464484
transform 1 0 107072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__S
timestamp 1666464484
transform -1 0 105280 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__I0
timestamp 1666464484
transform -1 0 105168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__I1
timestamp 1666464484
transform -1 0 107296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__S
timestamp 1666464484
transform 1 0 106176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__I0
timestamp 1666464484
transform 1 0 103488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__I1
timestamp 1666464484
transform 1 0 107520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__S
timestamp 1666464484
transform 1 0 107072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__I
timestamp 1666464484
transform -1 0 89152 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__I0
timestamp 1666464484
transform 1 0 96096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__I1
timestamp 1666464484
transform -1 0 97328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__I0
timestamp 1666464484
transform -1 0 96768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__I1
timestamp 1666464484
transform 1 0 96096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__S
timestamp 1666464484
transform 1 0 93744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__I0
timestamp 1666464484
transform -1 0 93296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__I1
timestamp 1666464484
transform -1 0 96096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__I0
timestamp 1666464484
transform 1 0 96432 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__I1
timestamp 1666464484
transform 1 0 95984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__S
timestamp 1666464484
transform -1 0 94080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__I0
timestamp 1666464484
transform -1 0 89600 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__I1
timestamp 1666464484
transform -1 0 93072 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__I
timestamp 1666464484
transform 1 0 85456 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__I0
timestamp 1666464484
transform -1 0 89936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__I1
timestamp 1666464484
transform -1 0 89488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__S
timestamp 1666464484
transform -1 0 87136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__I0
timestamp 1666464484
transform 1 0 91168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__I1
timestamp 1666464484
transform 1 0 92736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__I0
timestamp 1666464484
transform 1 0 89600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__I1
timestamp 1666464484
transform 1 0 89152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__S
timestamp 1666464484
transform -1 0 86688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__I
timestamp 1666464484
transform 1 0 74368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__I0
timestamp 1666464484
transform -1 0 76160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__I1
timestamp 1666464484
transform -1 0 78288 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__S
timestamp 1666464484
transform 1 0 79184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__I0
timestamp 1666464484
transform -1 0 79184 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__I1
timestamp 1666464484
transform 1 0 78512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__S
timestamp 1666464484
transform 1 0 78064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__I0
timestamp 1666464484
transform -1 0 77280 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__I1
timestamp 1666464484
transform -1 0 80416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__S
timestamp 1666464484
transform -1 0 76720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__I0
timestamp 1666464484
transform 1 0 75600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__I1
timestamp 1666464484
transform 1 0 78400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__S
timestamp 1666464484
transform 1 0 77952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__I0
timestamp 1666464484
transform -1 0 65968 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__I1
timestamp 1666464484
transform 1 0 67872 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__S
timestamp 1666464484
transform -1 0 64624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__I
timestamp 1666464484
transform -1 0 66416 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__I1
timestamp 1666464484
transform 1 0 67200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__I0
timestamp 1666464484
transform -1 0 65520 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__I1
timestamp 1666464484
transform 1 0 67424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__S
timestamp 1666464484
transform -1 0 66752 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__I1
timestamp 1666464484
transform -1 0 62944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__I
timestamp 1666464484
transform -1 0 63168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__I0
timestamp 1666464484
transform -1 0 62608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__I1
timestamp 1666464484
transform -1 0 65184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__S
timestamp 1666464484
transform -1 0 63840 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__I0
timestamp 1666464484
transform 1 0 66528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__I1
timestamp 1666464484
transform 1 0 66976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__I0
timestamp 1666464484
transform -1 0 62160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__I1
timestamp 1666464484
transform -1 0 64288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__S
timestamp 1666464484
transform 1 0 61600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__I0
timestamp 1666464484
transform 1 0 62048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__I1
timestamp 1666464484
transform 1 0 61600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__I0
timestamp 1666464484
transform -1 0 51632 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__I1
timestamp 1666464484
transform -1 0 53984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__S
timestamp 1666464484
transform -1 0 52864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__I
timestamp 1666464484
transform 1 0 52640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__I0
timestamp 1666464484
transform -1 0 55776 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__I1
timestamp 1666464484
transform 1 0 53648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__S
timestamp 1666464484
transform 1 0 52640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__I0
timestamp 1666464484
transform 1 0 49392 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__I1
timestamp 1666464484
transform -1 0 54880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__S
timestamp 1666464484
transform -1 0 54544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__I0
timestamp 1666464484
transform 1 0 53424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__I1
timestamp 1666464484
transform 1 0 55104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__S
timestamp 1666464484
transform 1 0 53536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__I
timestamp 1666464484
transform -1 0 59920 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__I0
timestamp 1666464484
transform 1 0 41776 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__I1
timestamp 1666464484
transform -1 0 45360 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__S
timestamp 1666464484
transform 1 0 44688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__I1
timestamp 1666464484
transform -1 0 44912 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__S
timestamp 1666464484
transform -1 0 45248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__I0
timestamp 1666464484
transform -1 0 46928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__I1
timestamp 1666464484
transform -1 0 45360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__S
timestamp 1666464484
transform 1 0 48160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__I0
timestamp 1666464484
transform 1 0 47488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__I1
timestamp 1666464484
transform 1 0 47936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__S
timestamp 1666464484
transform -1 0 47264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__I0
timestamp 1666464484
transform 1 0 29344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__I1
timestamp 1666464484
transform -1 0 31808 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__S
timestamp 1666464484
transform -1 0 31136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__I
timestamp 1666464484
transform -1 0 29680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__I1
timestamp 1666464484
transform 1 0 30352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__S
timestamp 1666464484
transform 1 0 29904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__I0
timestamp 1666464484
transform -1 0 29120 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__I1
timestamp 1666464484
transform -1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__S
timestamp 1666464484
transform -1 0 30688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__I1
timestamp 1666464484
transform 1 0 28000 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__S
timestamp 1666464484
transform -1 0 28672 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__I1
timestamp 1666464484
transform 1 0 19488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__S
timestamp 1666464484
transform -1 0 17584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__I1
timestamp 1666464484
transform 1 0 20496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__S
timestamp 1666464484
transform 1 0 20272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__I0
timestamp 1666464484
transform -1 0 17584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__I1
timestamp 1666464484
transform -1 0 19936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__S
timestamp 1666464484
transform -1 0 20384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__I1
timestamp 1666464484
transform 1 0 21504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__S
timestamp 1666464484
transform 1 0 19264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__A1
timestamp 1666464484
transform -1 0 16800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__A2
timestamp 1666464484
transform 1 0 16240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__A3
timestamp 1666464484
transform -1 0 7056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__A4
timestamp 1666464484
transform -1 0 9856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__288__I
timestamp 1666464484
transform 1 0 73248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__A2
timestamp 1666464484
transform 1 0 76160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A1
timestamp 1666464484
transform 1 0 53312 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A2
timestamp 1666464484
transform 1 0 54208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__I
timestamp 1666464484
transform -1 0 56000 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__I
timestamp 1666464484
transform -1 0 56448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__I
timestamp 1666464484
transform 1 0 29120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__I
timestamp 1666464484
transform -1 0 16016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__I
timestamp 1666464484
transform -1 0 21280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__I
timestamp 1666464484
transform 1 0 29568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__I
timestamp 1666464484
transform 1 0 30128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__I
timestamp 1666464484
transform 1 0 55888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__I
timestamp 1666464484
transform -1 0 63616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__I
timestamp 1666464484
transform 1 0 47600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__I
timestamp 1666464484
transform 1 0 46704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__I
timestamp 1666464484
transform -1 0 63168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__I
timestamp 1666464484
transform 1 0 58240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__I
timestamp 1666464484
transform 1 0 70224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__I
timestamp 1666464484
transform 1 0 62160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__I
timestamp 1666464484
transform 1 0 68096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__I
timestamp 1666464484
transform -1 0 65072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__I
timestamp 1666464484
transform 1 0 68208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__I
timestamp 1666464484
transform 1 0 84448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__I
timestamp 1666464484
transform -1 0 81424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__I
timestamp 1666464484
transform 1 0 80416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__I
timestamp 1666464484
transform -1 0 90048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__314__I
timestamp 1666464484
transform 1 0 90832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__I
timestamp 1666464484
transform 1 0 88480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__I
timestamp 1666464484
transform -1 0 99008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__I
timestamp 1666464484
transform -1 0 96656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__318__I
timestamp 1666464484
transform -1 0 103264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__I
timestamp 1666464484
transform -1 0 102816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__I
timestamp 1666464484
transform 1 0 119280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__321__I
timestamp 1666464484
transform -1 0 109200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__I
timestamp 1666464484
transform 1 0 110208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__323__I
timestamp 1666464484
transform 1 0 114912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__I
timestamp 1666464484
transform 1 0 116928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__I
timestamp 1666464484
transform -1 0 129136 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__I
timestamp 1666464484
transform 1 0 129808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__I
timestamp 1666464484
transform 1 0 16128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__I
timestamp 1666464484
transform -1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__I
timestamp 1666464484
transform 1 0 12656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__CLK
timestamp 1666464484
transform 1 0 18368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__CLK
timestamp 1666464484
transform 1 0 21504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__CLK
timestamp 1666464484
transform 1 0 28672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__CLK
timestamp 1666464484
transform 1 0 31696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__CLK
timestamp 1666464484
transform 1 0 47600 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__CLK
timestamp 1666464484
transform 1 0 45360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__CLK
timestamp 1666464484
transform 1 0 61264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__CLK
timestamp 1666464484
transform 1 0 57792 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__CLK
timestamp 1666464484
transform -1 0 60816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__CLK
timestamp 1666464484
transform 1 0 69328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__CLK
timestamp 1666464484
transform 1 0 60256 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__CLK
timestamp 1666464484
transform 1 0 69664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__CLK
timestamp 1666464484
transform 1 0 80416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__CLK
timestamp 1666464484
transform -1 0 79072 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__CLK
timestamp 1666464484
transform 1 0 85904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__CLK
timestamp 1666464484
transform 1 0 86800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__CLK
timestamp 1666464484
transform 1 0 95760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__CLK
timestamp 1666464484
transform 1 0 93856 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__CLK
timestamp 1666464484
transform 1 0 102592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__CLK
timestamp 1666464484
transform 1 0 102480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__CLK
timestamp 1666464484
transform 1 0 103936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__CLK
timestamp 1666464484
transform 1 0 104384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__CLK
timestamp 1666464484
transform 1 0 112336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__CLK
timestamp 1666464484
transform 1 0 114352 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__CLK
timestamp 1666464484
transform 1 0 126224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__CLK
timestamp 1666464484
transform 1 0 129360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__CLK
timestamp 1666464484
transform 1 0 121520 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__CLK
timestamp 1666464484
transform 1 0 120176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__D
timestamp 1666464484
transform -1 0 123872 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__CLK
timestamp 1666464484
transform 1 0 122192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__D
timestamp 1666464484
transform -1 0 127344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__CLK
timestamp 1666464484
transform 1 0 121184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__D
timestamp 1666464484
transform -1 0 126896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__CLK
timestamp 1666464484
transform 1 0 120176 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__CLK
timestamp 1666464484
transform 1 0 121968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__CLK
timestamp 1666464484
transform -1 0 21616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__D
timestamp 1666464484
transform 1 0 16912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__CLK
timestamp 1666464484
transform -1 0 11760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__372__CLK
timestamp 1666464484
transform 1 0 13664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__I
timestamp 1666464484
transform -1 0 6272 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__I
timestamp 1666464484
transform 1 0 9632 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__I
timestamp 1666464484
transform 1 0 13440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__I
timestamp 1666464484
transform -1 0 17136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__379__I
timestamp 1666464484
transform 1 0 21728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__380__I
timestamp 1666464484
transform 1 0 24192 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__I
timestamp 1666464484
transform 1 0 27104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__I
timestamp 1666464484
transform 1 0 29792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__I
timestamp 1666464484
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__I
timestamp 1666464484
transform 1 0 70112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__385__I
timestamp 1666464484
transform 1 0 25648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__I
timestamp 1666464484
transform 1 0 35056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__I
timestamp 1666464484
transform 1 0 38416 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__I
timestamp 1666464484
transform 1 0 41888 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__I
timestamp 1666464484
transform 1 0 51632 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__I
timestamp 1666464484
transform 1 0 51184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__I
timestamp 1666464484
transform 1 0 56112 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__I
timestamp 1666464484
transform 1 0 86576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__393__I
timestamp 1666464484
transform -1 0 7616 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__I
timestamp 1666464484
transform 1 0 10976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__I
timestamp 1666464484
transform 1 0 14784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__I
timestamp 1666464484
transform 1 0 19264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__I
timestamp 1666464484
transform 1 0 22400 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__I
timestamp 1666464484
transform 1 0 25536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__I
timestamp 1666464484
transform -1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__I
timestamp 1666464484
transform -1 0 31472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__I
timestamp 1666464484
transform 1 0 34160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__I
timestamp 1666464484
transform 1 0 36064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__I
timestamp 1666464484
transform 1 0 37968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__I
timestamp 1666464484
transform 1 0 39872 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__I
timestamp 1666464484
transform 1 0 41440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__I
timestamp 1666464484
transform 1 0 42896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__I
timestamp 1666464484
transform 1 0 57792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__I
timestamp 1666464484
transform 1 0 47376 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__I
timestamp 1666464484
transform -1 0 45696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__I
timestamp 1666464484
transform 1 0 48720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__I
timestamp 1666464484
transform 1 0 51968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__I
timestamp 1666464484
transform 1 0 55104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__I
timestamp 1666464484
transform -1 0 84672 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__I
timestamp 1666464484
transform 1 0 102592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__415__I
timestamp 1666464484
transform 1 0 110880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__I
timestamp 1666464484
transform -1 0 115584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__I
timestamp 1666464484
transform 1 0 114352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__418__I
timestamp 1666464484
transform 1 0 122080 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__I
timestamp 1666464484
transform 1 0 127344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__I
timestamp 1666464484
transform 1 0 126896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__I
timestamp 1666464484
transform 1 0 119280 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__I
timestamp 1666464484
transform -1 0 86240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__I
timestamp 1666464484
transform 1 0 80640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__424__I
timestamp 1666464484
transform 1 0 93408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__I
timestamp 1666464484
transform -1 0 72576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__I
timestamp 1666464484
transform 1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__I
timestamp 1666464484
transform -1 0 59696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__I
timestamp 1666464484
transform 1 0 90272 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__I
timestamp 1666464484
transform 1 0 38528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__I
timestamp 1666464484
transform 1 0 38080 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__431__I
timestamp 1666464484
transform -1 0 47376 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__I
timestamp 1666464484
transform 1 0 49168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__I
timestamp 1666464484
transform 1 0 56560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__I
timestamp 1666464484
transform 1 0 80192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__I
timestamp 1666464484
transform -1 0 101696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__I
timestamp 1666464484
transform 1 0 104384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__I
timestamp 1666464484
transform 1 0 106624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__I
timestamp 1666464484
transform 1 0 112224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__I
timestamp 1666464484
transform 1 0 111552 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__I
timestamp 1666464484
transform 1 0 113008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__I
timestamp 1666464484
transform 1 0 116256 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__I
timestamp 1666464484
transform 1 0 118496 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__I
timestamp 1666464484
transform 1 0 120288 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__I
timestamp 1666464484
transform 1 0 122752 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__I
timestamp 1666464484
transform 1 0 122976 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__I
timestamp 1666464484
transform 1 0 107968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__I
timestamp 1666464484
transform 1 0 128240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__I
timestamp 1666464484
transform 1 0 117488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__449__I
timestamp 1666464484
transform 1 0 133728 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__I
timestamp 1666464484
transform 1 0 127792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__I
timestamp 1666464484
transform 1 0 128688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__I
timestamp 1666464484
transform 1 0 130480 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__453__I
timestamp 1666464484
transform 1 0 134064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__I
timestamp 1666464484
transform 1 0 140784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__I
timestamp 1666464484
transform 1 0 142912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__456__I
timestamp 1666464484
transform 1 0 145488 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__I
timestamp 1666464484
transform 1 0 9632 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__I
timestamp 1666464484
transform 1 0 13552 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__I
timestamp 1666464484
transform 1 0 16464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__I
timestamp 1666464484
transform 1 0 18368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__461__I
timestamp 1666464484
transform 1 0 23296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__I
timestamp 1666464484
transform -1 0 20832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__I
timestamp 1666464484
transform 1 0 83888 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__I
timestamp 1666464484
transform 1 0 58688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_io_wbs_clk_I
timestamp 1666464484
transform 1 0 68544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_io_wbs_clk_I
timestamp 1666464484
transform 1 0 67088 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_io_wbs_clk_I
timestamp 1666464484
transform 1 0 70672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_io_wbs_clk_I
timestamp 1666464484
transform 1 0 72576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_io_wbs_clk_I
timestamp 1666464484
transform 1 0 79072 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1666464484
transform -1 0 8064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1666464484
transform 1 0 36848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1666464484
transform -1 0 37856 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1666464484
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1666464484
transform -1 0 42112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1666464484
transform -1 0 43904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1666464484
transform 1 0 46256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1666464484
transform -1 0 43344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1666464484
transform -1 0 48944 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1666464484
transform -1 0 50960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1666464484
transform -1 0 53536 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1666464484
transform 1 0 12208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1666464484
transform -1 0 54656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1666464484
transform -1 0 56112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1666464484
transform -1 0 58464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1666464484
transform -1 0 59360 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1666464484
transform -1 0 61824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1666464484
transform 1 0 64512 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1666464484
transform 1 0 65520 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1666464484
transform -1 0 67200 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1666464484
transform -1 0 68768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1666464484
transform 1 0 71008 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1666464484
transform 1 0 15680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1666464484
transform -1 0 72128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1666464484
transform 1 0 74592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1666464484
transform -1 0 19040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1666464484
transform 1 0 22848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1666464484
transform 1 0 25984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1666464484
transform -1 0 27776 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1666464484
transform -1 0 30464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1666464484
transform 1 0 33488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1666464484
transform 1 0 36064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1666464484
transform -1 0 78848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1666464484
transform -1 0 107744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1666464484
transform -1 0 109312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1666464484
transform -1 0 111328 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1666464484
transform 1 0 115808 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1666464484
transform -1 0 115024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1666464484
transform -1 0 117152 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1666464484
transform 1 0 120400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1666464484
transform -1 0 121072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1666464484
transform -1 0 122752 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1666464484
transform -1 0 124880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1666464484
transform -1 0 82432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1666464484
transform -1 0 126672 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1666464484
transform 1 0 129360 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1666464484
transform -1 0 131152 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1666464484
transform -1 0 131600 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1666464484
transform 1 0 132944 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1666464484
transform 1 0 136864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1666464484
transform -1 0 137424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1666464484
transform 1 0 138320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1666464484
transform 1 0 140336 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1666464484
transform -1 0 141568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1666464484
transform -1 0 86240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1666464484
transform -1 0 143584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1666464484
transform 1 0 146608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1666464484
transform -1 0 91840 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1666464484
transform -1 0 95648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1666464484
transform -1 0 97328 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1666464484
transform -1 0 99680 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1666464484
transform -1 0 101248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1666464484
transform -1 0 103936 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1666464484
transform -1 0 105728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1666464484
transform -1 0 57568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1666464484
transform -1 0 58912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1666464484
transform -1 0 23072 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1666464484
transform -1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1666464484
transform -1 0 34048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1666464484
transform 1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1666464484
transform 1 0 42560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1666464484
transform 1 0 47152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1666464484
transform -1 0 49952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1666464484
transform -1 0 51296 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1666464484
transform -1 0 6608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1666464484
transform -1 0 14560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1666464484
transform -1 0 58800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1666464484
transform 1 0 70560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1666464484
transform -1 0 69440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1666464484
transform 1 0 74928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1666464484
transform 1 0 79296 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1666464484
transform -1 0 81872 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1666464484
transform 1 0 86688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input84_I
timestamp 1666464484
transform 1 0 90608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input85_I
timestamp 1666464484
transform -1 0 93632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input86_I
timestamp 1666464484
transform -1 0 97664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input87_I
timestamp 1666464484
transform 1 0 22512 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input88_I
timestamp 1666464484
transform -1 0 101696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input89_I
timestamp 1666464484
transform 1 0 106624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input90_I
timestamp 1666464484
transform 1 0 111440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input91_I
timestamp 1666464484
transform -1 0 113792 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input92_I
timestamp 1666464484
transform -1 0 117376 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input93_I
timestamp 1666464484
transform -1 0 121856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input94_I
timestamp 1666464484
transform 1 0 131040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input95_I
timestamp 1666464484
transform 1 0 130256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input96_I
timestamp 1666464484
transform 1 0 134400 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input97_I
timestamp 1666464484
transform 1 0 137984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input98_I
timestamp 1666464484
transform -1 0 25088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input99_I
timestamp 1666464484
transform -1 0 141344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input100_I
timestamp 1666464484
transform -1 0 145376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input101_I
timestamp 1666464484
transform -1 0 31808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input102_I
timestamp 1666464484
transform -1 0 36960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input103_I
timestamp 1666464484
transform -1 0 40880 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input104_I
timestamp 1666464484
transform -1 0 44800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input105_I
timestamp 1666464484
transform -1 0 48832 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input106_I
timestamp 1666464484
transform -1 0 52416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input107_I
timestamp 1666464484
transform -1 0 56896 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input108_I
timestamp 1666464484
transform -1 0 5936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input109_I
timestamp 1666464484
transform -1 0 15008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input110_I
timestamp 1666464484
transform -1 0 22176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input111_I
timestamp 1666464484
transform -1 0 25760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input112_I
timestamp 1666464484
transform -1 0 33040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input113_I
timestamp 1666464484
transform 1 0 10080 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input114_I
timestamp 1666464484
transform -1 0 10976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output125_I
timestamp 1666464484
transform -1 0 81424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output126_I
timestamp 1666464484
transform -1 0 84448 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output127_I
timestamp 1666464484
transform -1 0 88032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output128_I
timestamp 1666464484
transform 1 0 91168 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output129_I
timestamp 1666464484
transform 1 0 96320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output130_I
timestamp 1666464484
transform 1 0 98336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output131_I
timestamp 1666464484
transform 1 0 100576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output132_I
timestamp 1666464484
transform 1 0 104160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output138_I
timestamp 1666464484
transform -1 0 43456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output145_I
timestamp 1666464484
transform -1 0 55888 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output146_I
timestamp 1666464484
transform -1 0 57568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output147_I
timestamp 1666464484
transform -1 0 59360 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output148_I
timestamp 1666464484
transform -1 0 60368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output149_I
timestamp 1666464484
transform -1 0 63056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output150_I
timestamp 1666464484
transform -1 0 64736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output151_I
timestamp 1666464484
transform -1 0 66528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output152_I
timestamp 1666464484
transform 1 0 68992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output153_I
timestamp 1666464484
transform -1 0 67872 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output154_I
timestamp 1666464484
transform -1 0 71680 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output157_I
timestamp 1666464484
transform -1 0 72800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output176_I
timestamp 1666464484
transform 1 0 81312 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output178_I
timestamp 1666464484
transform -1 0 127120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output180_I
timestamp 1666464484
transform -1 0 130256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output187_I
timestamp 1666464484
transform 1 0 87920 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output191_I
timestamp 1666464484
transform 1 0 93856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output192_I
timestamp 1666464484
transform -1 0 95200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output193_I
timestamp 1666464484
transform -1 0 98112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output194_I
timestamp 1666464484
transform -1 0 101248 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output195_I
timestamp 1666464484
transform -1 0 103600 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output196_I
timestamp 1666464484
transform -1 0 105280 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output197_I
timestamp 1666464484
transform -1 0 6272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output201_I
timestamp 1666464484
transform -1 0 70336 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output202_I
timestamp 1666464484
transform -1 0 71792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output203_I
timestamp 1666464484
transform -1 0 75712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output204_I
timestamp 1666464484
transform -1 0 82992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output205_I
timestamp 1666464484
transform 1 0 86352 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output206_I
timestamp 1666464484
transform 1 0 90048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output207_I
timestamp 1666464484
transform -1 0 94752 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output208_I
timestamp 1666464484
transform -1 0 98784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output210_I
timestamp 1666464484
transform -1 0 102816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output212_I
timestamp 1666464484
transform 1 0 111328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output214_I
timestamp 1666464484
transform -1 0 115808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output215_I
timestamp 1666464484
transform -1 0 123424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output216_I
timestamp 1666464484
transform -1 0 121408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output217_I
timestamp 1666464484
transform -1 0 131712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output218_I
timestamp 1666464484
transform 1 0 132944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output219_I
timestamp 1666464484
transform -1 0 135968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output221_I
timestamp 1666464484
transform -1 0 140000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output222_I
timestamp 1666464484
transform -1 0 144032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output224_I
timestamp 1666464484
transform 1 0 37184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output226_I
timestamp 1666464484
transform 1 0 45024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output227_I
timestamp 1666464484
transform 1 0 48160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output228_I
timestamp 1666464484
transform 1 0 53088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output229_I
timestamp 1666464484
transform 1 0 58128 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output230_I
timestamp 1666464484
transform 1 0 6048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output236_I
timestamp 1666464484
transform -1 0 81872 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output237_I
timestamp 1666464484
transform -1 0 84000 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output239_I
timestamp 1666464484
transform -1 0 90944 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41
timestamp 1666464484
transform 1 0 5936 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49
timestamp 1666464484
transform 1 0 6832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57
timestamp 1666464484
transform 1 0 7728 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1666464484
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 9408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82
timestamp 1666464484
transform 1 0 10528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86
timestamp 1666464484
transform 1 0 10976 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94
timestamp 1666464484
transform 1 0 11872 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100
timestamp 1666464484
transform 1 0 12544 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1666464484
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107
timestamp 1666464484
transform 1 0 13328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111
timestamp 1666464484
transform 1 0 13776 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_126
timestamp 1666464484
transform 1 0 15456 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_128
timestamp 1666464484
transform 1 0 15680 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131
timestamp 1666464484
transform 1 0 16016 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1666464484
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1666464484
transform 1 0 17248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_150
timestamp 1666464484
transform 1 0 18144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_158
timestamp 1666464484
transform 1 0 19040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1666464484
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_177
timestamp 1666464484
transform 1 0 21168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_181
timestamp 1666464484
transform 1 0 21616 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_183
timestamp 1666464484
transform 1 0 21840 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_190
timestamp 1666464484
transform 1 0 22624 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_194
timestamp 1666464484
transform 1 0 23072 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_202 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 23968 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1666464484
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_227
timestamp 1666464484
transform 1 0 26768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_231
timestamp 1666464484
transform 1 0 27216 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_238
timestamp 1666464484
transform 1 0 28000 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1666464484
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1666464484
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_254
timestamp 1666464484
transform 1 0 29792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_270
timestamp 1666464484
transform 1 0 31584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_278
timestamp 1666464484
transform 1 0 32480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1666464484
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_289
timestamp 1666464484
transform 1 0 33712 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_291
timestamp 1666464484
transform 1 0 33936 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_298
timestamp 1666464484
transform 1 0 34720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1666464484
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1666464484
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_324
timestamp 1666464484
transform 1 0 37632 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_326
timestamp 1666464484
transform 1 0 37856 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_333
timestamp 1666464484
transform 1 0 38640 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1666464484
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1666464484
transform 1 0 40768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_359
timestamp 1666464484
transform 1 0 41552 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_361
timestamp 1666464484
transform 1 0 41776 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_368
timestamp 1666464484
transform 1 0 42560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1666464484
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1666464484
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_394
timestamp 1666464484
transform 1 0 45472 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_396
timestamp 1666464484
transform 1 0 45696 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_403
timestamp 1666464484
transform 1 0 46480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1666464484
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_422
timestamp 1666464484
transform 1 0 48608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_430
timestamp 1666464484
transform 1 0 49504 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_434
timestamp 1666464484
transform 1 0 49952 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_442
timestamp 1666464484
transform 1 0 50848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_446
timestamp 1666464484
transform 1 0 51296 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1666464484
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_457
timestamp 1666464484
transform 1 0 52528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_459
timestamp 1666464484
transform 1 0 52752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_466
timestamp 1666464484
transform 1 0 53536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_483
timestamp 1666464484
transform 1 0 55440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1666464484
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1666464484
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_507
timestamp 1666464484
transform 1 0 58128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_509
timestamp 1666464484
transform 1 0 58352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_516
timestamp 1666464484
transform 1 0 59136 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_524
timestamp 1666464484
transform 1 0 60032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_527
timestamp 1666464484
transform 1 0 60368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_542
timestamp 1666464484
transform 1 0 62048 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_550
timestamp 1666464484
transform 1 0 62944 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_558
timestamp 1666464484
transform 1 0 63840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_562
timestamp 1666464484
transform 1 0 64288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_577
timestamp 1666464484
transform 1 0 65968 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_585
timestamp 1666464484
transform 1 0 66864 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_593
timestamp 1666464484
transform 1 0 67760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1666464484
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_612
timestamp 1666464484
transform 1 0 69888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_616
timestamp 1666464484
transform 1 0 70336 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_620
timestamp 1666464484
transform 1 0 70784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_624
timestamp 1666464484
transform 1 0 71232 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_626
timestamp 1666464484
transform 1 0 71456 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_629
timestamp 1666464484
transform 1 0 71792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_632
timestamp 1666464484
transform 1 0 72128 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_647
timestamp 1666464484
transform 1 0 73808 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_655
timestamp 1666464484
transform 1 0 74704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_659
timestamp 1666464484
transform 1 0 75152 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_661
timestamp 1666464484
transform 1 0 75376 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1666464484
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1666464484
transform 1 0 76048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_682
timestamp 1666464484
transform 1 0 77728 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_690
timestamp 1666464484
transform 1 0 78624 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_694
timestamp 1666464484
transform 1 0 79072 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_698
timestamp 1666464484
transform 1 0 79520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_702
timestamp 1666464484
transform 1 0 79968 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_717
timestamp 1666464484
transform 1 0 81648 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_725
timestamp 1666464484
transform 1 0 82544 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_729
timestamp 1666464484
transform 1 0 82992 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_733
timestamp 1666464484
transform 1 0 83440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_737
timestamp 1666464484
transform 1 0 83888 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_752
timestamp 1666464484
transform 1 0 85568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_760
timestamp 1666464484
transform 1 0 86464 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_764
timestamp 1666464484
transform 1 0 86912 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_768
timestamp 1666464484
transform 1 0 87360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_772
timestamp 1666464484
transform 1 0 87808 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_787
timestamp 1666464484
transform 1 0 89488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_795
timestamp 1666464484
transform 1 0 90384 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_799
timestamp 1666464484
transform 1 0 90832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_803
timestamp 1666464484
transform 1 0 91280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_807
timestamp 1666464484
transform 1 0 91728 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_822
timestamp 1666464484
transform 1 0 93408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_830
timestamp 1666464484
transform 1 0 94304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_834
timestamp 1666464484
transform 1 0 94752 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_838
timestamp 1666464484
transform 1 0 95200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_842
timestamp 1666464484
transform 1 0 95648 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_858
timestamp 1666464484
transform 1 0 97440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_866
timestamp 1666464484
transform 1 0 98336 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_870
timestamp 1666464484
transform 1 0 98784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_874
timestamp 1666464484
transform 1 0 99232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_877
timestamp 1666464484
transform 1 0 99568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_879
timestamp 1666464484
transform 1 0 99792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_894
timestamp 1666464484
transform 1 0 101472 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_902
timestamp 1666464484
transform 1 0 102368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_906
timestamp 1666464484
transform 1 0 102816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_912
timestamp 1666464484
transform 1 0 103488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_930
timestamp 1666464484
transform 1 0 105504 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_938
timestamp 1666464484
transform 1 0 106400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_942
timestamp 1666464484
transform 1 0 106848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_944
timestamp 1666464484
transform 1 0 107072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_947
timestamp 1666464484
transform 1 0 107408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_966
timestamp 1666464484
transform 1 0 109536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_974
timestamp 1666464484
transform 1 0 110432 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_978
timestamp 1666464484
transform 1 0 110880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_982
timestamp 1666464484
transform 1 0 111328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_985
timestamp 1666464484
transform 1 0 111664 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_987
timestamp 1666464484
transform 1 0 111888 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1002
timestamp 1666464484
transform 1 0 113568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1010
timestamp 1666464484
transform 1 0 114464 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1014
timestamp 1666464484
transform 1 0 114912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1017
timestamp 1666464484
transform 1 0 115248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1019
timestamp 1666464484
transform 1 0 115472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1022
timestamp 1666464484
transform 1 0 115808 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1038
timestamp 1666464484
transform 1 0 117600 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1046
timestamp 1666464484
transform 1 0 118496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1052
timestamp 1666464484
transform 1 0 119168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1055
timestamp 1666464484
transform 1 0 119504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1059
timestamp 1666464484
transform 1 0 119952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1074
timestamp 1666464484
transform 1 0 121632 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1082
timestamp 1666464484
transform 1 0 122528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1084
timestamp 1666464484
transform 1 0 122752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1087
timestamp 1666464484
transform 1 0 123088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1090
timestamp 1666464484
transform 1 0 123424 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1094
timestamp 1666464484
transform 1 0 123872 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1110
timestamp 1666464484
transform 1 0 125664 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1118
timestamp 1666464484
transform 1 0 126560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1122
timestamp 1666464484
transform 1 0 127008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1127
timestamp 1666464484
transform 1 0 127568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1131
timestamp 1666464484
transform 1 0 128016 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1146
timestamp 1666464484
transform 1 0 129696 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1154
timestamp 1666464484
transform 1 0 130592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1157
timestamp 1666464484
transform 1 0 130928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1160
timestamp 1666464484
transform 1 0 131264 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1164
timestamp 1666464484
transform 1 0 131712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1182
timestamp 1666464484
transform 1 0 133728 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1192
timestamp 1666464484
transform 1 0 134848 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1202
timestamp 1666464484
transform 1 0 135968 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1218
timestamp 1666464484
transform 1 0 137760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1222
timestamp 1666464484
transform 1 0 138208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1224
timestamp 1666464484
transform 1 0 138432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1227
timestamp 1666464484
transform 1 0 138768 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1235
timestamp 1666464484
transform 1 0 139664 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1238
timestamp 1666464484
transform 1 0 140000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1254
timestamp 1666464484
transform 1 0 141792 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1258
timestamp 1666464484
transform 1 0 142240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1262
timestamp 1666464484
transform 1 0 142688 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1270
timestamp 1666464484
transform 1 0 143584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1274
timestamp 1666464484
transform 1 0 144032 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1290
timestamp 1666464484
transform 1 0 145824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1294
timestamp 1666464484
transform 1 0 146272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1297 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 146608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_2
timestamp 1666464484
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_18
timestamp 1666464484
transform 1 0 3360 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_26
timestamp 1666464484
transform 1 0 4256 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_42
timestamp 1666464484
transform 1 0 6048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_44
timestamp 1666464484
transform 1 0 6272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_47
timestamp 1666464484
transform 1 0 6608 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_51
timestamp 1666464484
transform 1 0 7056 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_59
timestamp 1666464484
transform 1 0 7952 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1666464484
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1666464484
transform 1 0 9520 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_108
timestamp 1666464484
transform 1 0 13440 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_112
timestamp 1666464484
transform 1 0 13888 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_118
timestamp 1666464484
transform 1 0 14560 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_122
timestamp 1666464484
transform 1 0 15008 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_130
timestamp 1666464484
transform 1 0 15904 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_132
timestamp 1666464484
transform 1 0 16128 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_135
timestamp 1666464484
transform 1 0 16464 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1666464484
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1666464484
transform 1 0 17472 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_179
timestamp 1666464484
transform 1 0 21392 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_187
timestamp 1666464484
transform 1 0 22288 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_191
timestamp 1666464484
transform 1 0 22736 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_207
timestamp 1666464484
transform 1 0 24528 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_209
timestamp 1666464484
transform 1 0 24752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1666464484
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1666464484
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_218
timestamp 1666464484
transform 1 0 25760 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_226
timestamp 1666464484
transform 1 0 26656 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_228
timestamp 1666464484
transform 1 0 26880 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_235
timestamp 1666464484
transform 1 0 27664 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_241
timestamp 1666464484
transform 1 0 28336 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_243
timestamp 1666464484
transform 1 0 28560 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_246
timestamp 1666464484
transform 1 0 28896 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_250
timestamp 1666464484
transform 1 0 29344 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_254
timestamp 1666464484
transform 1 0 29792 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_272
timestamp 1666464484
transform 1 0 31808 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_280
timestamp 1666464484
transform 1 0 32704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1666464484
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_286
timestamp 1666464484
transform 1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_292
timestamp 1666464484
transform 1 0 34048 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_308
timestamp 1666464484
transform 1 0 35840 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_318
timestamp 1666464484
transform 1 0 36960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_322
timestamp 1666464484
transform 1 0 37408 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_330
timestamp 1666464484
transform 1 0 38304 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_332
timestamp 1666464484
transform 1 0 38528 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_335
timestamp 1666464484
transform 1 0 38864 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_353
timestamp 1666464484
transform 1 0 40880 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_357
timestamp 1666464484
transform 1 0 41328 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_365
timestamp 1666464484
transform 1 0 42224 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_367
timestamp 1666464484
transform 1 0 42448 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_370
timestamp 1666464484
transform 1 0 42784 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_388
timestamp 1666464484
transform 1 0 44800 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_392
timestamp 1666464484
transform 1 0 45248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_400
timestamp 1666464484
transform 1 0 46144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_404
timestamp 1666464484
transform 1 0 46592 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_407
timestamp 1666464484
transform 1 0 46928 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_411
timestamp 1666464484
transform 1 0 47376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_415
timestamp 1666464484
transform 1 0 47824 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_417
timestamp 1666464484
transform 1 0 48048 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_420
timestamp 1666464484
transform 1 0 48384 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_424
timestamp 1666464484
transform 1 0 48832 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_428
timestamp 1666464484
transform 1 0 49280 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_444
timestamp 1666464484
transform 1 0 51072 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_462
timestamp 1666464484
transform 1 0 53088 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_464
timestamp 1666464484
transform 1 0 53312 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_467
timestamp 1666464484
transform 1 0 53648 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_484
timestamp 1666464484
transform 1 0 55552 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_488
timestamp 1666464484
transform 1 0 56000 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1666464484
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_499
timestamp 1666464484
transform 1 0 57232 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_507
timestamp 1666464484
transform 1 0 58128 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_515
timestamp 1666464484
transform 1 0 59024 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1666464484
transform 1 0 64848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1666464484
transform 1 0 65184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_605
timestamp 1666464484
transform 1 0 69104 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_613
timestamp 1666464484
transform 1 0 70000 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_617
timestamp 1666464484
transform 1 0 70448 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_621
timestamp 1666464484
transform 1 0 70896 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_629
timestamp 1666464484
transform 1 0 71792 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_633
timestamp 1666464484
transform 1 0 72240 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_635
timestamp 1666464484
transform 1 0 72464 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_638
timestamp 1666464484
transform 1 0 72800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1666464484
transform 1 0 73136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_692
timestamp 1666464484
transform 1 0 78848 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_696
timestamp 1666464484
transform 1 0 79296 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_704
timestamp 1666464484
transform 1 0 80192 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_708
timestamp 1666464484
transform 1 0 80640 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_712
timestamp 1666464484
transform 1 0 81088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_716
timestamp 1666464484
transform 1 0 81536 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_719
timestamp 1666464484
transform 1 0 81872 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_751
timestamp 1666464484
transform 1 0 85456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_757
timestamp 1666464484
transform 1 0 86128 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_761
timestamp 1666464484
transform 1 0 86576 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_777
timestamp 1666464484
transform 1 0 88368 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_780
timestamp 1666464484
transform 1 0 88704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_783
timestamp 1666464484
transform 1 0 89040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_790
timestamp 1666464484
transform 1 0 89824 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_794
timestamp 1666464484
transform 1 0 90272 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_810
timestamp 1666464484
transform 1 0 92064 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_818
timestamp 1666464484
transform 1 0 92960 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_824
timestamp 1666464484
transform 1 0 93632 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_840
timestamp 1666464484
transform 1 0 95424 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_848
timestamp 1666464484
transform 1 0 96320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_854
timestamp 1666464484
transform 1 0 96992 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_860
timestamp 1666464484
transform 1 0 97664 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_892
timestamp 1666464484
transform 1 0 101248 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_896
timestamp 1666464484
transform 1 0 101696 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_912
timestamp 1666464484
transform 1 0 103488 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_918
timestamp 1666464484
transform 1 0 104160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_922
timestamp 1666464484
transform 1 0 104608 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_925
timestamp 1666464484
transform 1 0 104944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_960
timestamp 1666464484
transform 1 0 108864 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_976
timestamp 1666464484
transform 1 0 110656 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_980
timestamp 1666464484
transform 1 0 111104 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_984
timestamp 1666464484
transform 1 0 111552 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_992
timestamp 1666464484
transform 1 0 112448 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_996
timestamp 1666464484
transform 1 0 112896 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1000
timestamp 1666464484
transform 1 0 113344 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1004
timestamp 1666464484
transform 1 0 113792 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1008
timestamp 1666464484
transform 1 0 114240 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1011
timestamp 1666464484
transform 1 0 114576 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1047
timestamp 1666464484
transform 1 0 118608 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1055
timestamp 1666464484
transform 1 0 119504 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1063
timestamp 1666464484
transform 1 0 120400 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1067
timestamp 1666464484
transform 1 0 120848 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1069
timestamp 1666464484
transform 1 0 121072 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1072
timestamp 1666464484
transform 1 0 121408 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1076
timestamp 1666464484
transform 1 0 121856 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1078
timestamp 1666464484
transform 1 0 122080 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1081
timestamp 1666464484
transform 1 0 122416 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1117
timestamp 1666464484
transform 1 0 126448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1121
timestamp 1666464484
transform 1 0 126896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1128
timestamp 1666464484
transform 1 0 127680 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1134
timestamp 1666464484
transform 1 0 128352 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1138
timestamp 1666464484
transform 1 0 128800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1173
timestamp 1666464484
transform 1 0 132720 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1177
timestamp 1666464484
transform 1 0 133168 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1179
timestamp 1666464484
transform 1 0 133392 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1186
timestamp 1666464484
transform 1 0 134176 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1190
timestamp 1666464484
transform 1 0 134624 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1206
timestamp 1666464484
transform 1 0 136416 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1209
timestamp 1666464484
transform 1 0 136752 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1217
timestamp 1666464484
transform 1 0 137648 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1225
timestamp 1666464484
transform 1 0 138544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1229
timestamp 1666464484
transform 1 0 138992 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1245
timestamp 1666464484
transform 1 0 140784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1247
timestamp 1666464484
transform 1 0 141008 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1250
timestamp 1666464484
transform 1 0 141344 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1258
timestamp 1666464484
transform 1 0 142240 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1274
timestamp 1666464484
transform 1 0 144032 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1280
timestamp 1666464484
transform 1 0 144704 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1286
timestamp 1666464484
transform 1 0 145376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1294
timestamp 1666464484
transform 1 0 146272 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1310
timestamp 1666464484
transform 1 0 148064 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1312
timestamp 1666464484
transform 1 0 148288 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1666464484
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1666464484
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_37
timestamp 1666464484
transform 1 0 5488 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_41
timestamp 1666464484
transform 1 0 5936 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_44
timestamp 1666464484
transform 1 0 6272 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_52
timestamp 1666464484
transform 1 0 7168 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_54
timestamp 1666464484
transform 1 0 7392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_91
timestamp 1666464484
transform 1 0 11536 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_99
timestamp 1666464484
transform 1 0 12432 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_103
timestamp 1666464484
transform 1 0 12880 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1666464484
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_108
timestamp 1666464484
transform 1 0 13440 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_124
timestamp 1666464484
transform 1 0 15232 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_134
timestamp 1666464484
transform 1 0 16352 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_138
timestamp 1666464484
transform 1 0 16800 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_174
timestamp 1666464484
transform 1 0 20832 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1666464484
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_179
timestamp 1666464484
transform 1 0 21392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_182
timestamp 1666464484
transform 1 0 21728 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_186
timestamp 1666464484
transform 1 0 22176 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_202
timestamp 1666464484
transform 1 0 23968 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_244
timestamp 1666464484
transform 1 0 28672 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_250
timestamp 1666464484
transform 1 0 29344 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_255
timestamp 1666464484
transform 1 0 29904 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_259
timestamp 1666464484
transform 1 0 30352 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_291
timestamp 1666464484
transform 1 0 33936 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_307
timestamp 1666464484
transform 1 0 35728 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_315
timestamp 1666464484
transform 1 0 36624 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_321
timestamp 1666464484
transform 1 0 37296 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_353
timestamp 1666464484
transform 1 0 40880 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_388
timestamp 1666464484
transform 1 0 44800 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1666464484
transform 1 0 45248 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_395
timestamp 1666464484
transform 1 0 45584 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_399
timestamp 1666464484
transform 1 0 46032 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_405
timestamp 1666464484
transform 1 0 46704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_411
timestamp 1666464484
transform 1 0 47376 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_415
timestamp 1666464484
transform 1 0 47824 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_447
timestamp 1666464484
transform 1 0 51408 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_451
timestamp 1666464484
transform 1 0 51856 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_453
timestamp 1666464484
transform 1 0 52080 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_456
timestamp 1666464484
transform 1 0 52416 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1666464484
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_463
timestamp 1666464484
transform 1 0 53200 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_469
timestamp 1666464484
transform 1 0 53872 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_471
timestamp 1666464484
transform 1 0 54096 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_478
timestamp 1666464484
transform 1 0 54880 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_514
timestamp 1666464484
transform 1 0 58912 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_522
timestamp 1666464484
transform 1 0 59808 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_524
timestamp 1666464484
transform 1 0 60032 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1666464484
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_534
timestamp 1666464484
transform 1 0 61152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_585
timestamp 1666464484
transform 1 0 66864 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_589
timestamp 1666464484
transform 1 0 67312 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_595
timestamp 1666464484
transform 1 0 67984 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_599
timestamp 1666464484
transform 1 0 68432 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1666464484
transform 1 0 69104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_608
timestamp 1666464484
transform 1 0 69440 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_612
timestamp 1666464484
transform 1 0 69888 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_620
timestamp 1666464484
transform 1 0 70784 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_622
timestamp 1666464484
transform 1 0 71008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1666464484
transform 1 0 76720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_676
timestamp 1666464484
transform 1 0 77056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_711
timestamp 1666464484
transform 1 0 80976 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_727
timestamp 1666464484
transform 1 0 82768 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_735
timestamp 1666464484
transform 1 0 83664 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_739
timestamp 1666464484
transform 1 0 84112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_741
timestamp 1666464484
transform 1 0 84336 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_744
timestamp 1666464484
transform 1 0 84672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_747
timestamp 1666464484
transform 1 0 85008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_754
timestamp 1666464484
transform 1 0 85792 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_756
timestamp 1666464484
transform 1 0 86016 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_791
timestamp 1666464484
transform 1 0 89936 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_797
timestamp 1666464484
transform 1 0 90608 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_801
timestamp 1666464484
transform 1 0 91056 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_809
timestamp 1666464484
transform 1 0 91952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_813
timestamp 1666464484
transform 1 0 92400 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_815
timestamp 1666464484
transform 1 0 92624 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_818
timestamp 1666464484
transform 1 0 92960 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_828
timestamp 1666464484
transform 1 0 94080 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_864
timestamp 1666464484
transform 1 0 98112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_880
timestamp 1666464484
transform 1 0 99904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_884
timestamp 1666464484
transform 1 0 100352 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_886
timestamp 1666464484
transform 1 0 100576 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_889
timestamp 1666464484
transform 1 0 100912 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_897
timestamp 1666464484
transform 1 0 101808 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_901
timestamp 1666464484
transform 1 0 102256 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_903
timestamp 1666464484
transform 1 0 102480 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_906
timestamp 1666464484
transform 1 0 102816 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_942
timestamp 1666464484
transform 1 0 106848 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_950
timestamp 1666464484
transform 1 0 107744 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_956
timestamp 1666464484
transform 1 0 108416 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_960
timestamp 1666464484
transform 1 0 108864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_976
timestamp 1666464484
transform 1 0 110656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_980
timestamp 1666464484
transform 1 0 111104 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_984
timestamp 1666464484
transform 1 0 111552 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1000
timestamp 1666464484
transform 1 0 113344 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1008
timestamp 1666464484
transform 1 0 114240 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1012
timestamp 1666464484
transform 1 0 114688 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1016
timestamp 1666464484
transform 1 0 115136 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1022
timestamp 1666464484
transform 1 0 115808 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1028
timestamp 1666464484
transform 1 0 116480 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1031
timestamp 1666464484
transform 1 0 116816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1034
timestamp 1666464484
transform 1 0 117152 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1036
timestamp 1666464484
transform 1 0 117376 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1052
timestamp 1666464484
transform 1 0 119168 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1056
timestamp 1666464484
transform 1 0 119616 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1060
timestamp 1666464484
transform 1 0 120064 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1063
timestamp 1666464484
transform 1 0 120400 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1099
timestamp 1666464484
transform 1 0 124432 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1102
timestamp 1666464484
transform 1 0 124768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1137
timestamp 1666464484
transform 1 0 128688 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1145
timestamp 1666464484
transform 1 0 129584 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1153
timestamp 1666464484
transform 1 0 130480 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1159
timestamp 1666464484
transform 1 0 131152 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1163
timestamp 1666464484
transform 1 0 131600 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1166
timestamp 1666464484
transform 1 0 131936 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1170
timestamp 1666464484
transform 1 0 132384 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1173
timestamp 1666464484
transform 1 0 132720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1189
timestamp 1666464484
transform 1 0 134512 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1193
timestamp 1666464484
transform 1 0 134960 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1197
timestamp 1666464484
transform 1 0 135408 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1205
timestamp 1666464484
transform 1 0 136304 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1222
timestamp 1666464484
transform 1 0 138208 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1226
timestamp 1666464484
transform 1 0 138656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1230
timestamp 1666464484
transform 1 0 139104 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1234
timestamp 1666464484
transform 1 0 139552 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1238
timestamp 1666464484
transform 1 0 140000 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1244
timestamp 1666464484
transform 1 0 140672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1247 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 141008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1311
timestamp 1666464484
transform 1 0 148176 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1666464484
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1666464484
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1666464484
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1666464484
transform 1 0 9520 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_76
timestamp 1666464484
transform 1 0 9856 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_80
timestamp 1666464484
transform 1 0 10304 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_88
timestamp 1666464484
transform 1 0 11200 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_90
timestamp 1666464484
transform 1 0 11424 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_93
timestamp 1666464484
transform 1 0 11760 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_125
timestamp 1666464484
transform 1 0 15344 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_127
timestamp 1666464484
transform 1 0 15568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_134
timestamp 1666464484
transform 1 0 16352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_138
timestamp 1666464484
transform 1 0 16800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1666464484
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_144
timestamp 1666464484
transform 1 0 17472 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_160
timestamp 1666464484
transform 1 0 19264 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_168
timestamp 1666464484
transform 1 0 20160 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_174
timestamp 1666464484
transform 1 0 20832 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_178
timestamp 1666464484
transform 1 0 21280 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_182
timestamp 1666464484
transform 1 0 21728 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_198
timestamp 1666464484
transform 1 0 23520 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_206
timestamp 1666464484
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_210
timestamp 1666464484
transform 1 0 24864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1666464484
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_215
timestamp 1666464484
transform 1 0 25424 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_231
timestamp 1666464484
transform 1 0 27216 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_269
timestamp 1666464484
transform 1 0 31472 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_273
timestamp 1666464484
transform 1 0 31920 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_281
timestamp 1666464484
transform 1 0 32816 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1666464484
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_286
timestamp 1666464484
transform 1 0 33376 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_318
timestamp 1666464484
transform 1 0 36960 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_334
timestamp 1666464484
transform 1 0 38752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_337
timestamp 1666464484
transform 1 0 39088 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_345
timestamp 1666464484
transform 1 0 39984 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_353
timestamp 1666464484
transform 1 0 40880 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_357
timestamp 1666464484
transform 1 0 41328 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_373
timestamp 1666464484
transform 1 0 43120 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_411
timestamp 1666464484
transform 1 0 47376 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_415
timestamp 1666464484
transform 1 0 47824 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_423
timestamp 1666464484
transform 1 0 48720 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1666464484
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_428
timestamp 1666464484
transform 1 0 49280 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_460
timestamp 1666464484
transform 1 0 52864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_464
timestamp 1666464484
transform 1 0 53312 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_468
timestamp 1666464484
transform 1 0 53760 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_476
timestamp 1666464484
transform 1 0 54656 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_482
timestamp 1666464484
transform 1 0 55328 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_486
timestamp 1666464484
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_492
timestamp 1666464484
transform 1 0 56448 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1666464484
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_499
timestamp 1666464484
transform 1 0 57232 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_502
timestamp 1666464484
transform 1 0 57568 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_506
timestamp 1666464484
transform 1 0 58016 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_510
timestamp 1666464484
transform 1 0 58464 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_514
timestamp 1666464484
transform 1 0 58912 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_520
timestamp 1666464484
transform 1 0 59584 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_556
timestamp 1666464484
transform 1 0 63616 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_564
timestamp 1666464484
transform 1 0 64512 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_570
timestamp 1666464484
transform 1 0 65184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_605
timestamp 1666464484
transform 1 0 69104 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_609
timestamp 1666464484
transform 1 0 69552 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_625
timestamp 1666464484
transform 1 0 71344 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_633
timestamp 1666464484
transform 1 0 72240 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_637
timestamp 1666464484
transform 1 0 72688 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_641
timestamp 1666464484
transform 1 0 73136 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_649
timestamp 1666464484
transform 1 0 74032 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_653
timestamp 1666464484
transform 1 0 74480 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_655
timestamp 1666464484
transform 1 0 74704 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_662
timestamp 1666464484
transform 1 0 75488 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_698
timestamp 1666464484
transform 1 0 79520 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_704
timestamp 1666464484
transform 1 0 80192 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_708
timestamp 1666464484
transform 1 0 80640 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_712
timestamp 1666464484
transform 1 0 81088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_715
timestamp 1666464484
transform 1 0 81424 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_747
timestamp 1666464484
transform 1 0 85008 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_765
timestamp 1666464484
transform 1 0 87024 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_767
timestamp 1666464484
transform 1 0 87248 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_774
timestamp 1666464484
transform 1 0 88032 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_778
timestamp 1666464484
transform 1 0 88480 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_780
timestamp 1666464484
transform 1 0 88704 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_783
timestamp 1666464484
transform 1 0 89040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_788
timestamp 1666464484
transform 1 0 89600 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_792
timestamp 1666464484
transform 1 0 90048 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_824
timestamp 1666464484
transform 1 0 93632 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_832
timestamp 1666464484
transform 1 0 94528 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_834
timestamp 1666464484
transform 1 0 94752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_841
timestamp 1666464484
transform 1 0 95536 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_845
timestamp 1666464484
transform 1 0 95984 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_851
timestamp 1666464484
transform 1 0 96656 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_854
timestamp 1666464484
transform 1 0 96992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_859
timestamp 1666464484
transform 1 0 97552 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_863
timestamp 1666464484
transform 1 0 98000 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_868
timestamp 1666464484
transform 1 0 98560 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_872
timestamp 1666464484
transform 1 0 99008 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_906
timestamp 1666464484
transform 1 0 102816 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_910
timestamp 1666464484
transform 1 0 103264 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_916
timestamp 1666464484
transform 1 0 103936 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_922
timestamp 1666464484
transform 1 0 104608 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_925
timestamp 1666464484
transform 1 0 104944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_960
timestamp 1666464484
transform 1 0 108864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_966
timestamp 1666464484
transform 1 0 109536 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_970
timestamp 1666464484
transform 1 0 109984 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_974
timestamp 1666464484
transform 1 0 110432 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_986
timestamp 1666464484
transform 1 0 111776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_990
timestamp 1666464484
transform 1 0 112224 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_993
timestamp 1666464484
transform 1 0 112560 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_996
timestamp 1666464484
transform 1 0 112896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1031
timestamp 1666464484
transform 1 0 116816 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1035
timestamp 1666464484
transform 1 0 117264 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1042
timestamp 1666464484
transform 1 0 118048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1046
timestamp 1666464484
transform 1 0 118496 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1062
timestamp 1666464484
transform 1 0 120288 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1064
timestamp 1666464484
transform 1 0 120512 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1067
timestamp 1666464484
transform 1 0 120848 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1071
timestamp 1666464484
transform 1 0 121296 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1075
timestamp 1666464484
transform 1 0 121744 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1079
timestamp 1666464484
transform 1 0 122192 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1115
timestamp 1666464484
transform 1 0 126224 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1121
timestamp 1666464484
transform 1 0 126896 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1127
timestamp 1666464484
transform 1 0 127568 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1133
timestamp 1666464484
transform 1 0 128240 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1135
timestamp 1666464484
transform 1 0 128464 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1138
timestamp 1666464484
transform 1 0 128800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1145
timestamp 1666464484
transform 1 0 129584 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1149
timestamp 1666464484
transform 1 0 130032 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1153
timestamp 1666464484
transform 1 0 130480 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1161
timestamp 1666464484
transform 1 0 131376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1180
timestamp 1666464484
transform 1 0 133504 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1184
timestamp 1666464484
transform 1 0 133952 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1188
timestamp 1666464484
transform 1 0 134400 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1192
timestamp 1666464484
transform 1 0 134848 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1202
timestamp 1666464484
transform 1 0 135968 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1206
timestamp 1666464484
transform 1 0 136416 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1209
timestamp 1666464484
transform 1 0 136752 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1228
timestamp 1666464484
transform 1 0 138880 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1232
timestamp 1666464484
transform 1 0 139328 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1241
timestamp 1666464484
transform 1 0 140336 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1251
timestamp 1666464484
transform 1 0 141456 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1267
timestamp 1666464484
transform 1 0 143248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1275
timestamp 1666464484
transform 1 0 144144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1277
timestamp 1666464484
transform 1 0 144368 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_1280
timestamp 1666464484
transform 1 0 144704 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1312
timestamp 1666464484
transform 1 0 148288 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1666464484
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1666464484
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1666464484
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1666464484
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1666464484
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_108
timestamp 1666464484
transform 1 0 13440 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_116
timestamp 1666464484
transform 1 0 14336 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_152
timestamp 1666464484
transform 1 0 18368 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_169
timestamp 1666464484
transform 1 0 20272 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_173
timestamp 1666464484
transform 1 0 20720 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_179
timestamp 1666464484
transform 1 0 21392 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_211
timestamp 1666464484
transform 1 0 24976 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_219
timestamp 1666464484
transform 1 0 25872 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_226
timestamp 1666464484
transform 1 0 26656 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_234
timestamp 1666464484
transform 1 0 27552 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_244
timestamp 1666464484
transform 1 0 28672 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_250
timestamp 1666464484
transform 1 0 29344 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_253
timestamp 1666464484
transform 1 0 29680 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_317
timestamp 1666464484
transform 1 0 36848 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_321
timestamp 1666464484
transform 1 0 37296 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_353
timestamp 1666464484
transform 1 0 40880 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_367
timestamp 1666464484
transform 1 0 42448 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_369
timestamp 1666464484
transform 1 0 42672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_385
timestamp 1666464484
transform 1 0 44464 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1666464484
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_392
timestamp 1666464484
transform 1 0 45248 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_408
timestamp 1666464484
transform 1 0 47040 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_414
timestamp 1666464484
transform 1 0 47712 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_418
timestamp 1666464484
transform 1 0 48160 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_434
timestamp 1666464484
transform 1 0 49952 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_440
timestamp 1666464484
transform 1 0 50624 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_448
timestamp 1666464484
transform 1 0 51520 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_456
timestamp 1666464484
transform 1 0 52416 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1666464484
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_463
timestamp 1666464484
transform 1 0 53200 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_472
timestamp 1666464484
transform 1 0 54208 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_488
timestamp 1666464484
transform 1 0 56000 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_496
timestamp 1666464484
transform 1 0 56896 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1666464484
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_534
timestamp 1666464484
transform 1 0 61152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_537
timestamp 1666464484
transform 1 0 61488 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_543
timestamp 1666464484
transform 1 0 62160 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_579
timestamp 1666464484
transform 1 0 66192 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_587
timestamp 1666464484
transform 1 0 67088 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_589
timestamp 1666464484
transform 1 0 67312 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_594
timestamp 1666464484
transform 1 0 67872 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_598
timestamp 1666464484
transform 1 0 68320 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1666464484
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_605
timestamp 1666464484
transform 1 0 69104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_656
timestamp 1666464484
transform 1 0 74816 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1666464484
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_676
timestamp 1666464484
transform 1 0 77056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_683
timestamp 1666464484
transform 1 0 77840 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_687
timestamp 1666464484
transform 1 0 78288 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_691
timestamp 1666464484
transform 1 0 78736 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_695
timestamp 1666464484
transform 1 0 79184 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_727
timestamp 1666464484
transform 1 0 82768 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_743
timestamp 1666464484
transform 1 0 84560 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_747
timestamp 1666464484
transform 1 0 85008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_755
timestamp 1666464484
transform 1 0 85904 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_763
timestamp 1666464484
transform 1 0 86800 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_799
timestamp 1666464484
transform 1 0 90832 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_815
timestamp 1666464484
transform 1 0 92624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_818
timestamp 1666464484
transform 1 0 92960 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_828
timestamp 1666464484
transform 1 0 94080 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_836
timestamp 1666464484
transform 1 0 94976 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_872
timestamp 1666464484
transform 1 0 99008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_880
timestamp 1666464484
transform 1 0 99904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_884
timestamp 1666464484
transform 1 0 100352 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_886
timestamp 1666464484
transform 1 0 100576 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_889
timestamp 1666464484
transform 1 0 100912 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_897
timestamp 1666464484
transform 1 0 101808 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_901
timestamp 1666464484
transform 1 0 102256 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_905
timestamp 1666464484
transform 1 0 102704 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_941
timestamp 1666464484
transform 1 0 106736 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_949
timestamp 1666464484
transform 1 0 107632 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_957
timestamp 1666464484
transform 1 0 108528 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_960
timestamp 1666464484
transform 1 0 108864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_963
timestamp 1666464484
transform 1 0 109200 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_971
timestamp 1666464484
transform 1 0 110096 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_975
timestamp 1666464484
transform 1 0 110544 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_978
timestamp 1666464484
transform 1 0 110880 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1010
timestamp 1666464484
transform 1 0 114464 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1017
timestamp 1666464484
transform 1 0 115248 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1025
timestamp 1666464484
transform 1 0 116144 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1031
timestamp 1666464484
transform 1 0 116816 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1033
timestamp 1666464484
transform 1 0 117040 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1036
timestamp 1666464484
transform 1 0 117376 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1052
timestamp 1666464484
transform 1 0 119168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1060
timestamp 1666464484
transform 1 0 120064 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1063
timestamp 1666464484
transform 1 0 120400 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1099
timestamp 1666464484
transform 1 0 124432 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1102
timestamp 1666464484
transform 1 0 124768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1137
timestamp 1666464484
transform 1 0 128688 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1141
timestamp 1666464484
transform 1 0 129136 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1145
timestamp 1666464484
transform 1 0 129584 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1161
timestamp 1666464484
transform 1 0 131376 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1169
timestamp 1666464484
transform 1 0 132272 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1173
timestamp 1666464484
transform 1 0 132720 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1189
timestamp 1666464484
transform 1 0 134512 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1197
timestamp 1666464484
transform 1 0 135408 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1204
timestamp 1666464484
transform 1 0 136192 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1221
timestamp 1666464484
transform 1 0 138096 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1238
timestamp 1666464484
transform 1 0 140000 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1244
timestamp 1666464484
transform 1 0 140672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1247
timestamp 1666464484
transform 1 0 141008 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_1251
timestamp 1666464484
transform 1 0 141456 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1283
timestamp 1666464484
transform 1 0 145040 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1299
timestamp 1666464484
transform 1 0 146832 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1307
timestamp 1666464484
transform 1 0 147728 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1311
timestamp 1666464484
transform 1 0 148176 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1666464484
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1666464484
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1666464484
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1666464484
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1666464484
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1666464484
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_144
timestamp 1666464484
transform 1 0 17472 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_154
timestamp 1666464484
transform 1 0 18592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_158
timestamp 1666464484
transform 1 0 19040 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_162
timestamp 1666464484
transform 1 0 19488 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_166
timestamp 1666464484
transform 1 0 19936 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_168
timestamp 1666464484
transform 1 0 20160 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_171
timestamp 1666464484
transform 1 0 20496 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_203
timestamp 1666464484
transform 1 0 24080 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_211
timestamp 1666464484
transform 1 0 24976 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_215
timestamp 1666464484
transform 1 0 25424 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_219
timestamp 1666464484
transform 1 0 25872 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_236
timestamp 1666464484
transform 1 0 27776 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_253
timestamp 1666464484
transform 1 0 29680 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_257
timestamp 1666464484
transform 1 0 30128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_261
timestamp 1666464484
transform 1 0 30576 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_277
timestamp 1666464484
transform 1 0 32368 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_281
timestamp 1666464484
transform 1 0 32816 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1666464484
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1666464484
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1666464484
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1666464484
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_357
timestamp 1666464484
transform 1 0 41328 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_373
timestamp 1666464484
transform 1 0 43120 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_381
timestamp 1666464484
transform 1 0 44016 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_388
timestamp 1666464484
transform 1 0 44800 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_392
timestamp 1666464484
transform 1 0 45248 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_410
timestamp 1666464484
transform 1 0 47264 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1666464484
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1666464484
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1666464484
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_499
timestamp 1666464484
transform 1 0 57232 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_509
timestamp 1666464484
transform 1 0 58352 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_513
timestamp 1666464484
transform 1 0 58800 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_521
timestamp 1666464484
transform 1 0 59696 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_525
timestamp 1666464484
transform 1 0 60144 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_528
timestamp 1666464484
transform 1 0 60480 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_545
timestamp 1666464484
transform 1 0 62384 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_547
timestamp 1666464484
transform 1 0 62608 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_550
timestamp 1666464484
transform 1 0 62944 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1666464484
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_570
timestamp 1666464484
transform 1 0 65184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_586
timestamp 1666464484
transform 1 0 66976 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_590
timestamp 1666464484
transform 1 0 67424 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_622
timestamp 1666464484
transform 1 0 71008 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1666464484
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_641
timestamp 1666464484
transform 1 0 73136 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_657
timestamp 1666464484
transform 1 0 74928 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_661
timestamp 1666464484
transform 1 0 75376 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_665
timestamp 1666464484
transform 1 0 75824 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_682
timestamp 1666464484
transform 1 0 77728 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_686
timestamp 1666464484
transform 1 0 78176 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_690
timestamp 1666464484
transform 1 0 78624 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_706
timestamp 1666464484
transform 1 0 80416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_712
timestamp 1666464484
transform 1 0 81088 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_744
timestamp 1666464484
transform 1 0 84672 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_748
timestamp 1666464484
transform 1 0 85120 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_750
timestamp 1666464484
transform 1 0 85344 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_753
timestamp 1666464484
transform 1 0 85680 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_763
timestamp 1666464484
transform 1 0 86800 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_780
timestamp 1666464484
transform 1 0 88704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_783
timestamp 1666464484
transform 1 0 89040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_786
timestamp 1666464484
transform 1 0 89376 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_790
timestamp 1666464484
transform 1 0 89824 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_806
timestamp 1666464484
transform 1 0 91616 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_816
timestamp 1666464484
transform 1 0 92736 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_826
timestamp 1666464484
transform 1 0 93856 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_843
timestamp 1666464484
transform 1 0 95760 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_847
timestamp 1666464484
transform 1 0 96208 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_851
timestamp 1666464484
transform 1 0 96656 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_854
timestamp 1666464484
transform 1 0 96992 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_886
timestamp 1666464484
transform 1 0 100576 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_902
timestamp 1666464484
transform 1 0 102368 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_910
timestamp 1666464484
transform 1 0 103264 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_914
timestamp 1666464484
transform 1 0 103712 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_922
timestamp 1666464484
transform 1 0 104608 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_925
timestamp 1666464484
transform 1 0 104944 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_942
timestamp 1666464484
transform 1 0 106848 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_946
timestamp 1666464484
transform 1 0 107296 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_950
timestamp 1666464484
transform 1 0 107744 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_982
timestamp 1666464484
transform 1 0 111328 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_990
timestamp 1666464484
transform 1 0 112224 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_996
timestamp 1666464484
transform 1 0 112896 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1012
timestamp 1666464484
transform 1 0 114688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1016
timestamp 1666464484
transform 1 0 115136 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1020
timestamp 1666464484
transform 1 0 115584 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1037
timestamp 1666464484
transform 1 0 117488 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1041
timestamp 1666464484
transform 1 0 117936 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_1045
timestamp 1666464484
transform 1 0 118384 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1061
timestamp 1666464484
transform 1 0 120176 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1067
timestamp 1666464484
transform 1 0 120848 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1069
timestamp 1666464484
transform 1 0 121072 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1072
timestamp 1666464484
transform 1 0 121408 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1080
timestamp 1666464484
transform 1 0 122304 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1082
timestamp 1666464484
transform 1 0 122528 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1117
timestamp 1666464484
transform 1 0 126448 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1123
timestamp 1666464484
transform 1 0 127120 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1129
timestamp 1666464484
transform 1 0 127792 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1133
timestamp 1666464484
transform 1 0 128240 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1135
timestamp 1666464484
transform 1 0 128464 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1138
timestamp 1666464484
transform 1 0 128800 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1202
timestamp 1666464484
transform 1 0 135968 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1206
timestamp 1666464484
transform 1 0 136416 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1209
timestamp 1666464484
transform 1 0 136752 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1217
timestamp 1666464484
transform 1 0 137648 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1223
timestamp 1666464484
transform 1 0 138320 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1227
timestamp 1666464484
transform 1 0 138768 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_1231
timestamp 1666464484
transform 1 0 139216 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1263
timestamp 1666464484
transform 1 0 142800 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1271
timestamp 1666464484
transform 1 0 143696 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1275
timestamp 1666464484
transform 1 0 144144 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1277
timestamp 1666464484
transform 1 0 144368 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_1280
timestamp 1666464484
transform 1 0 144704 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1312
timestamp 1666464484
transform 1 0 148288 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1666464484
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1666464484
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1666464484
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1666464484
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1666464484
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1666464484
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1666464484
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1666464484
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_179
timestamp 1666464484
transform 1 0 21392 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_211
timestamp 1666464484
transform 1 0 24976 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_227
timestamp 1666464484
transform 1 0 26768 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_235
timestamp 1666464484
transform 1 0 27664 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_237
timestamp 1666464484
transform 1 0 27888 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_240
timestamp 1666464484
transform 1 0 28224 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_244
timestamp 1666464484
transform 1 0 28672 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1666464484
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1666464484
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1666464484
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1666464484
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1666464484
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1666464484
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1666464484
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1666464484
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1666464484
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1666464484
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_527
timestamp 1666464484
transform 1 0 60368 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_534
timestamp 1666464484
transform 1 0 61152 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_540
timestamp 1666464484
transform 1 0 61824 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_544
timestamp 1666464484
transform 1 0 62272 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_550
timestamp 1666464484
transform 1 0 62944 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_554
timestamp 1666464484
transform 1 0 63392 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_570
timestamp 1666464484
transform 1 0 65184 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_580
timestamp 1666464484
transform 1 0 66304 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_584
timestamp 1666464484
transform 1 0 66752 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_588
timestamp 1666464484
transform 1 0 67200 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_596
timestamp 1666464484
transform 1 0 68096 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_600
timestamp 1666464484
transform 1 0 68544 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1666464484
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1666464484
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_669
timestamp 1666464484
transform 1 0 76272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1666464484
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_676
timestamp 1666464484
transform 1 0 77056 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_740
timestamp 1666464484
transform 1 0 84224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_744
timestamp 1666464484
transform 1 0 84672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_747
timestamp 1666464484
transform 1 0 85008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_755
timestamp 1666464484
transform 1 0 85904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_759
timestamp 1666464484
transform 1 0 86352 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_762
timestamp 1666464484
transform 1 0 86688 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_766
timestamp 1666464484
transform 1 0 87136 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_783
timestamp 1666464484
transform 1 0 89040 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_787
timestamp 1666464484
transform 1 0 89488 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_791
timestamp 1666464484
transform 1 0 89936 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_807
timestamp 1666464484
transform 1 0 91728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_815
timestamp 1666464484
transform 1 0 92624 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_818
timestamp 1666464484
transform 1 0 92960 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_822
timestamp 1666464484
transform 1 0 93408 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_824
timestamp 1666464484
transform 1 0 93632 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_827
timestamp 1666464484
transform 1 0 93968 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_844
timestamp 1666464484
transform 1 0 95872 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_848
timestamp 1666464484
transform 1 0 96320 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_852
timestamp 1666464484
transform 1 0 96768 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_884
timestamp 1666464484
transform 1 0 100352 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_886
timestamp 1666464484
transform 1 0 100576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_889
timestamp 1666464484
transform 1 0 100912 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_905
timestamp 1666464484
transform 1 0 102704 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_913
timestamp 1666464484
transform 1 0 103600 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_917
timestamp 1666464484
transform 1 0 104048 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_925
timestamp 1666464484
transform 1 0 104944 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_942
timestamp 1666464484
transform 1 0 106848 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_946
timestamp 1666464484
transform 1 0 107296 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_954
timestamp 1666464484
transform 1 0 108192 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_960
timestamp 1666464484
transform 1 0 108864 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1024
timestamp 1666464484
transform 1 0 116032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1028
timestamp 1666464484
transform 1 0 116480 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_1031
timestamp 1666464484
transform 1 0 116816 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1063
timestamp 1666464484
transform 1 0 120400 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1071
timestamp 1666464484
transform 1 0 121296 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1077
timestamp 1666464484
transform 1 0 121968 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1094
timestamp 1666464484
transform 1 0 123872 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1098
timestamp 1666464484
transform 1 0 124320 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1102
timestamp 1666464484
transform 1 0 124768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1109
timestamp 1666464484
transform 1 0 125552 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1113
timestamp 1666464484
transform 1 0 126000 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1117
timestamp 1666464484
transform 1 0 126448 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1121
timestamp 1666464484
transform 1 0 126896 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_1125
timestamp 1666464484
transform 1 0 127344 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1157
timestamp 1666464484
transform 1 0 130928 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1165
timestamp 1666464484
transform 1 0 131824 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1169
timestamp 1666464484
transform 1 0 132272 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1173
timestamp 1666464484
transform 1 0 132720 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1237
timestamp 1666464484
transform 1 0 139888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1241
timestamp 1666464484
transform 1 0 140336 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1244
timestamp 1666464484
transform 1 0 140672 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1308
timestamp 1666464484
transform 1 0 147840 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1312
timestamp 1666464484
transform 1 0 148288 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1666464484
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1666464484
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1666464484
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1666464484
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1666464484
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1666464484
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1666464484
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1666464484
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1666464484
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1666464484
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1666464484
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1666464484
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1666464484
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1666464484
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1666464484
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1666464484
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1666464484
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1666464484
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1666464484
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1666464484
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1666464484
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_499
timestamp 1666464484
transform 1 0 57232 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_531
timestamp 1666464484
transform 1 0 60816 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_539
timestamp 1666464484
transform 1 0 61712 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_545
timestamp 1666464484
transform 1 0 62384 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_549
timestamp 1666464484
transform 1 0 62832 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_552
timestamp 1666464484
transform 1 0 63168 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_556
timestamp 1666464484
transform 1 0 63616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_560
timestamp 1666464484
transform 1 0 64064 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_562
timestamp 1666464484
transform 1 0 64288 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1666464484
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_570
timestamp 1666464484
transform 1 0 65184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_577
timestamp 1666464484
transform 1 0 65968 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_581
timestamp 1666464484
transform 1 0 66416 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_613
timestamp 1666464484
transform 1 0 70000 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_629
timestamp 1666464484
transform 1 0 71792 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_637
timestamp 1666464484
transform 1 0 72688 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_641
timestamp 1666464484
transform 1 0 73136 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_705
timestamp 1666464484
transform 1 0 80304 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_709
timestamp 1666464484
transform 1 0 80752 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_712
timestamp 1666464484
transform 1 0 81088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_776
timestamp 1666464484
transform 1 0 88256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_780
timestamp 1666464484
transform 1 0 88704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_783
timestamp 1666464484
transform 1 0 89040 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_847
timestamp 1666464484
transform 1 0 96208 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_851
timestamp 1666464484
transform 1 0 96656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_854
timestamp 1666464484
transform 1 0 96992 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_918
timestamp 1666464484
transform 1 0 104160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_922
timestamp 1666464484
transform 1 0 104608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_925
timestamp 1666464484
transform 1 0 104944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_928
timestamp 1666464484
transform 1 0 105280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_992
timestamp 1666464484
transform 1 0 112448 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_996
timestamp 1666464484
transform 1 0 112896 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1060
timestamp 1666464484
transform 1 0 120064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1064
timestamp 1666464484
transform 1 0 120512 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_1067
timestamp 1666464484
transform 1 0 120848 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1083
timestamp 1666464484
transform 1 0 122640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1089
timestamp 1666464484
transform 1 0 123312 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1106
timestamp 1666464484
transform 1 0 125216 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1110
timestamp 1666464484
transform 1 0 125664 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_1114
timestamp 1666464484
transform 1 0 126112 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1130
timestamp 1666464484
transform 1 0 127904 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1134
timestamp 1666464484
transform 1 0 128352 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1138
timestamp 1666464484
transform 1 0 128800 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1202
timestamp 1666464484
transform 1 0 135968 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1206
timestamp 1666464484
transform 1 0 136416 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1209
timestamp 1666464484
transform 1 0 136752 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1273
timestamp 1666464484
transform 1 0 143920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1277
timestamp 1666464484
transform 1 0 144368 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_1280
timestamp 1666464484
transform 1 0 144704 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1312
timestamp 1666464484
transform 1 0 148288 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1666464484
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1666464484
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1666464484
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1666464484
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1666464484
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1666464484
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1666464484
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1666464484
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1666464484
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1666464484
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1666464484
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1666464484
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1666464484
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1666464484
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1666464484
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1666464484
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1666464484
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1666464484
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1666464484
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1666464484
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1666464484
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1666464484
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1666464484
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_534
timestamp 1666464484
transform 1 0 61152 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_566
timestamp 1666464484
transform 1 0 64736 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_569
timestamp 1666464484
transform 1 0 65072 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_601
timestamp 1666464484
transform 1 0 68656 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1666464484
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_669
timestamp 1666464484
transform 1 0 76272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1666464484
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_676
timestamp 1666464484
transform 1 0 77056 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_740
timestamp 1666464484
transform 1 0 84224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_744
timestamp 1666464484
transform 1 0 84672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_747
timestamp 1666464484
transform 1 0 85008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_811
timestamp 1666464484
transform 1 0 92176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_815
timestamp 1666464484
transform 1 0 92624 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_818
timestamp 1666464484
transform 1 0 92960 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_882
timestamp 1666464484
transform 1 0 100128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_886
timestamp 1666464484
transform 1 0 100576 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_889
timestamp 1666464484
transform 1 0 100912 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_953
timestamp 1666464484
transform 1 0 108080 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_957
timestamp 1666464484
transform 1 0 108528 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_960
timestamp 1666464484
transform 1 0 108864 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1024
timestamp 1666464484
transform 1 0 116032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1028
timestamp 1666464484
transform 1 0 116480 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1031
timestamp 1666464484
transform 1 0 116816 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1095
timestamp 1666464484
transform 1 0 123984 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1099
timestamp 1666464484
transform 1 0 124432 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1102
timestamp 1666464484
transform 1 0 124768 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1166
timestamp 1666464484
transform 1 0 131936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1170
timestamp 1666464484
transform 1 0 132384 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1173
timestamp 1666464484
transform 1 0 132720 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1237
timestamp 1666464484
transform 1 0 139888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1241
timestamp 1666464484
transform 1 0 140336 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1244
timestamp 1666464484
transform 1 0 140672 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1308
timestamp 1666464484
transform 1 0 147840 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1312
timestamp 1666464484
transform 1 0 148288 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1666464484
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1666464484
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1666464484
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1666464484
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1666464484
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1666464484
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1666464484
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1666464484
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1666464484
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1666464484
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1666464484
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1666464484
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1666464484
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1666464484
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1666464484
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1666464484
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1666464484
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1666464484
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1666464484
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1666464484
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1666464484
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1666464484
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_563
timestamp 1666464484
transform 1 0 64400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1666464484
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1666464484
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1666464484
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1666464484
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_641
timestamp 1666464484
transform 1 0 73136 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_705
timestamp 1666464484
transform 1 0 80304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_709
timestamp 1666464484
transform 1 0 80752 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_712
timestamp 1666464484
transform 1 0 81088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_776
timestamp 1666464484
transform 1 0 88256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_780
timestamp 1666464484
transform 1 0 88704 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_783
timestamp 1666464484
transform 1 0 89040 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_847
timestamp 1666464484
transform 1 0 96208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_851
timestamp 1666464484
transform 1 0 96656 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_854
timestamp 1666464484
transform 1 0 96992 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_918
timestamp 1666464484
transform 1 0 104160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_922
timestamp 1666464484
transform 1 0 104608 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_925
timestamp 1666464484
transform 1 0 104944 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_989
timestamp 1666464484
transform 1 0 112112 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_993
timestamp 1666464484
transform 1 0 112560 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_996
timestamp 1666464484
transform 1 0 112896 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1060
timestamp 1666464484
transform 1 0 120064 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1064
timestamp 1666464484
transform 1 0 120512 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1067
timestamp 1666464484
transform 1 0 120848 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1131
timestamp 1666464484
transform 1 0 128016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1135
timestamp 1666464484
transform 1 0 128464 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1138
timestamp 1666464484
transform 1 0 128800 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1202
timestamp 1666464484
transform 1 0 135968 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1206
timestamp 1666464484
transform 1 0 136416 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1209
timestamp 1666464484
transform 1 0 136752 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1273
timestamp 1666464484
transform 1 0 143920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1277
timestamp 1666464484
transform 1 0 144368 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_1280
timestamp 1666464484
transform 1 0 144704 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1312
timestamp 1666464484
transform 1 0 148288 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1666464484
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1666464484
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1666464484
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1666464484
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1666464484
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1666464484
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1666464484
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1666464484
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1666464484
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1666464484
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1666464484
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1666464484
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1666464484
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1666464484
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1666464484
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1666464484
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1666464484
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1666464484
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1666464484
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1666464484
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1666464484
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1666464484
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1666464484
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1666464484
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_598
timestamp 1666464484
transform 1 0 68320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1666464484
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_605
timestamp 1666464484
transform 1 0 69104 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_669
timestamp 1666464484
transform 1 0 76272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1666464484
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_676
timestamp 1666464484
transform 1 0 77056 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_740
timestamp 1666464484
transform 1 0 84224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_744
timestamp 1666464484
transform 1 0 84672 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_747
timestamp 1666464484
transform 1 0 85008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_811
timestamp 1666464484
transform 1 0 92176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_815
timestamp 1666464484
transform 1 0 92624 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_818
timestamp 1666464484
transform 1 0 92960 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_882
timestamp 1666464484
transform 1 0 100128 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_886
timestamp 1666464484
transform 1 0 100576 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_889
timestamp 1666464484
transform 1 0 100912 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_953
timestamp 1666464484
transform 1 0 108080 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_957
timestamp 1666464484
transform 1 0 108528 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_960
timestamp 1666464484
transform 1 0 108864 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1024
timestamp 1666464484
transform 1 0 116032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1028
timestamp 1666464484
transform 1 0 116480 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1031
timestamp 1666464484
transform 1 0 116816 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1095
timestamp 1666464484
transform 1 0 123984 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1099
timestamp 1666464484
transform 1 0 124432 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1102
timestamp 1666464484
transform 1 0 124768 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1166
timestamp 1666464484
transform 1 0 131936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1170
timestamp 1666464484
transform 1 0 132384 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1173
timestamp 1666464484
transform 1 0 132720 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1237
timestamp 1666464484
transform 1 0 139888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1241
timestamp 1666464484
transform 1 0 140336 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1244
timestamp 1666464484
transform 1 0 140672 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1308
timestamp 1666464484
transform 1 0 147840 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1312
timestamp 1666464484
transform 1 0 148288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1666464484
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1666464484
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1666464484
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1666464484
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1666464484
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1666464484
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1666464484
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1666464484
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1666464484
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1666464484
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1666464484
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1666464484
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1666464484
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1666464484
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1666464484
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1666464484
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1666464484
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1666464484
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1666464484
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1666464484
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1666464484
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1666464484
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_563
timestamp 1666464484
transform 1 0 64400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1666464484
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1666464484
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1666464484
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1666464484
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_641
timestamp 1666464484
transform 1 0 73136 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_705
timestamp 1666464484
transform 1 0 80304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_709
timestamp 1666464484
transform 1 0 80752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_712
timestamp 1666464484
transform 1 0 81088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_776
timestamp 1666464484
transform 1 0 88256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_780
timestamp 1666464484
transform 1 0 88704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_783
timestamp 1666464484
transform 1 0 89040 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_847
timestamp 1666464484
transform 1 0 96208 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_851
timestamp 1666464484
transform 1 0 96656 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_854
timestamp 1666464484
transform 1 0 96992 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_918
timestamp 1666464484
transform 1 0 104160 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_922
timestamp 1666464484
transform 1 0 104608 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_925
timestamp 1666464484
transform 1 0 104944 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_989
timestamp 1666464484
transform 1 0 112112 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_993
timestamp 1666464484
transform 1 0 112560 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_996
timestamp 1666464484
transform 1 0 112896 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1060
timestamp 1666464484
transform 1 0 120064 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1064
timestamp 1666464484
transform 1 0 120512 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1067
timestamp 1666464484
transform 1 0 120848 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1131
timestamp 1666464484
transform 1 0 128016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1135
timestamp 1666464484
transform 1 0 128464 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1138
timestamp 1666464484
transform 1 0 128800 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1202
timestamp 1666464484
transform 1 0 135968 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1206
timestamp 1666464484
transform 1 0 136416 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1209
timestamp 1666464484
transform 1 0 136752 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1273
timestamp 1666464484
transform 1 0 143920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1277
timestamp 1666464484
transform 1 0 144368 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_1280
timestamp 1666464484
transform 1 0 144704 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1312
timestamp 1666464484
transform 1 0 148288 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1666464484
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1666464484
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1666464484
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1666464484
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1666464484
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1666464484
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1666464484
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1666464484
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1666464484
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1666464484
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1666464484
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1666464484
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1666464484
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1666464484
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1666464484
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1666464484
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1666464484
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1666464484
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1666464484
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1666464484
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1666464484
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1666464484
transform 1 0 60368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1666464484
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1666464484
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_598
timestamp 1666464484
transform 1 0 68320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1666464484
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1666464484
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_669
timestamp 1666464484
transform 1 0 76272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1666464484
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_676
timestamp 1666464484
transform 1 0 77056 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_740
timestamp 1666464484
transform 1 0 84224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_744
timestamp 1666464484
transform 1 0 84672 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_747
timestamp 1666464484
transform 1 0 85008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_811
timestamp 1666464484
transform 1 0 92176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_815
timestamp 1666464484
transform 1 0 92624 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_818
timestamp 1666464484
transform 1 0 92960 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_882
timestamp 1666464484
transform 1 0 100128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_886
timestamp 1666464484
transform 1 0 100576 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_889
timestamp 1666464484
transform 1 0 100912 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_953
timestamp 1666464484
transform 1 0 108080 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_957
timestamp 1666464484
transform 1 0 108528 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_960
timestamp 1666464484
transform 1 0 108864 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1024
timestamp 1666464484
transform 1 0 116032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1028
timestamp 1666464484
transform 1 0 116480 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1031
timestamp 1666464484
transform 1 0 116816 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1095
timestamp 1666464484
transform 1 0 123984 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1099
timestamp 1666464484
transform 1 0 124432 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1102
timestamp 1666464484
transform 1 0 124768 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1166
timestamp 1666464484
transform 1 0 131936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1170
timestamp 1666464484
transform 1 0 132384 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1173
timestamp 1666464484
transform 1 0 132720 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1237
timestamp 1666464484
transform 1 0 139888 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1241
timestamp 1666464484
transform 1 0 140336 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1244
timestamp 1666464484
transform 1 0 140672 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1308
timestamp 1666464484
transform 1 0 147840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1312
timestamp 1666464484
transform 1 0 148288 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1666464484
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1666464484
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1666464484
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1666464484
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1666464484
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1666464484
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1666464484
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1666464484
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1666464484
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1666464484
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1666464484
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1666464484
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1666464484
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1666464484
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1666464484
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1666464484
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1666464484
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1666464484
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1666464484
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1666464484
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1666464484
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_499
timestamp 1666464484
transform 1 0 57232 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_563
timestamp 1666464484
transform 1 0 64400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1666464484
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1666464484
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1666464484
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1666464484
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_641
timestamp 1666464484
transform 1 0 73136 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_705
timestamp 1666464484
transform 1 0 80304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_709
timestamp 1666464484
transform 1 0 80752 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_712
timestamp 1666464484
transform 1 0 81088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_776
timestamp 1666464484
transform 1 0 88256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_780
timestamp 1666464484
transform 1 0 88704 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_783
timestamp 1666464484
transform 1 0 89040 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_847
timestamp 1666464484
transform 1 0 96208 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_851
timestamp 1666464484
transform 1 0 96656 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_854
timestamp 1666464484
transform 1 0 96992 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_918
timestamp 1666464484
transform 1 0 104160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_922
timestamp 1666464484
transform 1 0 104608 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_925
timestamp 1666464484
transform 1 0 104944 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_989
timestamp 1666464484
transform 1 0 112112 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_993
timestamp 1666464484
transform 1 0 112560 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_996
timestamp 1666464484
transform 1 0 112896 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1060
timestamp 1666464484
transform 1 0 120064 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1064
timestamp 1666464484
transform 1 0 120512 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1067
timestamp 1666464484
transform 1 0 120848 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1131
timestamp 1666464484
transform 1 0 128016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1135
timestamp 1666464484
transform 1 0 128464 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1138
timestamp 1666464484
transform 1 0 128800 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1202
timestamp 1666464484
transform 1 0 135968 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1206
timestamp 1666464484
transform 1 0 136416 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1209
timestamp 1666464484
transform 1 0 136752 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1273
timestamp 1666464484
transform 1 0 143920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1277
timestamp 1666464484
transform 1 0 144368 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_1280
timestamp 1666464484
transform 1 0 144704 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1312
timestamp 1666464484
transform 1 0 148288 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1666464484
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1666464484
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1666464484
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1666464484
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1666464484
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1666464484
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1666464484
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1666464484
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1666464484
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1666464484
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1666464484
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1666464484
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1666464484
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1666464484
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1666464484
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1666464484
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1666464484
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1666464484
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1666464484
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1666464484
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_463
timestamp 1666464484
transform 1 0 53200 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1666464484
transform 1 0 60368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1666464484
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1666464484
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1666464484
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1666464484
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1666464484
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_669
timestamp 1666464484
transform 1 0 76272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1666464484
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_676
timestamp 1666464484
transform 1 0 77056 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_740
timestamp 1666464484
transform 1 0 84224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_744
timestamp 1666464484
transform 1 0 84672 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_747
timestamp 1666464484
transform 1 0 85008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_811
timestamp 1666464484
transform 1 0 92176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_815
timestamp 1666464484
transform 1 0 92624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_818
timestamp 1666464484
transform 1 0 92960 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_882
timestamp 1666464484
transform 1 0 100128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_886
timestamp 1666464484
transform 1 0 100576 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_889
timestamp 1666464484
transform 1 0 100912 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_953
timestamp 1666464484
transform 1 0 108080 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_957
timestamp 1666464484
transform 1 0 108528 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_960
timestamp 1666464484
transform 1 0 108864 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1024
timestamp 1666464484
transform 1 0 116032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1028
timestamp 1666464484
transform 1 0 116480 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1031
timestamp 1666464484
transform 1 0 116816 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1095
timestamp 1666464484
transform 1 0 123984 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1099
timestamp 1666464484
transform 1 0 124432 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1102
timestamp 1666464484
transform 1 0 124768 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1166
timestamp 1666464484
transform 1 0 131936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1170
timestamp 1666464484
transform 1 0 132384 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1173
timestamp 1666464484
transform 1 0 132720 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1237
timestamp 1666464484
transform 1 0 139888 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1241
timestamp 1666464484
transform 1 0 140336 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1244
timestamp 1666464484
transform 1 0 140672 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1308
timestamp 1666464484
transform 1 0 147840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1312
timestamp 1666464484
transform 1 0 148288 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1666464484
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1666464484
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1666464484
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1666464484
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1666464484
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1666464484
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1666464484
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1666464484
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1666464484
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1666464484
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1666464484
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1666464484
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1666464484
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1666464484
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1666464484
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1666464484
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1666464484
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1666464484
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1666464484
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1666464484
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1666464484
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1666464484
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1666464484
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1666464484
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1666464484
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1666464484
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1666464484
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_641
timestamp 1666464484
transform 1 0 73136 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_705
timestamp 1666464484
transform 1 0 80304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_709
timestamp 1666464484
transform 1 0 80752 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_712
timestamp 1666464484
transform 1 0 81088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_776
timestamp 1666464484
transform 1 0 88256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_780
timestamp 1666464484
transform 1 0 88704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_783
timestamp 1666464484
transform 1 0 89040 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_847
timestamp 1666464484
transform 1 0 96208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_851
timestamp 1666464484
transform 1 0 96656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_854
timestamp 1666464484
transform 1 0 96992 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_918
timestamp 1666464484
transform 1 0 104160 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_922
timestamp 1666464484
transform 1 0 104608 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_925
timestamp 1666464484
transform 1 0 104944 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_989
timestamp 1666464484
transform 1 0 112112 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_993
timestamp 1666464484
transform 1 0 112560 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_996
timestamp 1666464484
transform 1 0 112896 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1060
timestamp 1666464484
transform 1 0 120064 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1064
timestamp 1666464484
transform 1 0 120512 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1067
timestamp 1666464484
transform 1 0 120848 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1131
timestamp 1666464484
transform 1 0 128016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1135
timestamp 1666464484
transform 1 0 128464 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1138
timestamp 1666464484
transform 1 0 128800 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1202
timestamp 1666464484
transform 1 0 135968 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1206
timestamp 1666464484
transform 1 0 136416 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1209
timestamp 1666464484
transform 1 0 136752 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1273
timestamp 1666464484
transform 1 0 143920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1277
timestamp 1666464484
transform 1 0 144368 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_1280
timestamp 1666464484
transform 1 0 144704 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1312
timestamp 1666464484
transform 1 0 148288 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1666464484
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1666464484
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1666464484
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1666464484
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1666464484
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1666464484
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1666464484
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1666464484
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1666464484
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1666464484
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1666464484
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1666464484
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1666464484
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1666464484
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1666464484
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1666464484
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1666464484
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1666464484
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1666464484
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1666464484
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1666464484
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1666464484
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1666464484
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1666464484
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_598
timestamp 1666464484
transform 1 0 68320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1666464484
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_605
timestamp 1666464484
transform 1 0 69104 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_669
timestamp 1666464484
transform 1 0 76272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_673
timestamp 1666464484
transform 1 0 76720 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_676
timestamp 1666464484
transform 1 0 77056 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_740
timestamp 1666464484
transform 1 0 84224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_744
timestamp 1666464484
transform 1 0 84672 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_747
timestamp 1666464484
transform 1 0 85008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_811
timestamp 1666464484
transform 1 0 92176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_815
timestamp 1666464484
transform 1 0 92624 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_818
timestamp 1666464484
transform 1 0 92960 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_882
timestamp 1666464484
transform 1 0 100128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_886
timestamp 1666464484
transform 1 0 100576 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_889
timestamp 1666464484
transform 1 0 100912 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_953
timestamp 1666464484
transform 1 0 108080 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_957
timestamp 1666464484
transform 1 0 108528 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_960
timestamp 1666464484
transform 1 0 108864 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1024
timestamp 1666464484
transform 1 0 116032 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1028
timestamp 1666464484
transform 1 0 116480 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1031
timestamp 1666464484
transform 1 0 116816 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1095
timestamp 1666464484
transform 1 0 123984 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1099
timestamp 1666464484
transform 1 0 124432 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1102
timestamp 1666464484
transform 1 0 124768 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1166
timestamp 1666464484
transform 1 0 131936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1170
timestamp 1666464484
transform 1 0 132384 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1173
timestamp 1666464484
transform 1 0 132720 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1237
timestamp 1666464484
transform 1 0 139888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1241
timestamp 1666464484
transform 1 0 140336 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1244
timestamp 1666464484
transform 1 0 140672 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1308
timestamp 1666464484
transform 1 0 147840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1312
timestamp 1666464484
transform 1 0 148288 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1666464484
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1666464484
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1666464484
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1666464484
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1666464484
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1666464484
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1666464484
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1666464484
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1666464484
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1666464484
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1666464484
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1666464484
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1666464484
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1666464484
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1666464484
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1666464484
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1666464484
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1666464484
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1666464484
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1666464484
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1666464484
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1666464484
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_563
timestamp 1666464484
transform 1 0 64400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1666464484
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1666464484
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_634
timestamp 1666464484
transform 1 0 72352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1666464484
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_641
timestamp 1666464484
transform 1 0 73136 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_705
timestamp 1666464484
transform 1 0 80304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_709
timestamp 1666464484
transform 1 0 80752 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_712
timestamp 1666464484
transform 1 0 81088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_776
timestamp 1666464484
transform 1 0 88256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_780
timestamp 1666464484
transform 1 0 88704 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_783
timestamp 1666464484
transform 1 0 89040 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_847
timestamp 1666464484
transform 1 0 96208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_851
timestamp 1666464484
transform 1 0 96656 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_854
timestamp 1666464484
transform 1 0 96992 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_918
timestamp 1666464484
transform 1 0 104160 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_922
timestamp 1666464484
transform 1 0 104608 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_925
timestamp 1666464484
transform 1 0 104944 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_989
timestamp 1666464484
transform 1 0 112112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_993
timestamp 1666464484
transform 1 0 112560 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_996
timestamp 1666464484
transform 1 0 112896 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1060
timestamp 1666464484
transform 1 0 120064 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1064
timestamp 1666464484
transform 1 0 120512 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1067
timestamp 1666464484
transform 1 0 120848 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1131
timestamp 1666464484
transform 1 0 128016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1135
timestamp 1666464484
transform 1 0 128464 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1138
timestamp 1666464484
transform 1 0 128800 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1202
timestamp 1666464484
transform 1 0 135968 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1206
timestamp 1666464484
transform 1 0 136416 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1209
timestamp 1666464484
transform 1 0 136752 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1273
timestamp 1666464484
transform 1 0 143920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1277
timestamp 1666464484
transform 1 0 144368 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_1280
timestamp 1666464484
transform 1 0 144704 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1312
timestamp 1666464484
transform 1 0 148288 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1666464484
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1666464484
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1666464484
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1666464484
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1666464484
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1666464484
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1666464484
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1666464484
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1666464484
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1666464484
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1666464484
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1666464484
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1666464484
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1666464484
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1666464484
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1666464484
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1666464484
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1666464484
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1666464484
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1666464484
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_463
timestamp 1666464484
transform 1 0 53200 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_527
timestamp 1666464484
transform 1 0 60368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1666464484
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1666464484
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_598
timestamp 1666464484
transform 1 0 68320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1666464484
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_605
timestamp 1666464484
transform 1 0 69104 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_669
timestamp 1666464484
transform 1 0 76272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_673
timestamp 1666464484
transform 1 0 76720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_676
timestamp 1666464484
transform 1 0 77056 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_740
timestamp 1666464484
transform 1 0 84224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_744
timestamp 1666464484
transform 1 0 84672 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_747
timestamp 1666464484
transform 1 0 85008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_811
timestamp 1666464484
transform 1 0 92176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_815
timestamp 1666464484
transform 1 0 92624 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_818
timestamp 1666464484
transform 1 0 92960 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_882
timestamp 1666464484
transform 1 0 100128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_886
timestamp 1666464484
transform 1 0 100576 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_889
timestamp 1666464484
transform 1 0 100912 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_953
timestamp 1666464484
transform 1 0 108080 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_957
timestamp 1666464484
transform 1 0 108528 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_960
timestamp 1666464484
transform 1 0 108864 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1024
timestamp 1666464484
transform 1 0 116032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1028
timestamp 1666464484
transform 1 0 116480 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1031
timestamp 1666464484
transform 1 0 116816 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1095
timestamp 1666464484
transform 1 0 123984 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1099
timestamp 1666464484
transform 1 0 124432 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1102
timestamp 1666464484
transform 1 0 124768 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1166
timestamp 1666464484
transform 1 0 131936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1170
timestamp 1666464484
transform 1 0 132384 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1173
timestamp 1666464484
transform 1 0 132720 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1237
timestamp 1666464484
transform 1 0 139888 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1241
timestamp 1666464484
transform 1 0 140336 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1244
timestamp 1666464484
transform 1 0 140672 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1308
timestamp 1666464484
transform 1 0 147840 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1312
timestamp 1666464484
transform 1 0 148288 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1666464484
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1666464484
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1666464484
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1666464484
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1666464484
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1666464484
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1666464484
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1666464484
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1666464484
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1666464484
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1666464484
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1666464484
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1666464484
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1666464484
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1666464484
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1666464484
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1666464484
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1666464484
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1666464484
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1666464484
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1666464484
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1666464484
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_563
timestamp 1666464484
transform 1 0 64400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1666464484
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1666464484
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1666464484
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1666464484
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_641
timestamp 1666464484
transform 1 0 73136 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_705
timestamp 1666464484
transform 1 0 80304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_709
timestamp 1666464484
transform 1 0 80752 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_712
timestamp 1666464484
transform 1 0 81088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_776
timestamp 1666464484
transform 1 0 88256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_780
timestamp 1666464484
transform 1 0 88704 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_783
timestamp 1666464484
transform 1 0 89040 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_847
timestamp 1666464484
transform 1 0 96208 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_851
timestamp 1666464484
transform 1 0 96656 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_854
timestamp 1666464484
transform 1 0 96992 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_918
timestamp 1666464484
transform 1 0 104160 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_922
timestamp 1666464484
transform 1 0 104608 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_925
timestamp 1666464484
transform 1 0 104944 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_989
timestamp 1666464484
transform 1 0 112112 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_993
timestamp 1666464484
transform 1 0 112560 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_996
timestamp 1666464484
transform 1 0 112896 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1060
timestamp 1666464484
transform 1 0 120064 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1064
timestamp 1666464484
transform 1 0 120512 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1067
timestamp 1666464484
transform 1 0 120848 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1131
timestamp 1666464484
transform 1 0 128016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1135
timestamp 1666464484
transform 1 0 128464 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1138
timestamp 1666464484
transform 1 0 128800 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1202
timestamp 1666464484
transform 1 0 135968 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1206
timestamp 1666464484
transform 1 0 136416 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1209
timestamp 1666464484
transform 1 0 136752 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1273
timestamp 1666464484
transform 1 0 143920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1277
timestamp 1666464484
transform 1 0 144368 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_1280
timestamp 1666464484
transform 1 0 144704 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1312
timestamp 1666464484
transform 1 0 148288 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1666464484
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1666464484
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1666464484
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1666464484
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1666464484
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1666464484
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1666464484
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1666464484
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1666464484
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1666464484
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1666464484
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1666464484
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1666464484
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1666464484
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1666464484
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1666464484
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1666464484
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1666464484
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1666464484
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1666464484
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1666464484
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_527
timestamp 1666464484
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1666464484
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1666464484
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_598
timestamp 1666464484
transform 1 0 68320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1666464484
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_605
timestamp 1666464484
transform 1 0 69104 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_669
timestamp 1666464484
transform 1 0 76272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_673
timestamp 1666464484
transform 1 0 76720 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_676
timestamp 1666464484
transform 1 0 77056 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_740
timestamp 1666464484
transform 1 0 84224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_744
timestamp 1666464484
transform 1 0 84672 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_747
timestamp 1666464484
transform 1 0 85008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_811
timestamp 1666464484
transform 1 0 92176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_815
timestamp 1666464484
transform 1 0 92624 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_818
timestamp 1666464484
transform 1 0 92960 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_882
timestamp 1666464484
transform 1 0 100128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_886
timestamp 1666464484
transform 1 0 100576 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_889
timestamp 1666464484
transform 1 0 100912 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_953
timestamp 1666464484
transform 1 0 108080 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_957
timestamp 1666464484
transform 1 0 108528 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_960
timestamp 1666464484
transform 1 0 108864 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1024
timestamp 1666464484
transform 1 0 116032 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1028
timestamp 1666464484
transform 1 0 116480 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1031
timestamp 1666464484
transform 1 0 116816 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1095
timestamp 1666464484
transform 1 0 123984 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1099
timestamp 1666464484
transform 1 0 124432 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1102
timestamp 1666464484
transform 1 0 124768 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1166
timestamp 1666464484
transform 1 0 131936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1170
timestamp 1666464484
transform 1 0 132384 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1173
timestamp 1666464484
transform 1 0 132720 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1237
timestamp 1666464484
transform 1 0 139888 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1241
timestamp 1666464484
transform 1 0 140336 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1244
timestamp 1666464484
transform 1 0 140672 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1308
timestamp 1666464484
transform 1 0 147840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1312
timestamp 1666464484
transform 1 0 148288 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1666464484
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1666464484
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1666464484
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1666464484
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1666464484
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1666464484
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1666464484
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1666464484
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1666464484
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1666464484
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1666464484
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1666464484
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1666464484
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1666464484
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1666464484
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1666464484
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1666464484
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1666464484
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1666464484
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1666464484
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1666464484
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1666464484
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_563
timestamp 1666464484
transform 1 0 64400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1666464484
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1666464484
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_634
timestamp 1666464484
transform 1 0 72352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1666464484
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_641
timestamp 1666464484
transform 1 0 73136 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_705
timestamp 1666464484
transform 1 0 80304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_709
timestamp 1666464484
transform 1 0 80752 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_712
timestamp 1666464484
transform 1 0 81088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_776
timestamp 1666464484
transform 1 0 88256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_780
timestamp 1666464484
transform 1 0 88704 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_783
timestamp 1666464484
transform 1 0 89040 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_847
timestamp 1666464484
transform 1 0 96208 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_851
timestamp 1666464484
transform 1 0 96656 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_854
timestamp 1666464484
transform 1 0 96992 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_918
timestamp 1666464484
transform 1 0 104160 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_922
timestamp 1666464484
transform 1 0 104608 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_925
timestamp 1666464484
transform 1 0 104944 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_989
timestamp 1666464484
transform 1 0 112112 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_993
timestamp 1666464484
transform 1 0 112560 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_996
timestamp 1666464484
transform 1 0 112896 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1060
timestamp 1666464484
transform 1 0 120064 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1064
timestamp 1666464484
transform 1 0 120512 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1067
timestamp 1666464484
transform 1 0 120848 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1131
timestamp 1666464484
transform 1 0 128016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1135
timestamp 1666464484
transform 1 0 128464 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1138
timestamp 1666464484
transform 1 0 128800 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1202
timestamp 1666464484
transform 1 0 135968 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1206
timestamp 1666464484
transform 1 0 136416 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1209
timestamp 1666464484
transform 1 0 136752 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1273
timestamp 1666464484
transform 1 0 143920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1277
timestamp 1666464484
transform 1 0 144368 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_1280
timestamp 1666464484
transform 1 0 144704 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1312
timestamp 1666464484
transform 1 0 148288 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1666464484
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1666464484
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1666464484
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1666464484
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1666464484
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1666464484
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1666464484
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1666464484
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1666464484
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1666464484
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1666464484
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1666464484
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1666464484
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1666464484
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1666464484
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1666464484
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1666464484
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1666464484
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1666464484
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1666464484
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1666464484
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_527
timestamp 1666464484
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1666464484
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1666464484
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_598
timestamp 1666464484
transform 1 0 68320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1666464484
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_605
timestamp 1666464484
transform 1 0 69104 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_669
timestamp 1666464484
transform 1 0 76272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_673
timestamp 1666464484
transform 1 0 76720 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_676
timestamp 1666464484
transform 1 0 77056 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_740
timestamp 1666464484
transform 1 0 84224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_744
timestamp 1666464484
transform 1 0 84672 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_747
timestamp 1666464484
transform 1 0 85008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_811
timestamp 1666464484
transform 1 0 92176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_815
timestamp 1666464484
transform 1 0 92624 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_818
timestamp 1666464484
transform 1 0 92960 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_882
timestamp 1666464484
transform 1 0 100128 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_886
timestamp 1666464484
transform 1 0 100576 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_889
timestamp 1666464484
transform 1 0 100912 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_953
timestamp 1666464484
transform 1 0 108080 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_957
timestamp 1666464484
transform 1 0 108528 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_960
timestamp 1666464484
transform 1 0 108864 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1024
timestamp 1666464484
transform 1 0 116032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1028
timestamp 1666464484
transform 1 0 116480 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1031
timestamp 1666464484
transform 1 0 116816 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1095
timestamp 1666464484
transform 1 0 123984 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1099
timestamp 1666464484
transform 1 0 124432 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1102
timestamp 1666464484
transform 1 0 124768 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1166
timestamp 1666464484
transform 1 0 131936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1170
timestamp 1666464484
transform 1 0 132384 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1173
timestamp 1666464484
transform 1 0 132720 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1237
timestamp 1666464484
transform 1 0 139888 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1241
timestamp 1666464484
transform 1 0 140336 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1244
timestamp 1666464484
transform 1 0 140672 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1308
timestamp 1666464484
transform 1 0 147840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1312
timestamp 1666464484
transform 1 0 148288 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1666464484
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1666464484
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1666464484
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1666464484
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1666464484
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1666464484
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1666464484
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1666464484
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1666464484
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1666464484
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1666464484
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1666464484
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1666464484
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1666464484
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1666464484
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1666464484
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1666464484
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1666464484
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1666464484
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1666464484
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1666464484
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1666464484
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_563
timestamp 1666464484
transform 1 0 64400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1666464484
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1666464484
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_634
timestamp 1666464484
transform 1 0 72352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1666464484
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_641
timestamp 1666464484
transform 1 0 73136 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_705
timestamp 1666464484
transform 1 0 80304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_709
timestamp 1666464484
transform 1 0 80752 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_712
timestamp 1666464484
transform 1 0 81088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_776
timestamp 1666464484
transform 1 0 88256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_780
timestamp 1666464484
transform 1 0 88704 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_783
timestamp 1666464484
transform 1 0 89040 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_847
timestamp 1666464484
transform 1 0 96208 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_851
timestamp 1666464484
transform 1 0 96656 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_854
timestamp 1666464484
transform 1 0 96992 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_918
timestamp 1666464484
transform 1 0 104160 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_922
timestamp 1666464484
transform 1 0 104608 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_925
timestamp 1666464484
transform 1 0 104944 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_989
timestamp 1666464484
transform 1 0 112112 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_993
timestamp 1666464484
transform 1 0 112560 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_996
timestamp 1666464484
transform 1 0 112896 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1060
timestamp 1666464484
transform 1 0 120064 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1064
timestamp 1666464484
transform 1 0 120512 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1067
timestamp 1666464484
transform 1 0 120848 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1131
timestamp 1666464484
transform 1 0 128016 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1135
timestamp 1666464484
transform 1 0 128464 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1138
timestamp 1666464484
transform 1 0 128800 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1202
timestamp 1666464484
transform 1 0 135968 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1206
timestamp 1666464484
transform 1 0 136416 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1209
timestamp 1666464484
transform 1 0 136752 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1273
timestamp 1666464484
transform 1 0 143920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1277
timestamp 1666464484
transform 1 0 144368 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_1280
timestamp 1666464484
transform 1 0 144704 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1312
timestamp 1666464484
transform 1 0 148288 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1666464484
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1666464484
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1666464484
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1666464484
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1666464484
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1666464484
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1666464484
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1666464484
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1666464484
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1666464484
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1666464484
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1666464484
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1666464484
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1666464484
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1666464484
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1666464484
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1666464484
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1666464484
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1666464484
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1666464484
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1666464484
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_527
timestamp 1666464484
transform 1 0 60368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1666464484
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1666464484
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_598
timestamp 1666464484
transform 1 0 68320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1666464484
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_605
timestamp 1666464484
transform 1 0 69104 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_669
timestamp 1666464484
transform 1 0 76272 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1666464484
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_676
timestamp 1666464484
transform 1 0 77056 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_740
timestamp 1666464484
transform 1 0 84224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_744
timestamp 1666464484
transform 1 0 84672 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_747
timestamp 1666464484
transform 1 0 85008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_811
timestamp 1666464484
transform 1 0 92176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_815
timestamp 1666464484
transform 1 0 92624 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_818
timestamp 1666464484
transform 1 0 92960 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_882
timestamp 1666464484
transform 1 0 100128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_886
timestamp 1666464484
transform 1 0 100576 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_889
timestamp 1666464484
transform 1 0 100912 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_953
timestamp 1666464484
transform 1 0 108080 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_957
timestamp 1666464484
transform 1 0 108528 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_960
timestamp 1666464484
transform 1 0 108864 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1024
timestamp 1666464484
transform 1 0 116032 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1028
timestamp 1666464484
transform 1 0 116480 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1031
timestamp 1666464484
transform 1 0 116816 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1095
timestamp 1666464484
transform 1 0 123984 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1099
timestamp 1666464484
transform 1 0 124432 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1102
timestamp 1666464484
transform 1 0 124768 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1166
timestamp 1666464484
transform 1 0 131936 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1170
timestamp 1666464484
transform 1 0 132384 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1173
timestamp 1666464484
transform 1 0 132720 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1237
timestamp 1666464484
transform 1 0 139888 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1241
timestamp 1666464484
transform 1 0 140336 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1244
timestamp 1666464484
transform 1 0 140672 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1308
timestamp 1666464484
transform 1 0 147840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1312
timestamp 1666464484
transform 1 0 148288 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1666464484
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1666464484
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1666464484
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1666464484
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1666464484
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1666464484
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1666464484
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1666464484
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1666464484
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1666464484
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1666464484
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1666464484
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1666464484
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1666464484
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1666464484
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1666464484
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1666464484
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1666464484
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1666464484
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1666464484
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1666464484
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1666464484
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_563
timestamp 1666464484
transform 1 0 64400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1666464484
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1666464484
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1666464484
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1666464484
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_641
timestamp 1666464484
transform 1 0 73136 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_705
timestamp 1666464484
transform 1 0 80304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_709
timestamp 1666464484
transform 1 0 80752 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_712
timestamp 1666464484
transform 1 0 81088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_776
timestamp 1666464484
transform 1 0 88256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_780
timestamp 1666464484
transform 1 0 88704 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_783
timestamp 1666464484
transform 1 0 89040 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_847
timestamp 1666464484
transform 1 0 96208 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_851
timestamp 1666464484
transform 1 0 96656 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_854
timestamp 1666464484
transform 1 0 96992 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_918
timestamp 1666464484
transform 1 0 104160 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_922
timestamp 1666464484
transform 1 0 104608 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_925
timestamp 1666464484
transform 1 0 104944 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_989
timestamp 1666464484
transform 1 0 112112 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_993
timestamp 1666464484
transform 1 0 112560 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_996
timestamp 1666464484
transform 1 0 112896 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1060
timestamp 1666464484
transform 1 0 120064 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1064
timestamp 1666464484
transform 1 0 120512 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1067
timestamp 1666464484
transform 1 0 120848 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1131
timestamp 1666464484
transform 1 0 128016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1135
timestamp 1666464484
transform 1 0 128464 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1138
timestamp 1666464484
transform 1 0 128800 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1202
timestamp 1666464484
transform 1 0 135968 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1206
timestamp 1666464484
transform 1 0 136416 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1209
timestamp 1666464484
transform 1 0 136752 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1273
timestamp 1666464484
transform 1 0 143920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1277
timestamp 1666464484
transform 1 0 144368 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_1280
timestamp 1666464484
transform 1 0 144704 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1312
timestamp 1666464484
transform 1 0 148288 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1666464484
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1666464484
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1666464484
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1666464484
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1666464484
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1666464484
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1666464484
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1666464484
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1666464484
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1666464484
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1666464484
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1666464484
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1666464484
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1666464484
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1666464484
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1666464484
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1666464484
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1666464484
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1666464484
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1666464484
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1666464484
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_527
timestamp 1666464484
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1666464484
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1666464484
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_598
timestamp 1666464484
transform 1 0 68320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1666464484
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605
timestamp 1666464484
transform 1 0 69104 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_669
timestamp 1666464484
transform 1 0 76272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1666464484
transform 1 0 76720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_676
timestamp 1666464484
transform 1 0 77056 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_740
timestamp 1666464484
transform 1 0 84224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_744
timestamp 1666464484
transform 1 0 84672 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_747
timestamp 1666464484
transform 1 0 85008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_811
timestamp 1666464484
transform 1 0 92176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_815
timestamp 1666464484
transform 1 0 92624 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_818
timestamp 1666464484
transform 1 0 92960 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_882
timestamp 1666464484
transform 1 0 100128 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_886
timestamp 1666464484
transform 1 0 100576 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_889
timestamp 1666464484
transform 1 0 100912 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_953
timestamp 1666464484
transform 1 0 108080 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_957
timestamp 1666464484
transform 1 0 108528 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_960
timestamp 1666464484
transform 1 0 108864 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1024
timestamp 1666464484
transform 1 0 116032 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1028
timestamp 1666464484
transform 1 0 116480 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1031
timestamp 1666464484
transform 1 0 116816 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1095
timestamp 1666464484
transform 1 0 123984 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1099
timestamp 1666464484
transform 1 0 124432 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1102
timestamp 1666464484
transform 1 0 124768 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1166
timestamp 1666464484
transform 1 0 131936 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1170
timestamp 1666464484
transform 1 0 132384 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1173
timestamp 1666464484
transform 1 0 132720 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1237
timestamp 1666464484
transform 1 0 139888 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1241
timestamp 1666464484
transform 1 0 140336 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1244
timestamp 1666464484
transform 1 0 140672 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1308
timestamp 1666464484
transform 1 0 147840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1312
timestamp 1666464484
transform 1 0 148288 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1666464484
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1666464484
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1666464484
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1666464484
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1666464484
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1666464484
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1666464484
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1666464484
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1666464484
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1666464484
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1666464484
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1666464484
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1666464484
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1666464484
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1666464484
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1666464484
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1666464484
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1666464484
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1666464484
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1666464484
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1666464484
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1666464484
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_563
timestamp 1666464484
transform 1 0 64400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1666464484
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1666464484
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1666464484
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1666464484
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_641
timestamp 1666464484
transform 1 0 73136 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_705
timestamp 1666464484
transform 1 0 80304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_709
timestamp 1666464484
transform 1 0 80752 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_712
timestamp 1666464484
transform 1 0 81088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_776
timestamp 1666464484
transform 1 0 88256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_780
timestamp 1666464484
transform 1 0 88704 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_783
timestamp 1666464484
transform 1 0 89040 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_847
timestamp 1666464484
transform 1 0 96208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_851
timestamp 1666464484
transform 1 0 96656 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_854
timestamp 1666464484
transform 1 0 96992 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_918
timestamp 1666464484
transform 1 0 104160 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_922
timestamp 1666464484
transform 1 0 104608 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_925
timestamp 1666464484
transform 1 0 104944 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_989
timestamp 1666464484
transform 1 0 112112 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_993
timestamp 1666464484
transform 1 0 112560 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_996
timestamp 1666464484
transform 1 0 112896 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1060
timestamp 1666464484
transform 1 0 120064 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1064
timestamp 1666464484
transform 1 0 120512 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1067
timestamp 1666464484
transform 1 0 120848 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1131
timestamp 1666464484
transform 1 0 128016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1135
timestamp 1666464484
transform 1 0 128464 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1138
timestamp 1666464484
transform 1 0 128800 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1202
timestamp 1666464484
transform 1 0 135968 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1206
timestamp 1666464484
transform 1 0 136416 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1209
timestamp 1666464484
transform 1 0 136752 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1273
timestamp 1666464484
transform 1 0 143920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1277
timestamp 1666464484
transform 1 0 144368 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_1280
timestamp 1666464484
transform 1 0 144704 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1312
timestamp 1666464484
transform 1 0 148288 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1666464484
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1666464484
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1666464484
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1666464484
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1666464484
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1666464484
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1666464484
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1666464484
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1666464484
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1666464484
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1666464484
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1666464484
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1666464484
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1666464484
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1666464484
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1666464484
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1666464484
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1666464484
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1666464484
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1666464484
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1666464484
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_527
timestamp 1666464484
transform 1 0 60368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1666464484
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1666464484
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1666464484
transform 1 0 68320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1666464484
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1666464484
transform 1 0 69104 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_669
timestamp 1666464484
transform 1 0 76272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1666464484
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_676
timestamp 1666464484
transform 1 0 77056 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_740
timestamp 1666464484
transform 1 0 84224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_744
timestamp 1666464484
transform 1 0 84672 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_747
timestamp 1666464484
transform 1 0 85008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_811
timestamp 1666464484
transform 1 0 92176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_815
timestamp 1666464484
transform 1 0 92624 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_818
timestamp 1666464484
transform 1 0 92960 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_882
timestamp 1666464484
transform 1 0 100128 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_886
timestamp 1666464484
transform 1 0 100576 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_889
timestamp 1666464484
transform 1 0 100912 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_953
timestamp 1666464484
transform 1 0 108080 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_957
timestamp 1666464484
transform 1 0 108528 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_960
timestamp 1666464484
transform 1 0 108864 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1024
timestamp 1666464484
transform 1 0 116032 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1028
timestamp 1666464484
transform 1 0 116480 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1031
timestamp 1666464484
transform 1 0 116816 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1095
timestamp 1666464484
transform 1 0 123984 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1099
timestamp 1666464484
transform 1 0 124432 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1102
timestamp 1666464484
transform 1 0 124768 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1166
timestamp 1666464484
transform 1 0 131936 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1170
timestamp 1666464484
transform 1 0 132384 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1173
timestamp 1666464484
transform 1 0 132720 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1237
timestamp 1666464484
transform 1 0 139888 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1241
timestamp 1666464484
transform 1 0 140336 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1244
timestamp 1666464484
transform 1 0 140672 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1308
timestamp 1666464484
transform 1 0 147840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1312
timestamp 1666464484
transform 1 0 148288 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1666464484
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1666464484
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1666464484
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1666464484
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1666464484
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1666464484
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1666464484
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1666464484
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1666464484
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1666464484
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1666464484
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1666464484
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1666464484
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1666464484
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1666464484
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1666464484
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1666464484
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1666464484
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1666464484
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1666464484
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1666464484
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1666464484
transform 1 0 57232 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_563
timestamp 1666464484
transform 1 0 64400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1666464484
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1666464484
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1666464484
transform 1 0 72352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1666464484
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_641
timestamp 1666464484
transform 1 0 73136 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_705
timestamp 1666464484
transform 1 0 80304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_709
timestamp 1666464484
transform 1 0 80752 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_712
timestamp 1666464484
transform 1 0 81088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_776
timestamp 1666464484
transform 1 0 88256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_780
timestamp 1666464484
transform 1 0 88704 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_783
timestamp 1666464484
transform 1 0 89040 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_847
timestamp 1666464484
transform 1 0 96208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_851
timestamp 1666464484
transform 1 0 96656 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_854
timestamp 1666464484
transform 1 0 96992 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_918
timestamp 1666464484
transform 1 0 104160 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_922
timestamp 1666464484
transform 1 0 104608 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_925
timestamp 1666464484
transform 1 0 104944 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_989
timestamp 1666464484
transform 1 0 112112 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_993
timestamp 1666464484
transform 1 0 112560 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_996
timestamp 1666464484
transform 1 0 112896 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1060
timestamp 1666464484
transform 1 0 120064 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1064
timestamp 1666464484
transform 1 0 120512 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1067
timestamp 1666464484
transform 1 0 120848 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1131
timestamp 1666464484
transform 1 0 128016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1135
timestamp 1666464484
transform 1 0 128464 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1138
timestamp 1666464484
transform 1 0 128800 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1202
timestamp 1666464484
transform 1 0 135968 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1206
timestamp 1666464484
transform 1 0 136416 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1209
timestamp 1666464484
transform 1 0 136752 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1273
timestamp 1666464484
transform 1 0 143920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1277
timestamp 1666464484
transform 1 0 144368 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_1280
timestamp 1666464484
transform 1 0 144704 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1312
timestamp 1666464484
transform 1 0 148288 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1666464484
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1666464484
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1666464484
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1666464484
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1666464484
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1666464484
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1666464484
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1666464484
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1666464484
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1666464484
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1666464484
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1666464484
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1666464484
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1666464484
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1666464484
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1666464484
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1666464484
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1666464484
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1666464484
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1666464484
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1666464484
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1666464484
transform 1 0 60368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1666464484
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1666464484
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1666464484
transform 1 0 68320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1666464484
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1666464484
transform 1 0 69104 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_669
timestamp 1666464484
transform 1 0 76272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1666464484
transform 1 0 76720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_676
timestamp 1666464484
transform 1 0 77056 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_740
timestamp 1666464484
transform 1 0 84224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_744
timestamp 1666464484
transform 1 0 84672 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_747
timestamp 1666464484
transform 1 0 85008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_811
timestamp 1666464484
transform 1 0 92176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_815
timestamp 1666464484
transform 1 0 92624 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_818
timestamp 1666464484
transform 1 0 92960 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_882
timestamp 1666464484
transform 1 0 100128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_886
timestamp 1666464484
transform 1 0 100576 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_889
timestamp 1666464484
transform 1 0 100912 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_953
timestamp 1666464484
transform 1 0 108080 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_957
timestamp 1666464484
transform 1 0 108528 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_960
timestamp 1666464484
transform 1 0 108864 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1024
timestamp 1666464484
transform 1 0 116032 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1028
timestamp 1666464484
transform 1 0 116480 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1031
timestamp 1666464484
transform 1 0 116816 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1095
timestamp 1666464484
transform 1 0 123984 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1099
timestamp 1666464484
transform 1 0 124432 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1102
timestamp 1666464484
transform 1 0 124768 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1166
timestamp 1666464484
transform 1 0 131936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1170
timestamp 1666464484
transform 1 0 132384 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1173
timestamp 1666464484
transform 1 0 132720 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1237
timestamp 1666464484
transform 1 0 139888 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1241
timestamp 1666464484
transform 1 0 140336 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1244
timestamp 1666464484
transform 1 0 140672 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1308
timestamp 1666464484
transform 1 0 147840 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1312
timestamp 1666464484
transform 1 0 148288 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1666464484
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1666464484
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1666464484
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1666464484
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1666464484
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1666464484
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1666464484
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1666464484
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1666464484
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1666464484
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1666464484
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1666464484
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1666464484
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1666464484
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1666464484
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1666464484
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1666464484
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1666464484
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1666464484
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1666464484
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1666464484
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1666464484
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1666464484
transform 1 0 64400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1666464484
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1666464484
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1666464484
transform 1 0 72352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1666464484
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_641
timestamp 1666464484
transform 1 0 73136 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_705
timestamp 1666464484
transform 1 0 80304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_709
timestamp 1666464484
transform 1 0 80752 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_712
timestamp 1666464484
transform 1 0 81088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_776
timestamp 1666464484
transform 1 0 88256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_780
timestamp 1666464484
transform 1 0 88704 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_783
timestamp 1666464484
transform 1 0 89040 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_847
timestamp 1666464484
transform 1 0 96208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_851
timestamp 1666464484
transform 1 0 96656 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_854
timestamp 1666464484
transform 1 0 96992 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_918
timestamp 1666464484
transform 1 0 104160 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_922
timestamp 1666464484
transform 1 0 104608 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_925
timestamp 1666464484
transform 1 0 104944 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_989
timestamp 1666464484
transform 1 0 112112 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_993
timestamp 1666464484
transform 1 0 112560 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_996
timestamp 1666464484
transform 1 0 112896 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1060
timestamp 1666464484
transform 1 0 120064 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1064
timestamp 1666464484
transform 1 0 120512 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1067
timestamp 1666464484
transform 1 0 120848 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1131
timestamp 1666464484
transform 1 0 128016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1135
timestamp 1666464484
transform 1 0 128464 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1138
timestamp 1666464484
transform 1 0 128800 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1202
timestamp 1666464484
transform 1 0 135968 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1206
timestamp 1666464484
transform 1 0 136416 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1209
timestamp 1666464484
transform 1 0 136752 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1273
timestamp 1666464484
transform 1 0 143920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1277
timestamp 1666464484
transform 1 0 144368 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_1280
timestamp 1666464484
transform 1 0 144704 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1312
timestamp 1666464484
transform 1 0 148288 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1666464484
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1666464484
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1666464484
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1666464484
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1666464484
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1666464484
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1666464484
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1666464484
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1666464484
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1666464484
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1666464484
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1666464484
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1666464484
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1666464484
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1666464484
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1666464484
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1666464484
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1666464484
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1666464484
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1666464484
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1666464484
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1666464484
transform 1 0 60368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1666464484
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1666464484
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1666464484
transform 1 0 68320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1666464484
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1666464484
transform 1 0 69104 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_669
timestamp 1666464484
transform 1 0 76272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1666464484
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_676
timestamp 1666464484
transform 1 0 77056 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_740
timestamp 1666464484
transform 1 0 84224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_744
timestamp 1666464484
transform 1 0 84672 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_747
timestamp 1666464484
transform 1 0 85008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_811
timestamp 1666464484
transform 1 0 92176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_815
timestamp 1666464484
transform 1 0 92624 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_818
timestamp 1666464484
transform 1 0 92960 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_882
timestamp 1666464484
transform 1 0 100128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_886
timestamp 1666464484
transform 1 0 100576 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_889
timestamp 1666464484
transform 1 0 100912 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_953
timestamp 1666464484
transform 1 0 108080 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_957
timestamp 1666464484
transform 1 0 108528 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_960
timestamp 1666464484
transform 1 0 108864 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1024
timestamp 1666464484
transform 1 0 116032 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1028
timestamp 1666464484
transform 1 0 116480 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1031
timestamp 1666464484
transform 1 0 116816 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1095
timestamp 1666464484
transform 1 0 123984 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1099
timestamp 1666464484
transform 1 0 124432 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1102
timestamp 1666464484
transform 1 0 124768 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1166
timestamp 1666464484
transform 1 0 131936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1170
timestamp 1666464484
transform 1 0 132384 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1173
timestamp 1666464484
transform 1 0 132720 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1237
timestamp 1666464484
transform 1 0 139888 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1241
timestamp 1666464484
transform 1 0 140336 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1244
timestamp 1666464484
transform 1 0 140672 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1308
timestamp 1666464484
transform 1 0 147840 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1312
timestamp 1666464484
transform 1 0 148288 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1666464484
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1666464484
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1666464484
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1666464484
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1666464484
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1666464484
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1666464484
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1666464484
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1666464484
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1666464484
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1666464484
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1666464484
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1666464484
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1666464484
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1666464484
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1666464484
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1666464484
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1666464484
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1666464484
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1666464484
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1666464484
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1666464484
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1666464484
transform 1 0 64400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1666464484
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1666464484
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1666464484
transform 1 0 72352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1666464484
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_641
timestamp 1666464484
transform 1 0 73136 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_705
timestamp 1666464484
transform 1 0 80304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_709
timestamp 1666464484
transform 1 0 80752 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_712
timestamp 1666464484
transform 1 0 81088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_776
timestamp 1666464484
transform 1 0 88256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_780
timestamp 1666464484
transform 1 0 88704 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_783
timestamp 1666464484
transform 1 0 89040 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_847
timestamp 1666464484
transform 1 0 96208 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_851
timestamp 1666464484
transform 1 0 96656 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_854
timestamp 1666464484
transform 1 0 96992 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_918
timestamp 1666464484
transform 1 0 104160 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_922
timestamp 1666464484
transform 1 0 104608 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_925
timestamp 1666464484
transform 1 0 104944 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_989
timestamp 1666464484
transform 1 0 112112 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_993
timestamp 1666464484
transform 1 0 112560 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_996
timestamp 1666464484
transform 1 0 112896 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1060
timestamp 1666464484
transform 1 0 120064 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1064
timestamp 1666464484
transform 1 0 120512 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1067
timestamp 1666464484
transform 1 0 120848 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1131
timestamp 1666464484
transform 1 0 128016 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1135
timestamp 1666464484
transform 1 0 128464 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1138
timestamp 1666464484
transform 1 0 128800 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1202
timestamp 1666464484
transform 1 0 135968 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1206
timestamp 1666464484
transform 1 0 136416 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1209
timestamp 1666464484
transform 1 0 136752 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1273
timestamp 1666464484
transform 1 0 143920 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1277
timestamp 1666464484
transform 1 0 144368 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_1280
timestamp 1666464484
transform 1 0 144704 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1312
timestamp 1666464484
transform 1 0 148288 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1666464484
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1666464484
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1666464484
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1666464484
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1666464484
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1666464484
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1666464484
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1666464484
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1666464484
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1666464484
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1666464484
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1666464484
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1666464484
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1666464484
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1666464484
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1666464484
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1666464484
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1666464484
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1666464484
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1666464484
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1666464484
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1666464484
transform 1 0 60368 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1666464484
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1666464484
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1666464484
transform 1 0 68320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1666464484
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_605
timestamp 1666464484
transform 1 0 69104 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_669
timestamp 1666464484
transform 1 0 76272 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1666464484
transform 1 0 76720 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_676
timestamp 1666464484
transform 1 0 77056 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_740
timestamp 1666464484
transform 1 0 84224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_744
timestamp 1666464484
transform 1 0 84672 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_747
timestamp 1666464484
transform 1 0 85008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_811
timestamp 1666464484
transform 1 0 92176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_815
timestamp 1666464484
transform 1 0 92624 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_818
timestamp 1666464484
transform 1 0 92960 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_882
timestamp 1666464484
transform 1 0 100128 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_886
timestamp 1666464484
transform 1 0 100576 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_889
timestamp 1666464484
transform 1 0 100912 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_953
timestamp 1666464484
transform 1 0 108080 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_957
timestamp 1666464484
transform 1 0 108528 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_960
timestamp 1666464484
transform 1 0 108864 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1024
timestamp 1666464484
transform 1 0 116032 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1028
timestamp 1666464484
transform 1 0 116480 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1031
timestamp 1666464484
transform 1 0 116816 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1095
timestamp 1666464484
transform 1 0 123984 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1099
timestamp 1666464484
transform 1 0 124432 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1102
timestamp 1666464484
transform 1 0 124768 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1166
timestamp 1666464484
transform 1 0 131936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1170
timestamp 1666464484
transform 1 0 132384 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1173
timestamp 1666464484
transform 1 0 132720 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1237
timestamp 1666464484
transform 1 0 139888 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1241
timestamp 1666464484
transform 1 0 140336 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1244
timestamp 1666464484
transform 1 0 140672 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1308
timestamp 1666464484
transform 1 0 147840 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1312
timestamp 1666464484
transform 1 0 148288 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1666464484
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1666464484
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1666464484
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1666464484
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1666464484
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1666464484
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1666464484
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1666464484
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1666464484
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1666464484
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1666464484
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1666464484
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1666464484
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1666464484
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1666464484
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1666464484
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1666464484
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1666464484
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1666464484
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1666464484
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1666464484
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1666464484
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1666464484
transform 1 0 64400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1666464484
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1666464484
transform 1 0 65184 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1666464484
transform 1 0 72352 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1666464484
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_641
timestamp 1666464484
transform 1 0 73136 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_705
timestamp 1666464484
transform 1 0 80304 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_709
timestamp 1666464484
transform 1 0 80752 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_712
timestamp 1666464484
transform 1 0 81088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_776
timestamp 1666464484
transform 1 0 88256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_780
timestamp 1666464484
transform 1 0 88704 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_783
timestamp 1666464484
transform 1 0 89040 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_847
timestamp 1666464484
transform 1 0 96208 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_851
timestamp 1666464484
transform 1 0 96656 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_854
timestamp 1666464484
transform 1 0 96992 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_918
timestamp 1666464484
transform 1 0 104160 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_922
timestamp 1666464484
transform 1 0 104608 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_925
timestamp 1666464484
transform 1 0 104944 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_989
timestamp 1666464484
transform 1 0 112112 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_993
timestamp 1666464484
transform 1 0 112560 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_996
timestamp 1666464484
transform 1 0 112896 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1060
timestamp 1666464484
transform 1 0 120064 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1064
timestamp 1666464484
transform 1 0 120512 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1067
timestamp 1666464484
transform 1 0 120848 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1131
timestamp 1666464484
transform 1 0 128016 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1135
timestamp 1666464484
transform 1 0 128464 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1138
timestamp 1666464484
transform 1 0 128800 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1202
timestamp 1666464484
transform 1 0 135968 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1206
timestamp 1666464484
transform 1 0 136416 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1209
timestamp 1666464484
transform 1 0 136752 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1273
timestamp 1666464484
transform 1 0 143920 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1277
timestamp 1666464484
transform 1 0 144368 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_1280
timestamp 1666464484
transform 1 0 144704 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1312
timestamp 1666464484
transform 1 0 148288 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1666464484
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1666464484
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1666464484
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1666464484
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1666464484
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1666464484
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1666464484
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1666464484
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1666464484
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1666464484
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1666464484
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1666464484
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1666464484
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1666464484
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1666464484
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1666464484
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1666464484
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1666464484
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1666464484
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1666464484
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1666464484
transform 1 0 53200 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1666464484
transform 1 0 60368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1666464484
transform 1 0 60816 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1666464484
transform 1 0 61152 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_598
timestamp 1666464484
transform 1 0 68320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1666464484
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1666464484
transform 1 0 69104 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_669
timestamp 1666464484
transform 1 0 76272 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1666464484
transform 1 0 76720 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_676
timestamp 1666464484
transform 1 0 77056 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_740
timestamp 1666464484
transform 1 0 84224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_744
timestamp 1666464484
transform 1 0 84672 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_747
timestamp 1666464484
transform 1 0 85008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_811
timestamp 1666464484
transform 1 0 92176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_815
timestamp 1666464484
transform 1 0 92624 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_818
timestamp 1666464484
transform 1 0 92960 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_882
timestamp 1666464484
transform 1 0 100128 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_886
timestamp 1666464484
transform 1 0 100576 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_889
timestamp 1666464484
transform 1 0 100912 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_953
timestamp 1666464484
transform 1 0 108080 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_957
timestamp 1666464484
transform 1 0 108528 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_960
timestamp 1666464484
transform 1 0 108864 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1024
timestamp 1666464484
transform 1 0 116032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1028
timestamp 1666464484
transform 1 0 116480 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1031
timestamp 1666464484
transform 1 0 116816 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1095
timestamp 1666464484
transform 1 0 123984 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1099
timestamp 1666464484
transform 1 0 124432 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1102
timestamp 1666464484
transform 1 0 124768 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1166
timestamp 1666464484
transform 1 0 131936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1170
timestamp 1666464484
transform 1 0 132384 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1173
timestamp 1666464484
transform 1 0 132720 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1237
timestamp 1666464484
transform 1 0 139888 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1241
timestamp 1666464484
transform 1 0 140336 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1244
timestamp 1666464484
transform 1 0 140672 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1308
timestamp 1666464484
transform 1 0 147840 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1312
timestamp 1666464484
transform 1 0 148288 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1666464484
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1666464484
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1666464484
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1666464484
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1666464484
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1666464484
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1666464484
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1666464484
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1666464484
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1666464484
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1666464484
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1666464484
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1666464484
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1666464484
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1666464484
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1666464484
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1666464484
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1666464484
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_428
timestamp 1666464484
transform 1 0 49280 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_460
timestamp 1666464484
transform 1 0 52864 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_466
timestamp 1666464484
transform 1 0 53536 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_482
timestamp 1666464484
transform 1 0 55328 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_490
timestamp 1666464484
transform 1 0 56224 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_494
timestamp 1666464484
transform 1 0 56672 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1666464484
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_499
timestamp 1666464484
transform 1 0 57232 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_531
timestamp 1666464484
transform 1 0 60816 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_539
timestamp 1666464484
transform 1 0 61712 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_543
timestamp 1666464484
transform 1 0 62160 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_547
timestamp 1666464484
transform 1 0 62608 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_551
timestamp 1666464484
transform 1 0 63056 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1666464484
transform 1 0 64848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1666464484
transform 1 0 65184 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_634
timestamp 1666464484
transform 1 0 72352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1666464484
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_641
timestamp 1666464484
transform 1 0 73136 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_705
timestamp 1666464484
transform 1 0 80304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_709
timestamp 1666464484
transform 1 0 80752 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_712
timestamp 1666464484
transform 1 0 81088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_776
timestamp 1666464484
transform 1 0 88256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_780
timestamp 1666464484
transform 1 0 88704 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_783
timestamp 1666464484
transform 1 0 89040 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_847
timestamp 1666464484
transform 1 0 96208 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_851
timestamp 1666464484
transform 1 0 96656 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_854
timestamp 1666464484
transform 1 0 96992 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_918
timestamp 1666464484
transform 1 0 104160 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_922
timestamp 1666464484
transform 1 0 104608 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_925
timestamp 1666464484
transform 1 0 104944 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_941
timestamp 1666464484
transform 1 0 106736 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_949
timestamp 1666464484
transform 1 0 107632 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_955
timestamp 1666464484
transform 1 0 108304 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_987
timestamp 1666464484
transform 1 0 111888 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_991
timestamp 1666464484
transform 1 0 112336 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_993
timestamp 1666464484
transform 1 0 112560 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_996
timestamp 1666464484
transform 1 0 112896 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1060
timestamp 1666464484
transform 1 0 120064 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1064
timestamp 1666464484
transform 1 0 120512 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1067
timestamp 1666464484
transform 1 0 120848 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1131
timestamp 1666464484
transform 1 0 128016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1135
timestamp 1666464484
transform 1 0 128464 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1138
timestamp 1666464484
transform 1 0 128800 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1202
timestamp 1666464484
transform 1 0 135968 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1206
timestamp 1666464484
transform 1 0 136416 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1209
timestamp 1666464484
transform 1 0 136752 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1273
timestamp 1666464484
transform 1 0 143920 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1277
timestamp 1666464484
transform 1 0 144368 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_1280
timestamp 1666464484
transform 1 0 144704 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1312
timestamp 1666464484
transform 1 0 148288 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1666464484
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1666464484
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1666464484
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1666464484
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1666464484
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_108
timestamp 1666464484
transform 1 0 13440 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_140
timestamp 1666464484
transform 1 0 17024 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_142
timestamp 1666464484
transform 1 0 17248 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_145
timestamp 1666464484
transform 1 0 17584 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_149
timestamp 1666464484
transform 1 0 18032 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_151
timestamp 1666464484
transform 1 0 18256 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_154
timestamp 1666464484
transform 1 0 18592 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_158
timestamp 1666464484
transform 1 0 19040 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_162
timestamp 1666464484
transform 1 0 19488 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_166
timestamp 1666464484
transform 1 0 19936 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_170
timestamp 1666464484
transform 1 0 20384 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_174
timestamp 1666464484
transform 1 0 20832 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1666464484
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1666464484
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1666464484
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1666464484
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_250
timestamp 1666464484
transform 1 0 29344 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_258
timestamp 1666464484
transform 1 0 30240 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_262
timestamp 1666464484
transform 1 0 30688 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_266
timestamp 1666464484
transform 1 0 31136 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_298
timestamp 1666464484
transform 1 0 34720 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1666464484
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1666464484
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_321
timestamp 1666464484
transform 1 0 37296 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_325
timestamp 1666464484
transform 1 0 37744 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_329
timestamp 1666464484
transform 1 0 38192 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_333
timestamp 1666464484
transform 1 0 38640 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_365
timestamp 1666464484
transform 1 0 42224 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_381
timestamp 1666464484
transform 1 0 44016 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1666464484
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_392
timestamp 1666464484
transform 1 0 45248 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_400
timestamp 1666464484
transform 1 0 46144 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_403
timestamp 1666464484
transform 1 0 46480 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_407
timestamp 1666464484
transform 1 0 46928 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_423
timestamp 1666464484
transform 1 0 48720 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_429
timestamp 1666464484
transform 1 0 49392 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_445
timestamp 1666464484
transform 1 0 51184 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_449
timestamp 1666464484
transform 1 0 51632 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_451
timestamp 1666464484
transform 1 0 51856 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_454
timestamp 1666464484
transform 1 0 52192 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1666464484
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_463
timestamp 1666464484
transform 1 0 53200 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_466
timestamp 1666464484
transform 1 0 53536 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_470
timestamp 1666464484
transform 1 0 53984 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_472
timestamp 1666464484
transform 1 0 54208 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_475
timestamp 1666464484
transform 1 0 54544 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_507
timestamp 1666464484
transform 1 0 58128 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_515
timestamp 1666464484
transform 1 0 59024 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_518
timestamp 1666464484
transform 1 0 59360 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_522
timestamp 1666464484
transform 1 0 59808 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_524
timestamp 1666464484
transform 1 0 60032 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_527
timestamp 1666464484
transform 1 0 60368 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1666464484
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_534
timestamp 1666464484
transform 1 0 61152 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_540
timestamp 1666464484
transform 1 0 61824 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_548
timestamp 1666464484
transform 1 0 62720 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_552
timestamp 1666464484
transform 1 0 63168 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_558
timestamp 1666464484
transform 1 0 63840 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_562
timestamp 1666464484
transform 1 0 64288 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_566
timestamp 1666464484
transform 1 0 64736 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_570
timestamp 1666464484
transform 1 0 65184 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_572
timestamp 1666464484
transform 1 0 65408 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_575
timestamp 1666464484
transform 1 0 65744 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_591
timestamp 1666464484
transform 1 0 67536 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_599
timestamp 1666464484
transform 1 0 68432 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_605
timestamp 1666464484
transform 1 0 69104 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_637
timestamp 1666464484
transform 1 0 72688 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_645
timestamp 1666464484
transform 1 0 73584 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_648
timestamp 1666464484
transform 1 0 73920 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_652
timestamp 1666464484
transform 1 0 74368 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_656
timestamp 1666464484
transform 1 0 74816 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_664
timestamp 1666464484
transform 1 0 75712 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_668
timestamp 1666464484
transform 1 0 76160 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_672
timestamp 1666464484
transform 1 0 76608 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_676
timestamp 1666464484
transform 1 0 77056 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_740
timestamp 1666464484
transform 1 0 84224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_744
timestamp 1666464484
transform 1 0 84672 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_747
timestamp 1666464484
transform 1 0 85008 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_763
timestamp 1666464484
transform 1 0 86800 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_771
timestamp 1666464484
transform 1 0 87696 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_774
timestamp 1666464484
transform 1 0 88032 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_784
timestamp 1666464484
transform 1 0 89152 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_788
timestamp 1666464484
transform 1 0 89600 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_804
timestamp 1666464484
transform 1 0 91392 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_808
timestamp 1666464484
transform 1 0 91840 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_818
timestamp 1666464484
transform 1 0 92960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_821
timestamp 1666464484
transform 1 0 93296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_885
timestamp 1666464484
transform 1 0 100464 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_889
timestamp 1666464484
transform 1 0 100912 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_921
timestamp 1666464484
transform 1 0 104496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_927
timestamp 1666464484
transform 1 0 105168 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_931
timestamp 1666464484
transform 1 0 105616 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_934
timestamp 1666464484
transform 1 0 105952 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_938
timestamp 1666464484
transform 1 0 106400 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_942
timestamp 1666464484
transform 1 0 106848 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_946
timestamp 1666464484
transform 1 0 107296 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_950
timestamp 1666464484
transform 1 0 107744 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_954
timestamp 1666464484
transform 1 0 108192 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_960
timestamp 1666464484
transform 1 0 108864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_963
timestamp 1666464484
transform 1 0 109200 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_967
timestamp 1666464484
transform 1 0 109648 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_969
timestamp 1666464484
transform 1 0 109872 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_972
timestamp 1666464484
transform 1 0 110208 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_976
timestamp 1666464484
transform 1 0 110656 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_980
timestamp 1666464484
transform 1 0 111104 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_1012
timestamp 1666464484
transform 1 0 114688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1028
timestamp 1666464484
transform 1 0 116480 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1031
timestamp 1666464484
transform 1 0 116816 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1095
timestamp 1666464484
transform 1 0 123984 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1099
timestamp 1666464484
transform 1 0 124432 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_1102
timestamp 1666464484
transform 1 0 124768 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1110
timestamp 1666464484
transform 1 0 125664 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1114
timestamp 1666464484
transform 1 0 126112 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1116
timestamp 1666464484
transform 1 0 126336 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1119
timestamp 1666464484
transform 1 0 126672 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_1123
timestamp 1666464484
transform 1 0 127120 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1131
timestamp 1666464484
transform 1 0 128016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1135
timestamp 1666464484
transform 1 0 128464 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1139
timestamp 1666464484
transform 1 0 128912 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1147
timestamp 1666464484
transform 1 0 129808 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1151
timestamp 1666464484
transform 1 0 130256 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1155
timestamp 1666464484
transform 1 0 130704 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1159
timestamp 1666464484
transform 1 0 131152 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_1163
timestamp 1666464484
transform 1 0 131600 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1173
timestamp 1666464484
transform 1 0 132720 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1237
timestamp 1666464484
transform 1 0 139888 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1241
timestamp 1666464484
transform 1 0 140336 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1244
timestamp 1666464484
transform 1 0 140672 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1308
timestamp 1666464484
transform 1 0 147840 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1312
timestamp 1666464484
transform 1 0 148288 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_2
timestamp 1666464484
transform 1 0 1568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_34
timestamp 1666464484
transform 1 0 5152 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_50
timestamp 1666464484
transform 1 0 6944 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_56
timestamp 1666464484
transform 1 0 7616 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_60
timestamp 1666464484
transform 1 0 8064 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_68
timestamp 1666464484
transform 1 0 8960 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1666464484
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_73
timestamp 1666464484
transform 1 0 9520 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_76
timestamp 1666464484
transform 1 0 9856 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_92
timestamp 1666464484
transform 1 0 11648 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_96
timestamp 1666464484
transform 1 0 12096 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_99
timestamp 1666464484
transform 1 0 12432 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_107
timestamp 1666464484
transform 1 0 13328 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_110
timestamp 1666464484
transform 1 0 13664 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_118
timestamp 1666464484
transform 1 0 14560 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_122
timestamp 1666464484
transform 1 0 15008 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_126
timestamp 1666464484
transform 1 0 15456 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_130
timestamp 1666464484
transform 1 0 15904 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_134
timestamp 1666464484
transform 1 0 16352 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_137
timestamp 1666464484
transform 1 0 16688 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1666464484
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_144
timestamp 1666464484
transform 1 0 17472 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_154
timestamp 1666464484
transform 1 0 18592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_164
timestamp 1666464484
transform 1 0 19712 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_172
timestamp 1666464484
transform 1 0 20608 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_180
timestamp 1666464484
transform 1 0 21504 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_184
timestamp 1666464484
transform 1 0 21952 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_190
timestamp 1666464484
transform 1 0 22624 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_194
timestamp 1666464484
transform 1 0 23072 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_198
timestamp 1666464484
transform 1 0 23520 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_202
timestamp 1666464484
transform 1 0 23968 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_206
timestamp 1666464484
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_210
timestamp 1666464484
transform 1 0 24864 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1666464484
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_215
timestamp 1666464484
transform 1 0 25424 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_218
timestamp 1666464484
transform 1 0 25760 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_222
timestamp 1666464484
transform 1 0 26208 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_232
timestamp 1666464484
transform 1 0 27328 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_236
timestamp 1666464484
transform 1 0 27776 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_244
timestamp 1666464484
transform 1 0 28672 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_248
timestamp 1666464484
transform 1 0 29120 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_252
timestamp 1666464484
transform 1 0 29568 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_256
timestamp 1666464484
transform 1 0 30016 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_260
timestamp 1666464484
transform 1 0 30464 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_268
timestamp 1666464484
transform 1 0 31360 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_272
timestamp 1666464484
transform 1 0 31808 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_276
timestamp 1666464484
transform 1 0 32256 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1666464484
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1666464484
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_286
timestamp 1666464484
transform 1 0 33376 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_289
timestamp 1666464484
transform 1 0 33712 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_295
timestamp 1666464484
transform 1 0 34384 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_299
timestamp 1666464484
transform 1 0 34832 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_303
timestamp 1666464484
transform 1 0 35280 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_307
timestamp 1666464484
transform 1 0 35728 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_309
timestamp 1666464484
transform 1 0 35952 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_312
timestamp 1666464484
transform 1 0 36288 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_316
timestamp 1666464484
transform 1 0 36736 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_319
timestamp 1666464484
transform 1 0 37072 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_327
timestamp 1666464484
transform 1 0 37968 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_331
timestamp 1666464484
transform 1 0 38416 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_334
timestamp 1666464484
transform 1 0 38752 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_342
timestamp 1666464484
transform 1 0 39648 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_346
timestamp 1666464484
transform 1 0 40096 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_352
timestamp 1666464484
transform 1 0 40768 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1666464484
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_357
timestamp 1666464484
transform 1 0 41328 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_360
timestamp 1666464484
transform 1 0 41664 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_364
timestamp 1666464484
transform 1 0 42112 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_368
timestamp 1666464484
transform 1 0 42560 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_370
timestamp 1666464484
transform 1 0 42784 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_373
timestamp 1666464484
transform 1 0 43120 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_381
timestamp 1666464484
transform 1 0 44016 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_385
timestamp 1666464484
transform 1 0 44464 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_389
timestamp 1666464484
transform 1 0 44912 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_393
timestamp 1666464484
transform 1 0 45360 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_401
timestamp 1666464484
transform 1 0 46256 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_409
timestamp 1666464484
transform 1 0 47152 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_413
timestamp 1666464484
transform 1 0 47600 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_417
timestamp 1666464484
transform 1 0 48048 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_420
timestamp 1666464484
transform 1 0 48384 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_422
timestamp 1666464484
transform 1 0 48608 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1666464484
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_428
timestamp 1666464484
transform 1 0 49280 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_436
timestamp 1666464484
transform 1 0 50176 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_440
timestamp 1666464484
transform 1 0 50624 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_443
timestamp 1666464484
transform 1 0 50960 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_447
timestamp 1666464484
transform 1 0 51408 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_451
timestamp 1666464484
transform 1 0 51856 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_459
timestamp 1666464484
transform 1 0 52752 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_467
timestamp 1666464484
transform 1 0 53648 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_471
timestamp 1666464484
transform 1 0 54096 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_474
timestamp 1666464484
transform 1 0 54432 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_478
timestamp 1666464484
transform 1 0 54880 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_482
timestamp 1666464484
transform 1 0 55328 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_484
timestamp 1666464484
transform 1 0 55552 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_487
timestamp 1666464484
transform 1 0 55888 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_491
timestamp 1666464484
transform 1 0 56336 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_495
timestamp 1666464484
transform 1 0 56784 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_499
timestamp 1666464484
transform 1 0 57232 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_502
timestamp 1666464484
transform 1 0 57568 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_506
timestamp 1666464484
transform 1 0 58016 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_510
timestamp 1666464484
transform 1 0 58464 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_514
timestamp 1666464484
transform 1 0 58912 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_518
timestamp 1666464484
transform 1 0 59360 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_520
timestamp 1666464484
transform 1 0 59584 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_523
timestamp 1666464484
transform 1 0 59920 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_527
timestamp 1666464484
transform 1 0 60368 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_531
timestamp 1666464484
transform 1 0 60816 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_541
timestamp 1666464484
transform 1 0 61936 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_549
timestamp 1666464484
transform 1 0 62832 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_551
timestamp 1666464484
transform 1 0 63056 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_560
timestamp 1666464484
transform 1 0 64064 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_566
timestamp 1666464484
transform 1 0 64736 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_570
timestamp 1666464484
transform 1 0 65184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_573
timestamp 1666464484
transform 1 0 65520 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_577
timestamp 1666464484
transform 1 0 65968 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_579
timestamp 1666464484
transform 1 0 66192 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_582
timestamp 1666464484
transform 1 0 66528 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_592
timestamp 1666464484
transform 1 0 67648 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_596
timestamp 1666464484
transform 1 0 68096 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_606
timestamp 1666464484
transform 1 0 69216 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_622
timestamp 1666464484
transform 1 0 71008 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_630
timestamp 1666464484
transform 1 0 71904 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_634
timestamp 1666464484
transform 1 0 72352 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1666464484
transform 1 0 72800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_641
timestamp 1666464484
transform 1 0 73136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_644
timestamp 1666464484
transform 1 0 73472 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_650
timestamp 1666464484
transform 1 0 74144 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_654
timestamp 1666464484
transform 1 0 74592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_660
timestamp 1666464484
transform 1 0 75264 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_666
timestamp 1666464484
transform 1 0 75936 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_670
timestamp 1666464484
transform 1 0 76384 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_674
timestamp 1666464484
transform 1 0 76832 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_678
timestamp 1666464484
transform 1 0 77280 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_682
timestamp 1666464484
transform 1 0 77728 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_684
timestamp 1666464484
transform 1 0 77952 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_687
timestamp 1666464484
transform 1 0 78288 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_689
timestamp 1666464484
transform 1 0 78512 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_692
timestamp 1666464484
transform 1 0 78848 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_700
timestamp 1666464484
transform 1 0 79744 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_708
timestamp 1666464484
transform 1 0 80640 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_712
timestamp 1666464484
transform 1 0 81088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_715
timestamp 1666464484
transform 1 0 81424 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_719
timestamp 1666464484
transform 1 0 81872 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_721
timestamp 1666464484
transform 1 0 82096 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_724
timestamp 1666464484
transform 1 0 82432 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_732
timestamp 1666464484
transform 1 0 83328 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_738
timestamp 1666464484
transform 1 0 84000 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_742
timestamp 1666464484
transform 1 0 84448 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_750
timestamp 1666464484
transform 1 0 85344 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_754
timestamp 1666464484
transform 1 0 85792 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_758
timestamp 1666464484
transform 1 0 86240 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_760
timestamp 1666464484
transform 1 0 86464 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_763
timestamp 1666464484
transform 1 0 86800 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_767
timestamp 1666464484
transform 1 0 87248 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_770
timestamp 1666464484
transform 1 0 87584 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_780
timestamp 1666464484
transform 1 0 88704 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_783
timestamp 1666464484
transform 1 0 89040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_792
timestamp 1666464484
transform 1 0 90048 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_796
timestamp 1666464484
transform 1 0 90496 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_800
timestamp 1666464484
transform 1 0 90944 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_804
timestamp 1666464484
transform 1 0 91392 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_820
timestamp 1666464484
transform 1 0 93184 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_824
timestamp 1666464484
transform 1 0 93632 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_828
timestamp 1666464484
transform 1 0 94080 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_838
timestamp 1666464484
transform 1 0 95200 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_842
timestamp 1666464484
transform 1 0 95648 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_846
timestamp 1666464484
transform 1 0 96096 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_850
timestamp 1666464484
transform 1 0 96544 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_854
timestamp 1666464484
transform 1 0 96992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_857
timestamp 1666464484
transform 1 0 97328 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_889
timestamp 1666464484
transform 1 0 100912 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_897
timestamp 1666464484
transform 1 0 101808 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_901
timestamp 1666464484
transform 1 0 102256 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_903
timestamp 1666464484
transform 1 0 102480 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_906
timestamp 1666464484
transform 1 0 102816 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_910
timestamp 1666464484
transform 1 0 103264 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_913
timestamp 1666464484
transform 1 0 103600 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_917
timestamp 1666464484
transform 1 0 104048 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_919
timestamp 1666464484
transform 1 0 104272 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_922
timestamp 1666464484
transform 1 0 104608 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_925
timestamp 1666464484
transform 1 0 104944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_928
timestamp 1666464484
transform 1 0 105280 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_932
timestamp 1666464484
transform 1 0 105728 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_940
timestamp 1666464484
transform 1 0 106624 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_948
timestamp 1666464484
transform 1 0 107520 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_956
timestamp 1666464484
transform 1 0 108416 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_960
timestamp 1666464484
transform 1 0 108864 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_964
timestamp 1666464484
transform 1 0 109312 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_972
timestamp 1666464484
transform 1 0 110208 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_978
timestamp 1666464484
transform 1 0 110880 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_982
timestamp 1666464484
transform 1 0 111328 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_986
timestamp 1666464484
transform 1 0 111776 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_996
timestamp 1666464484
transform 1 0 112896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_999
timestamp 1666464484
transform 1 0 113232 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1007
timestamp 1666464484
transform 1 0 114128 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1011
timestamp 1666464484
transform 1 0 114576 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_1015
timestamp 1666464484
transform 1 0 115024 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1031
timestamp 1666464484
transform 1 0 116816 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1035
timestamp 1666464484
transform 1 0 117264 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_1039
timestamp 1666464484
transform 1 0 117712 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1047
timestamp 1666464484
transform 1 0 118608 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1051
timestamp 1666464484
transform 1 0 119056 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_1055
timestamp 1666464484
transform 1 0 119504 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1063
timestamp 1666464484
transform 1 0 120400 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_1067
timestamp 1666464484
transform 1 0 120848 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1075
timestamp 1666464484
transform 1 0 121744 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1077
timestamp 1666464484
transform 1 0 121968 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1080
timestamp 1666464484
transform 1 0 122304 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1084
timestamp 1666464484
transform 1 0 122752 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1088
timestamp 1666464484
transform 1 0 123200 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_1092
timestamp 1666464484
transform 1 0 123648 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1100
timestamp 1666464484
transform 1 0 124544 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1103
timestamp 1666464484
transform 1 0 124880 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1107
timestamp 1666464484
transform 1 0 125328 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1111
timestamp 1666464484
transform 1 0 125776 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1119
timestamp 1666464484
transform 1 0 126672 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1123
timestamp 1666464484
transform 1 0 127120 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1127
timestamp 1666464484
transform 1 0 127568 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1131
timestamp 1666464484
transform 1 0 128016 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1135
timestamp 1666464484
transform 1 0 128464 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1138
timestamp 1666464484
transform 1 0 128800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1145
timestamp 1666464484
transform 1 0 129584 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1153
timestamp 1666464484
transform 1 0 130480 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1161
timestamp 1666464484
transform 1 0 131376 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1169
timestamp 1666464484
transform 1 0 132272 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1173
timestamp 1666464484
transform 1 0 132720 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_1177
timestamp 1666464484
transform 1 0 133168 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1187
timestamp 1666464484
transform 1 0 134288 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1191
timestamp 1666464484
transform 1 0 134736 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1193
timestamp 1666464484
transform 1 0 134960 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1196
timestamp 1666464484
transform 1 0 135296 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1200
timestamp 1666464484
transform 1 0 135744 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1204
timestamp 1666464484
transform 1 0 136192 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1206
timestamp 1666464484
transform 1 0 136416 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1209
timestamp 1666464484
transform 1 0 136752 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1215
timestamp 1666464484
transform 1 0 137424 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1221
timestamp 1666464484
transform 1 0 138096 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1225
timestamp 1666464484
transform 1 0 138544 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1229
timestamp 1666464484
transform 1 0 138992 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1233
timestamp 1666464484
transform 1 0 139440 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1235
timestamp 1666464484
transform 1 0 139664 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1238
timestamp 1666464484
transform 1 0 140000 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1240
timestamp 1666464484
transform 1 0 140224 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1243
timestamp 1666464484
transform 1 0 140560 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1247
timestamp 1666464484
transform 1 0 141008 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1249
timestamp 1666464484
transform 1 0 141232 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1252
timestamp 1666464484
transform 1 0 141568 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_1260
timestamp 1666464484
transform 1 0 142464 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_1270
timestamp 1666464484
transform 1 0 143584 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_1280
timestamp 1666464484
transform 1 0 144704 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1312
timestamp 1666464484
transform 1 0 148288 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1666464484
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1666464484
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_37
timestamp 1666464484
transform 1 0 5488 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_41
timestamp 1666464484
transform 1 0 5936 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_44
timestamp 1666464484
transform 1 0 6272 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_52
timestamp 1666464484
transform 1 0 7168 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_60
timestamp 1666464484
transform 1 0 8064 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_68
timestamp 1666464484
transform 1 0 8960 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_84
timestamp 1666464484
transform 1 0 10752 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_88
timestamp 1666464484
transform 1 0 11200 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_90
timestamp 1666464484
transform 1 0 11424 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_97
timestamp 1666464484
transform 1 0 12208 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1666464484
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_108
timestamp 1666464484
transform 1 0 13440 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_111
timestamp 1666464484
transform 1 0 13776 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_113
timestamp 1666464484
transform 1 0 14000 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_120
timestamp 1666464484
transform 1 0 14784 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_128
timestamp 1666464484
transform 1 0 15680 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_136
timestamp 1666464484
transform 1 0 16576 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_144
timestamp 1666464484
transform 1 0 17472 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_160
timestamp 1666464484
transform 1 0 19264 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1666464484
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_179
timestamp 1666464484
transform 1 0 21392 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_181
timestamp 1666464484
transform 1 0 21616 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_188
timestamp 1666464484
transform 1 0 22400 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_196
timestamp 1666464484
transform 1 0 23296 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_204
timestamp 1666464484
transform 1 0 24192 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_212
timestamp 1666464484
transform 1 0 25088 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_220
timestamp 1666464484
transform 1 0 25984 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_230
timestamp 1666464484
transform 1 0 27104 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_234
timestamp 1666464484
transform 1 0 27552 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_241
timestamp 1666464484
transform 1 0 28336 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_245
timestamp 1666464484
transform 1 0 28784 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1666464484
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_250
timestamp 1666464484
transform 1 0 29344 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_257
timestamp 1666464484
transform 1 0 30128 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_265
timestamp 1666464484
transform 1 0 31024 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_269
timestamp 1666464484
transform 1 0 31472 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_277
timestamp 1666464484
transform 1 0 32368 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_285
timestamp 1666464484
transform 1 0 33264 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_293
timestamp 1666464484
transform 1 0 34160 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_301
timestamp 1666464484
transform 1 0 35056 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_303
timestamp 1666464484
transform 1 0 35280 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_310
timestamp 1666464484
transform 1 0 36064 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1666464484
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_321
timestamp 1666464484
transform 1 0 37296 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_323
timestamp 1666464484
transform 1 0 37520 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_326
timestamp 1666464484
transform 1 0 37856 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_334
timestamp 1666464484
transform 1 0 38752 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_342
timestamp 1666464484
transform 1 0 39648 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_350
timestamp 1666464484
transform 1 0 40544 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_358
timestamp 1666464484
transform 1 0 41440 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_364
timestamp 1666464484
transform 1 0 42112 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_372
timestamp 1666464484
transform 1 0 43008 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_376
timestamp 1666464484
transform 1 0 43456 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_380
timestamp 1666464484
transform 1 0 43904 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_388
timestamp 1666464484
transform 1 0 44800 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_392
timestamp 1666464484
transform 1 0 45248 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_407
timestamp 1666464484
transform 1 0 46928 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_411
timestamp 1666464484
transform 1 0 47376 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_419
timestamp 1666464484
transform 1 0 48272 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_427
timestamp 1666464484
transform 1 0 49168 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_435
timestamp 1666464484
transform 1 0 50064 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_437
timestamp 1666464484
transform 1 0 50288 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_444
timestamp 1666464484
transform 1 0 51072 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_452
timestamp 1666464484
transform 1 0 51968 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1666464484
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_463
timestamp 1666464484
transform 1 0 53200 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_472
timestamp 1666464484
transform 1 0 54208 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_476
timestamp 1666464484
transform 1 0 54656 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_484
timestamp 1666464484
transform 1 0 55552 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_486
timestamp 1666464484
transform 1 0 55776 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_489
timestamp 1666464484
transform 1 0 56112 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_497
timestamp 1666464484
transform 1 0 57008 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_505
timestamp 1666464484
transform 1 0 57904 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_509
timestamp 1666464484
transform 1 0 58352 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_516
timestamp 1666464484
transform 1 0 59136 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_518
timestamp 1666464484
transform 1 0 59360 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_521
timestamp 1666464484
transform 1 0 59696 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_534
timestamp 1666464484
transform 1 0 61152 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_540
timestamp 1666464484
transform 1 0 61824 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_548
timestamp 1666464484
transform 1 0 62720 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_564
timestamp 1666464484
transform 1 0 64512 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_580
timestamp 1666464484
transform 1 0 66304 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_584
timestamp 1666464484
transform 1 0 66752 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_588
timestamp 1666464484
transform 1 0 67200 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_596
timestamp 1666464484
transform 1 0 68096 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1666464484
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_605
timestamp 1666464484
transform 1 0 69104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_612
timestamp 1666464484
transform 1 0 69888 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_616
timestamp 1666464484
transform 1 0 70336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_620
timestamp 1666464484
transform 1 0 70784 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_624
timestamp 1666464484
transform 1 0 71232 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_628
timestamp 1666464484
transform 1 0 71680 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_632
timestamp 1666464484
transform 1 0 72128 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_636
timestamp 1666464484
transform 1 0 72576 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_644
timestamp 1666464484
transform 1 0 73472 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_652
timestamp 1666464484
transform 1 0 74368 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_662
timestamp 1666464484
transform 1 0 75488 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_669
timestamp 1666464484
transform 1 0 76272 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1666464484
transform 1 0 76720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_676
timestamp 1666464484
transform 1 0 77056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_691
timestamp 1666464484
transform 1 0 78736 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_695
timestamp 1666464484
transform 1 0 79184 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_702
timestamp 1666464484
transform 1 0 79968 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_706
timestamp 1666464484
transform 1 0 80416 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_710
timestamp 1666464484
transform 1 0 80864 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_716
timestamp 1666464484
transform 1 0 81536 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_732
timestamp 1666464484
transform 1 0 83328 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_740
timestamp 1666464484
transform 1 0 84224 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_744
timestamp 1666464484
transform 1 0 84672 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_747
timestamp 1666464484
transform 1 0 85008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_754
timestamp 1666464484
transform 1 0 85792 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_758
timestamp 1666464484
transform 1 0 86240 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_762
timestamp 1666464484
transform 1 0 86688 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_769
timestamp 1666464484
transform 1 0 87472 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_773
timestamp 1666464484
transform 1 0 87920 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_788
timestamp 1666464484
transform 1 0 89600 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_804
timestamp 1666464484
transform 1 0 91392 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_808
timestamp 1666464484
transform 1 0 91840 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_815
timestamp 1666464484
transform 1 0 92624 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_818
timestamp 1666464484
transform 1 0 92960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_833
timestamp 1666464484
transform 1 0 94640 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_837
timestamp 1666464484
transform 1 0 95088 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_852
timestamp 1666464484
transform 1 0 96768 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_860
timestamp 1666464484
transform 1 0 97664 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_864
timestamp 1666464484
transform 1 0 98112 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_868
timestamp 1666464484
transform 1 0 98560 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_878
timestamp 1666464484
transform 1 0 99680 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_886
timestamp 1666464484
transform 1 0 100576 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_889
timestamp 1666464484
transform 1 0 100912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_892
timestamp 1666464484
transform 1 0 101248 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_896
timestamp 1666464484
transform 1 0 101696 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_904
timestamp 1666464484
transform 1 0 102592 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_912
timestamp 1666464484
transform 1 0 103488 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_916
timestamp 1666464484
transform 1 0 103936 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_924
timestamp 1666464484
transform 1 0 104832 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_940
timestamp 1666464484
transform 1 0 106624 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_956
timestamp 1666464484
transform 1 0 108416 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_960
timestamp 1666464484
transform 1 0 108864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_975
timestamp 1666464484
transform 1 0 110544 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_979
timestamp 1666464484
transform 1 0 110992 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_981
timestamp 1666464484
transform 1 0 111216 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_988
timestamp 1666464484
transform 1 0 112000 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_992
timestamp 1666464484
transform 1 0 112448 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_996
timestamp 1666464484
transform 1 0 112896 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1003
timestamp 1666464484
transform 1 0 113680 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1011
timestamp 1666464484
transform 1 0 114576 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1013
timestamp 1666464484
transform 1 0 114800 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1020
timestamp 1666464484
transform 1 0 115584 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1024
timestamp 1666464484
transform 1 0 116032 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1028
timestamp 1666464484
transform 1 0 116480 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1031
timestamp 1666464484
transform 1 0 116816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1034
timestamp 1666464484
transform 1 0 117152 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1038
timestamp 1666464484
transform 1 0 117600 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1045
timestamp 1666464484
transform 1 0 118384 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1053
timestamp 1666464484
transform 1 0 119280 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1061
timestamp 1666464484
transform 1 0 120176 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1065
timestamp 1666464484
transform 1 0 120624 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1069
timestamp 1666464484
transform 1 0 121072 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1071
timestamp 1666464484
transform 1 0 121296 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1078
timestamp 1666464484
transform 1 0 122080 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1086
timestamp 1666464484
transform 1 0 122976 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1094
timestamp 1666464484
transform 1 0 123872 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1098
timestamp 1666464484
transform 1 0 124320 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1102
timestamp 1666464484
transform 1 0 124768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1109
timestamp 1666464484
transform 1 0 125552 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1117
timestamp 1666464484
transform 1 0 126448 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1125
timestamp 1666464484
transform 1 0 127344 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1133
timestamp 1666464484
transform 1 0 128240 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1141
timestamp 1666464484
transform 1 0 129136 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1145
timestamp 1666464484
transform 1 0 129584 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1149
timestamp 1666464484
transform 1 0 130032 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1164
timestamp 1666464484
transform 1 0 131712 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1168
timestamp 1666464484
transform 1 0 132160 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1170
timestamp 1666464484
transform 1 0 132384 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1173
timestamp 1666464484
transform 1 0 132720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1180
timestamp 1666464484
transform 1 0 133504 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1184
timestamp 1666464484
transform 1 0 133952 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1186
timestamp 1666464484
transform 1 0 134176 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1193
timestamp 1666464484
transform 1 0 134960 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1197
timestamp 1666464484
transform 1 0 135408 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1212
timestamp 1666464484
transform 1 0 137088 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1228
timestamp 1666464484
transform 1 0 138880 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1232
timestamp 1666464484
transform 1 0 139328 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1234
timestamp 1666464484
transform 1 0 139552 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1241
timestamp 1666464484
transform 1 0 140336 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1244
timestamp 1666464484
transform 1 0 140672 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1251
timestamp 1666464484
transform 1 0 141456 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1255
timestamp 1666464484
transform 1 0 141904 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1262
timestamp 1666464484
transform 1 0 142688 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1266
timestamp 1666464484
transform 1 0 143136 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_1276
timestamp 1666464484
transform 1 0 144256 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1284
timestamp 1666464484
transform 1 0 145152 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1286
timestamp 1666464484
transform 1 0 145376 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_1289
timestamp 1666464484
transform 1 0 145712 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_1305
timestamp 1666464484
transform 1 0 147504 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_2
timestamp 1666464484
transform 1 0 1568 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_34
timestamp 1666464484
transform 1 0 5152 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_44
timestamp 1666464484
transform 1 0 6272 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_60
timestamp 1666464484
transform 1 0 8064 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1666464484
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_73
timestamp 1666464484
transform 1 0 9520 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_76
timestamp 1666464484
transform 1 0 9856 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_84
timestamp 1666464484
transform 1 0 10752 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_100
timestamp 1666464484
transform 1 0 12544 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_108
timestamp 1666464484
transform 1 0 13440 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_124
timestamp 1666464484
transform 1 0 15232 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_126
timestamp 1666464484
transform 1 0 15456 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1666464484
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_144
timestamp 1666464484
transform 1 0 17472 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_160
timestamp 1666464484
transform 1 0 19264 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_164
timestamp 1666464484
transform 1 0 19712 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_172
timestamp 1666464484
transform 1 0 20608 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_188
timestamp 1666464484
transform 1 0 22400 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_196
timestamp 1666464484
transform 1 0 23296 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1666464484
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_215
timestamp 1666464484
transform 1 0 25424 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_219
timestamp 1666464484
transform 1 0 25872 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_227
timestamp 1666464484
transform 1 0 26768 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_243
timestamp 1666464484
transform 1 0 28560 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_260
timestamp 1666464484
transform 1 0 30464 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_276
timestamp 1666464484
transform 1 0 32256 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_280
timestamp 1666464484
transform 1 0 32704 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_286
timestamp 1666464484
transform 1 0 33376 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_301
timestamp 1666464484
transform 1 0 35056 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_309
timestamp 1666464484
transform 1 0 35952 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_324
timestamp 1666464484
transform 1 0 37632 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_330
timestamp 1666464484
transform 1 0 38304 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_338
timestamp 1666464484
transform 1 0 39200 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_346
timestamp 1666464484
transform 1 0 40096 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1666464484
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_357
timestamp 1666464484
transform 1 0 41328 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_363
timestamp 1666464484
transform 1 0 42000 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_371
timestamp 1666464484
transform 1 0 42896 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_375
timestamp 1666464484
transform 1 0 43344 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_392
timestamp 1666464484
transform 1 0 45248 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_396
timestamp 1666464484
transform 1 0 45696 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_404
timestamp 1666464484
transform 1 0 46592 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_420
timestamp 1666464484
transform 1 0 48384 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_422
timestamp 1666464484
transform 1 0 48608 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1666464484
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_428
timestamp 1666464484
transform 1 0 49280 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_431
timestamp 1666464484
transform 1 0 49616 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_447
timestamp 1666464484
transform 1 0 51408 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_464
timestamp 1666464484
transform 1 0 53312 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_472
timestamp 1666464484
transform 1 0 54208 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_480
timestamp 1666464484
transform 1 0 55104 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1666464484
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_499
timestamp 1666464484
transform 1 0 57232 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_507
timestamp 1666464484
transform 1 0 58128 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_509
timestamp 1666464484
transform 1 0 58352 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_516
timestamp 1666464484
transform 1 0 59136 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_532
timestamp 1666464484
transform 1 0 60928 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_540
timestamp 1666464484
transform 1 0 61824 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_542
timestamp 1666464484
transform 1 0 62048 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_558
timestamp 1666464484
transform 1 0 63840 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_566
timestamp 1666464484
transform 1 0 64736 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_570
timestamp 1666464484
transform 1 0 65184 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_572
timestamp 1666464484
transform 1 0 65408 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_588
timestamp 1666464484
transform 1 0 67200 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_604
timestamp 1666464484
transform 1 0 68992 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_614
timestamp 1666464484
transform 1 0 70112 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_622
timestamp 1666464484
transform 1 0 71008 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1666464484
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_641
timestamp 1666464484
transform 1 0 73136 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_643
timestamp 1666464484
transform 1 0 73360 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_650
timestamp 1666464484
transform 1 0 74144 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_667
timestamp 1666464484
transform 1 0 76048 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_686
timestamp 1666464484
transform 1 0 78176 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_702
timestamp 1666464484
transform 1 0 79968 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_706
timestamp 1666464484
transform 1 0 80416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_712
timestamp 1666464484
transform 1 0 81088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_727
timestamp 1666464484
transform 1 0 82768 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_735
timestamp 1666464484
transform 1 0 83664 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_739
timestamp 1666464484
transform 1 0 84112 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_741
timestamp 1666464484
transform 1 0 84336 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_756
timestamp 1666464484
transform 1 0 86016 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_764
timestamp 1666464484
transform 1 0 86912 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_780
timestamp 1666464484
transform 1 0 88704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_783
timestamp 1666464484
transform 1 0 89040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_799
timestamp 1666464484
transform 1 0 90832 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_815
timestamp 1666464484
transform 1 0 92624 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_819
timestamp 1666464484
transform 1 0 93072 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_836
timestamp 1666464484
transform 1 0 94976 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_844
timestamp 1666464484
transform 1 0 95872 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_848
timestamp 1666464484
transform 1 0 96320 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_854
timestamp 1666464484
transform 1 0 96992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_857
timestamp 1666464484
transform 1 0 97328 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_861
timestamp 1666464484
transform 1 0 97776 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_876
timestamp 1666464484
transform 1 0 99456 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_884
timestamp 1666464484
transform 1 0 100352 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_888
timestamp 1666464484
transform 1 0 100800 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_892
timestamp 1666464484
transform 1 0 101248 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_900
timestamp 1666464484
transform 1 0 102144 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_916
timestamp 1666464484
transform 1 0 103936 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_920
timestamp 1666464484
transform 1 0 104384 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_922
timestamp 1666464484
transform 1 0 104608 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_925
timestamp 1666464484
transform 1 0 104944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_932
timestamp 1666464484
transform 1 0 105728 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_949
timestamp 1666464484
transform 1 0 107632 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_957
timestamp 1666464484
transform 1 0 108528 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_976
timestamp 1666464484
transform 1 0 110656 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_984
timestamp 1666464484
transform 1 0 111552 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_992
timestamp 1666464484
transform 1 0 112448 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_996
timestamp 1666464484
transform 1 0 112896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1003
timestamp 1666464484
transform 1 0 113680 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1005
timestamp 1666464484
transform 1 0 113904 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1020
timestamp 1666464484
transform 1 0 115584 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1028
timestamp 1666464484
transform 1 0 116480 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1036
timestamp 1666464484
transform 1 0 117376 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1052
timestamp 1666464484
transform 1 0 119168 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1060
timestamp 1666464484
transform 1 0 120064 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1064
timestamp 1666464484
transform 1 0 120512 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1067
timestamp 1666464484
transform 1 0 120848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1074
timestamp 1666464484
transform 1 0 121632 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1082
timestamp 1666464484
transform 1 0 122528 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1086
timestamp 1666464484
transform 1 0 122976 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1088
timestamp 1666464484
transform 1 0 123200 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1104
timestamp 1666464484
transform 1 0 124992 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1120
timestamp 1666464484
transform 1 0 126784 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1132
timestamp 1666464484
transform 1 0 128128 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1138
timestamp 1666464484
transform 1 0 128800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1147
timestamp 1666464484
transform 1 0 129808 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1151
timestamp 1666464484
transform 1 0 130256 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1153
timestamp 1666464484
transform 1 0 130480 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1169
timestamp 1666464484
transform 1 0 132272 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1177
timestamp 1666464484
transform 1 0 133168 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1181
timestamp 1666464484
transform 1 0 133616 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1196
timestamp 1666464484
transform 1 0 135296 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1204
timestamp 1666464484
transform 1 0 136192 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1206
timestamp 1666464484
transform 1 0 136416 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1209
timestamp 1666464484
transform 1 0 136752 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1212
timestamp 1666464484
transform 1 0 137088 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1214
timestamp 1666464484
transform 1 0 137312 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1221
timestamp 1666464484
transform 1 0 138096 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1238
timestamp 1666464484
transform 1 0 140000 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1255
timestamp 1666464484
transform 1 0 141904 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1259
timestamp 1666464484
transform 1 0 142352 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1261
timestamp 1666464484
transform 1 0 142576 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1276
timestamp 1666464484
transform 1 0 144256 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1280
timestamp 1666464484
transform 1 0 144704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1287
timestamp 1666464484
transform 1 0 145488 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1295
timestamp 1666464484
transform 1 0 146384 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_1299
timestamp 1666464484
transform 1 0 146832 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1307
timestamp 1666464484
transform 1 0 147728 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1311
timestamp 1666464484
transform 1 0 148176 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_2
timestamp 1666464484
transform 1 0 1568 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_18
timestamp 1666464484
transform 1 0 3360 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_26
timestamp 1666464484
transform 1 0 4256 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1666464484
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_37
timestamp 1666464484
transform 1 0 5488 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_52
timestamp 1666464484
transform 1 0 7168 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_68
timestamp 1666464484
transform 1 0 8960 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_72
timestamp 1666464484
transform 1 0 9408 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_88
timestamp 1666464484
transform 1 0 11200 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_104
timestamp 1666464484
transform 1 0 12992 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_107
timestamp 1666464484
transform 1 0 13328 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_123
timestamp 1666464484
transform 1 0 15120 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 16912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_142
timestamp 1666464484
transform 1 0 17248 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_145
timestamp 1666464484
transform 1 0 17584 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_153
timestamp 1666464484
transform 1 0 18480 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_170
timestamp 1666464484
transform 1 0 20384 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_174
timestamp 1666464484
transform 1 0 20832 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_177
timestamp 1666464484
transform 1 0 21168 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_193
timestamp 1666464484
transform 1 0 22960 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_209
timestamp 1666464484
transform 1 0 24752 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_212
timestamp 1666464484
transform 1 0 25088 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_228
timestamp 1666464484
transform 1 0 26880 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_244
timestamp 1666464484
transform 1 0 28672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1666464484
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_263
timestamp 1666464484
transform 1 0 30800 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_279
timestamp 1666464484
transform 1 0 32592 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_282
timestamp 1666464484
transform 1 0 32928 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_292
timestamp 1666464484
transform 1 0 34048 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_308
timestamp 1666464484
transform 1 0 35840 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_312
timestamp 1666464484
transform 1 0 36288 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_314
timestamp 1666464484
transform 1 0 36512 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_317
timestamp 1666464484
transform 1 0 36848 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_333
timestamp 1666464484
transform 1 0 38640 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_349
timestamp 1666464484
transform 1 0 40432 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_352
timestamp 1666464484
transform 1 0 40768 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_368
timestamp 1666464484
transform 1 0 42560 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_384
timestamp 1666464484
transform 1 0 44352 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_387
timestamp 1666464484
transform 1 0 44688 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_393
timestamp 1666464484
transform 1 0 45360 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_401
timestamp 1666464484
transform 1 0 46256 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_418
timestamp 1666464484
transform 1 0 48160 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_422
timestamp 1666464484
transform 1 0 48608 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_437
timestamp 1666464484
transform 1 0 50288 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_439
timestamp 1666464484
transform 1 0 50512 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_454
timestamp 1666464484
transform 1 0 52192 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_457
timestamp 1666464484
transform 1 0 52528 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_473
timestamp 1666464484
transform 1 0 54320 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_489
timestamp 1666464484
transform 1 0 56112 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_492
timestamp 1666464484
transform 1 0 56448 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_500
timestamp 1666464484
transform 1 0 57344 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_516
timestamp 1666464484
transform 1 0 59136 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_524
timestamp 1666464484
transform 1 0 60032 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_527
timestamp 1666464484
transform 1 0 60368 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_542
timestamp 1666464484
transform 1 0 62048 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_559
timestamp 1666464484
transform 1 0 63952 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_562
timestamp 1666464484
transform 1 0 64288 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_565
timestamp 1666464484
transform 1 0 64624 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_573
timestamp 1666464484
transform 1 0 65520 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_590
timestamp 1666464484
transform 1 0 67424 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_594
timestamp 1666464484
transform 1 0 67872 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_597
timestamp 1666464484
transform 1 0 68208 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_612
timestamp 1666464484
transform 1 0 69888 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_628
timestamp 1666464484
transform 1 0 71680 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_632
timestamp 1666464484
transform 1 0 72128 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_647
timestamp 1666464484
transform 1 0 73808 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_664
timestamp 1666464484
transform 1 0 75712 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_667
timestamp 1666464484
transform 1 0 76048 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_669
timestamp 1666464484
transform 1 0 76272 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_685
timestamp 1666464484
transform 1 0 78064 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_693
timestamp 1666464484
transform 1 0 78960 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_697
timestamp 1666464484
transform 1 0 79408 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_699
timestamp 1666464484
transform 1 0 79632 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_702
timestamp 1666464484
transform 1 0 79968 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_717
timestamp 1666464484
transform 1 0 81648 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_733
timestamp 1666464484
transform 1 0 83440 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_737
timestamp 1666464484
transform 1 0 83888 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_752
timestamp 1666464484
transform 1 0 85568 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_768
timestamp 1666464484
transform 1 0 87360 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_772
timestamp 1666464484
transform 1 0 87808 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_775
timestamp 1666464484
transform 1 0 88144 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_792
timestamp 1666464484
transform 1 0 90048 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_800
timestamp 1666464484
transform 1 0 90944 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_804
timestamp 1666464484
transform 1 0 91392 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_807
timestamp 1666464484
transform 1 0 91728 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_814
timestamp 1666464484
transform 1 0 92512 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_818
timestamp 1666464484
transform 1 0 92960 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_820
timestamp 1666464484
transform 1 0 93184 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_836
timestamp 1666464484
transform 1 0 94976 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_842
timestamp 1666464484
transform 1 0 95648 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_857
timestamp 1666464484
transform 1 0 97328 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_873
timestamp 1666464484
transform 1 0 99120 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_877
timestamp 1666464484
transform 1 0 99568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_892
timestamp 1666464484
transform 1 0 101248 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_908
timestamp 1666464484
transform 1 0 103040 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_912
timestamp 1666464484
transform 1 0 103488 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_927
timestamp 1666464484
transform 1 0 105168 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_944
timestamp 1666464484
transform 1 0 107072 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_947
timestamp 1666464484
transform 1 0 107408 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_950
timestamp 1666464484
transform 1 0 107744 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_954
timestamp 1666464484
transform 1 0 108192 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_970
timestamp 1666464484
transform 1 0 109984 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_978
timestamp 1666464484
transform 1 0 110880 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_982
timestamp 1666464484
transform 1 0 111328 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_997
timestamp 1666464484
transform 1 0 113008 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1013
timestamp 1666464484
transform 1 0 114800 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1017
timestamp 1666464484
transform 1 0 115248 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1020
timestamp 1666464484
transform 1 0 115584 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1036
timestamp 1666464484
transform 1 0 117376 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1044
timestamp 1666464484
transform 1 0 118272 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1048
timestamp 1666464484
transform 1 0 118720 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1052
timestamp 1666464484
transform 1 0 119168 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1068
timestamp 1666464484
transform 1 0 120960 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1084
timestamp 1666464484
transform 1 0 122752 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1087
timestamp 1666464484
transform 1 0 123088 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1103
timestamp 1666464484
transform 1 0 124880 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1119
timestamp 1666464484
transform 1 0 126672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1122
timestamp 1666464484
transform 1 0 127008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1137
timestamp 1666464484
transform 1 0 128688 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1153
timestamp 1666464484
transform 1 0 130480 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1157
timestamp 1666464484
transform 1 0 130928 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1173
timestamp 1666464484
transform 1 0 132720 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1189
timestamp 1666464484
transform 1 0 134512 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1192
timestamp 1666464484
transform 1 0 134848 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1195
timestamp 1666464484
transform 1 0 135184 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1197
timestamp 1666464484
transform 1 0 135408 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1213
timestamp 1666464484
transform 1 0 137200 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1221
timestamp 1666464484
transform 1 0 138096 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1227
timestamp 1666464484
transform 1 0 138768 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1243
timestamp 1666464484
transform 1 0 140560 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1259
timestamp 1666464484
transform 1 0 142352 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1262
timestamp 1666464484
transform 1 0 142688 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1277
timestamp 1666464484
transform 1 0 144368 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1293
timestamp 1666464484
transform 1 0 146160 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_1297
timestamp 1666464484
transform 1 0 146608 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1666464484
transform -1 0 148624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1666464484
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1666464484
transform -1 0 148624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1666464484
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1666464484
transform -1 0 148624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1666464484
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1666464484
transform -1 0 148624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1666464484
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1666464484
transform -1 0 148624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1666464484
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1666464484
transform -1 0 148624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1666464484
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1666464484
transform -1 0 148624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1666464484
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1666464484
transform -1 0 148624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1666464484
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1666464484
transform -1 0 148624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1666464484
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1666464484
transform -1 0 148624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1666464484
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1666464484
transform -1 0 148624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1666464484
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1666464484
transform -1 0 148624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1666464484
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1666464484
transform -1 0 148624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1666464484
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1666464484
transform -1 0 148624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1666464484
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1666464484
transform -1 0 148624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1666464484
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1666464484
transform -1 0 148624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1666464484
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1666464484
transform -1 0 148624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1666464484
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1666464484
transform -1 0 148624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1666464484
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1666464484
transform -1 0 148624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1666464484
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1666464484
transform -1 0 148624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1666464484
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1666464484
transform -1 0 148624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1666464484
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1666464484
transform -1 0 148624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1666464484
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1666464484
transform -1 0 148624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1666464484
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1666464484
transform -1 0 148624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1666464484
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1666464484
transform -1 0 148624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1666464484
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1666464484
transform -1 0 148624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1666464484
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1666464484
transform -1 0 148624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1666464484
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1666464484
transform -1 0 148624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1666464484
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1666464484
transform -1 0 148624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1666464484
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1666464484
transform -1 0 148624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1666464484
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1666464484
transform -1 0 148624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1666464484
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1666464484
transform -1 0 148624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1666464484
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1666464484
transform -1 0 148624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1666464484
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1666464484
transform -1 0 148624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1666464484
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1666464484
transform -1 0 148624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1666464484
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1666464484
transform -1 0 148624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1666464484
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1666464484
transform -1 0 148624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1666464484
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1666464484
transform -1 0 148624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1666464484
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1666464484
transform -1 0 148624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1666464484
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1666464484
transform -1 0 148624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1666464484
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1666464484
transform -1 0 148624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1666464484
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1666464484
transform -1 0 148624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1666464484
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1666464484
transform -1 0 148624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1666464484
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1666464484
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1666464484
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1666464484
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1666464484
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1666464484
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1666464484
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1666464484
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1666464484
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1666464484
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1666464484
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1666464484
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1666464484
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1666464484
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1666464484
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1666464484
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1666464484
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1666464484
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1666464484
transform 1 0 79744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1666464484
transform 1 0 83664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1666464484
transform 1 0 87584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1666464484
transform 1 0 91504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1666464484
transform 1 0 95424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1666464484
transform 1 0 99344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1666464484
transform 1 0 103264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1666464484
transform 1 0 107184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1666464484
transform 1 0 111104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1666464484
transform 1 0 115024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1666464484
transform 1 0 118944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1666464484
transform 1 0 122864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1666464484
transform 1 0 126784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1666464484
transform 1 0 130704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1666464484
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1666464484
transform 1 0 138544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1666464484
transform 1 0 142464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1666464484
transform 1 0 146384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1666464484
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1666464484
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1666464484
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1666464484
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1666464484
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1666464484
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1666464484
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1666464484
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1666464484
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1666464484
transform 1 0 80864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1666464484
transform 1 0 88816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1666464484
transform 1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1666464484
transform 1 0 104720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1666464484
transform 1 0 112672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1666464484
transform 1 0 120624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1666464484
transform 1 0 128576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1666464484
transform 1 0 136528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1666464484
transform 1 0 144480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1666464484
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1666464484
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1666464484
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1666464484
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1666464484
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1666464484
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1666464484
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1666464484
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1666464484
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1666464484
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1666464484
transform 1 0 84784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1666464484
transform 1 0 92736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1666464484
transform 1 0 100688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1666464484
transform 1 0 108640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1666464484
transform 1 0 116592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1666464484
transform 1 0 124544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1666464484
transform 1 0 132496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1666464484
transform 1 0 140448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1666464484
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1666464484
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1666464484
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1666464484
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1666464484
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1666464484
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1666464484
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1666464484
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1666464484
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1666464484
transform 1 0 80864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1666464484
transform 1 0 88816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1666464484
transform 1 0 96768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1666464484
transform 1 0 104720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1666464484
transform 1 0 112672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1666464484
transform 1 0 120624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1666464484
transform 1 0 128576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1666464484
transform 1 0 136528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1666464484
transform 1 0 144480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1666464484
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1666464484
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1666464484
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1666464484
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1666464484
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1666464484
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1666464484
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1666464484
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1666464484
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1666464484
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1666464484
transform 1 0 84784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1666464484
transform 1 0 92736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1666464484
transform 1 0 100688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1666464484
transform 1 0 108640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1666464484
transform 1 0 116592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1666464484
transform 1 0 124544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1666464484
transform 1 0 132496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1666464484
transform 1 0 140448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1666464484
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1666464484
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1666464484
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1666464484
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1666464484
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1666464484
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1666464484
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1666464484
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1666464484
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1666464484
transform 1 0 80864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1666464484
transform 1 0 88816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1666464484
transform 1 0 96768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1666464484
transform 1 0 104720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1666464484
transform 1 0 112672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1666464484
transform 1 0 120624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1666464484
transform 1 0 128576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1666464484
transform 1 0 136528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1666464484
transform 1 0 144480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1666464484
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1666464484
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1666464484
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1666464484
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1666464484
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1666464484
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1666464484
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1666464484
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1666464484
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1666464484
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1666464484
transform 1 0 84784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1666464484
transform 1 0 92736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1666464484
transform 1 0 100688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1666464484
transform 1 0 108640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1666464484
transform 1 0 116592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1666464484
transform 1 0 124544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1666464484
transform 1 0 132496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1666464484
transform 1 0 140448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1666464484
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1666464484
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1666464484
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1666464484
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1666464484
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1666464484
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1666464484
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1666464484
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1666464484
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1666464484
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1666464484
transform 1 0 88816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1666464484
transform 1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1666464484
transform 1 0 104720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1666464484
transform 1 0 112672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1666464484
transform 1 0 120624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1666464484
transform 1 0 128576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1666464484
transform 1 0 136528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1666464484
transform 1 0 144480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1666464484
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1666464484
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1666464484
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1666464484
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1666464484
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1666464484
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1666464484
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1666464484
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1666464484
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1666464484
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1666464484
transform 1 0 84784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1666464484
transform 1 0 92736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1666464484
transform 1 0 100688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1666464484
transform 1 0 108640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1666464484
transform 1 0 116592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1666464484
transform 1 0 124544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1666464484
transform 1 0 132496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1666464484
transform 1 0 140448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1666464484
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1666464484
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1666464484
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1666464484
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1666464484
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1666464484
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1666464484
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1666464484
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1666464484
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1666464484
transform 1 0 80864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1666464484
transform 1 0 88816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1666464484
transform 1 0 96768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1666464484
transform 1 0 104720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1666464484
transform 1 0 112672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1666464484
transform 1 0 120624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1666464484
transform 1 0 128576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1666464484
transform 1 0 136528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1666464484
transform 1 0 144480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1666464484
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1666464484
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1666464484
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1666464484
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1666464484
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1666464484
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1666464484
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1666464484
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1666464484
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1666464484
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1666464484
transform 1 0 84784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1666464484
transform 1 0 92736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1666464484
transform 1 0 100688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1666464484
transform 1 0 108640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1666464484
transform 1 0 116592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1666464484
transform 1 0 124544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1666464484
transform 1 0 132496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1666464484
transform 1 0 140448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1666464484
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1666464484
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1666464484
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1666464484
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1666464484
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1666464484
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1666464484
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1666464484
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1666464484
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1666464484
transform 1 0 80864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1666464484
transform 1 0 88816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1666464484
transform 1 0 96768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1666464484
transform 1 0 104720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1666464484
transform 1 0 112672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1666464484
transform 1 0 120624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1666464484
transform 1 0 128576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1666464484
transform 1 0 136528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1666464484
transform 1 0 144480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1666464484
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1666464484
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1666464484
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1666464484
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1666464484
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1666464484
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1666464484
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1666464484
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1666464484
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1666464484
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1666464484
transform 1 0 84784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1666464484
transform 1 0 92736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1666464484
transform 1 0 100688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1666464484
transform 1 0 108640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1666464484
transform 1 0 116592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1666464484
transform 1 0 124544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1666464484
transform 1 0 132496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1666464484
transform 1 0 140448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1666464484
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1666464484
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1666464484
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1666464484
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1666464484
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1666464484
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1666464484
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1666464484
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1666464484
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1666464484
transform 1 0 80864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1666464484
transform 1 0 88816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1666464484
transform 1 0 96768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1666464484
transform 1 0 104720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1666464484
transform 1 0 112672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1666464484
transform 1 0 120624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1666464484
transform 1 0 128576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1666464484
transform 1 0 136528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1666464484
transform 1 0 144480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1666464484
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1666464484
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1666464484
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1666464484
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1666464484
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1666464484
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1666464484
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1666464484
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1666464484
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1666464484
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1666464484
transform 1 0 84784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1666464484
transform 1 0 92736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1666464484
transform 1 0 100688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1666464484
transform 1 0 108640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1666464484
transform 1 0 116592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1666464484
transform 1 0 124544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1666464484
transform 1 0 132496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1666464484
transform 1 0 140448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1666464484
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1666464484
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1666464484
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1666464484
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1666464484
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1666464484
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1666464484
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1666464484
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1666464484
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1666464484
transform 1 0 80864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1666464484
transform 1 0 88816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1666464484
transform 1 0 96768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1666464484
transform 1 0 104720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1666464484
transform 1 0 112672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1666464484
transform 1 0 120624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1666464484
transform 1 0 128576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1666464484
transform 1 0 136528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1666464484
transform 1 0 144480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1666464484
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1666464484
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1666464484
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1666464484
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1666464484
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1666464484
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1666464484
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1666464484
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1666464484
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1666464484
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1666464484
transform 1 0 84784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1666464484
transform 1 0 92736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1666464484
transform 1 0 100688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1666464484
transform 1 0 108640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1666464484
transform 1 0 116592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1666464484
transform 1 0 124544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1666464484
transform 1 0 132496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1666464484
transform 1 0 140448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1666464484
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1666464484
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1666464484
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1666464484
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1666464484
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1666464484
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1666464484
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1666464484
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1666464484
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1666464484
transform 1 0 80864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1666464484
transform 1 0 88816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1666464484
transform 1 0 96768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1666464484
transform 1 0 104720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1666464484
transform 1 0 112672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1666464484
transform 1 0 120624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1666464484
transform 1 0 128576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1666464484
transform 1 0 136528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1666464484
transform 1 0 144480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1666464484
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1666464484
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1666464484
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1666464484
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1666464484
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1666464484
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1666464484
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1666464484
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1666464484
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1666464484
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1666464484
transform 1 0 84784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1666464484
transform 1 0 92736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1666464484
transform 1 0 100688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1666464484
transform 1 0 108640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1666464484
transform 1 0 116592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1666464484
transform 1 0 124544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1666464484
transform 1 0 132496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1666464484
transform 1 0 140448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1666464484
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1666464484
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1666464484
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1666464484
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1666464484
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1666464484
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1666464484
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1666464484
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1666464484
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1666464484
transform 1 0 80864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1666464484
transform 1 0 88816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1666464484
transform 1 0 96768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1666464484
transform 1 0 104720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1666464484
transform 1 0 112672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1666464484
transform 1 0 120624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1666464484
transform 1 0 128576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1666464484
transform 1 0 136528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1666464484
transform 1 0 144480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1666464484
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1666464484
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1666464484
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1666464484
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1666464484
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1666464484
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1666464484
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1666464484
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1666464484
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1666464484
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1666464484
transform 1 0 84784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1666464484
transform 1 0 92736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1666464484
transform 1 0 100688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1666464484
transform 1 0 108640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1666464484
transform 1 0 116592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1666464484
transform 1 0 124544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1666464484
transform 1 0 132496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1666464484
transform 1 0 140448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1666464484
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1666464484
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1666464484
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1666464484
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1666464484
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1666464484
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1666464484
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1666464484
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1666464484
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1666464484
transform 1 0 80864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1666464484
transform 1 0 88816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1666464484
transform 1 0 96768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1666464484
transform 1 0 104720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1666464484
transform 1 0 112672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1666464484
transform 1 0 120624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1666464484
transform 1 0 128576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1666464484
transform 1 0 136528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1666464484
transform 1 0 144480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1666464484
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1666464484
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1666464484
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1666464484
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1666464484
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1666464484
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1666464484
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1666464484
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1666464484
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1666464484
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1666464484
transform 1 0 84784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1666464484
transform 1 0 92736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1666464484
transform 1 0 100688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1666464484
transform 1 0 108640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1666464484
transform 1 0 116592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1666464484
transform 1 0 124544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1666464484
transform 1 0 132496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1666464484
transform 1 0 140448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1666464484
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1666464484
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1666464484
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1666464484
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1666464484
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1666464484
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1666464484
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1666464484
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1666464484
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1666464484
transform 1 0 80864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1666464484
transform 1 0 88816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1666464484
transform 1 0 96768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1666464484
transform 1 0 104720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1666464484
transform 1 0 112672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1666464484
transform 1 0 120624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1666464484
transform 1 0 128576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1666464484
transform 1 0 136528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1666464484
transform 1 0 144480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1666464484
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1666464484
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1666464484
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1666464484
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1666464484
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1666464484
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1666464484
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1666464484
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1666464484
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1666464484
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1666464484
transform 1 0 84784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1666464484
transform 1 0 92736 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1666464484
transform 1 0 100688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1666464484
transform 1 0 108640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1666464484
transform 1 0 116592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1666464484
transform 1 0 124544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1666464484
transform 1 0 132496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1666464484
transform 1 0 140448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1666464484
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1666464484
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1666464484
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1666464484
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1666464484
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1666464484
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1666464484
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1666464484
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1666464484
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1666464484
transform 1 0 80864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1666464484
transform 1 0 88816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1666464484
transform 1 0 96768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1666464484
transform 1 0 104720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1666464484
transform 1 0 112672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1666464484
transform 1 0 120624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1666464484
transform 1 0 128576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1666464484
transform 1 0 136528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1666464484
transform 1 0 144480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1666464484
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1666464484
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1666464484
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1666464484
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1666464484
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1666464484
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1666464484
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1666464484
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1666464484
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1666464484
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1666464484
transform 1 0 84784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1666464484
transform 1 0 92736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1666464484
transform 1 0 100688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1666464484
transform 1 0 108640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1666464484
transform 1 0 116592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1666464484
transform 1 0 124544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1666464484
transform 1 0 132496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1666464484
transform 1 0 140448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1666464484
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1666464484
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1666464484
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1666464484
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1666464484
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1666464484
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1666464484
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1666464484
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1666464484
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1666464484
transform 1 0 80864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1666464484
transform 1 0 88816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1666464484
transform 1 0 96768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1666464484
transform 1 0 104720 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1666464484
transform 1 0 112672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1666464484
transform 1 0 120624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1666464484
transform 1 0 128576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1666464484
transform 1 0 136528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1666464484
transform 1 0 144480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1666464484
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1666464484
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1666464484
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1666464484
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1666464484
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1666464484
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1666464484
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1666464484
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1666464484
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1666464484
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1666464484
transform 1 0 84784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1666464484
transform 1 0 92736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1666464484
transform 1 0 100688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1666464484
transform 1 0 108640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1666464484
transform 1 0 116592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1666464484
transform 1 0 124544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1666464484
transform 1 0 132496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1666464484
transform 1 0 140448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1666464484
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1666464484
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1666464484
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1666464484
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1666464484
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1666464484
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1666464484
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1666464484
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1666464484
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1666464484
transform 1 0 80864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1666464484
transform 1 0 88816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1666464484
transform 1 0 96768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1666464484
transform 1 0 104720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1666464484
transform 1 0 112672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1666464484
transform 1 0 120624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1666464484
transform 1 0 128576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1666464484
transform 1 0 136528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1666464484
transform 1 0 144480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1666464484
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1666464484
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1666464484
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1666464484
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1666464484
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1666464484
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1666464484
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1666464484
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1666464484
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1666464484
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1666464484
transform 1 0 84784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1666464484
transform 1 0 92736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1666464484
transform 1 0 100688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1666464484
transform 1 0 108640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1666464484
transform 1 0 116592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1666464484
transform 1 0 124544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1666464484
transform 1 0 132496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1666464484
transform 1 0 140448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1666464484
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1666464484
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1666464484
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1666464484
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1666464484
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1666464484
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1666464484
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1666464484
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1666464484
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1666464484
transform 1 0 80864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1666464484
transform 1 0 88816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1666464484
transform 1 0 96768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1666464484
transform 1 0 104720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1666464484
transform 1 0 112672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1666464484
transform 1 0 120624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1666464484
transform 1 0 128576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1666464484
transform 1 0 136528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1666464484
transform 1 0 144480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1666464484
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1666464484
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1666464484
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1666464484
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1666464484
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1666464484
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1666464484
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1666464484
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1666464484
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1666464484
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1666464484
transform 1 0 84784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1666464484
transform 1 0 92736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1666464484
transform 1 0 100688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1666464484
transform 1 0 108640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1666464484
transform 1 0 116592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1666464484
transform 1 0 124544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1666464484
transform 1 0 132496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1666464484
transform 1 0 140448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1666464484
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1666464484
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1666464484
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1666464484
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1666464484
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1666464484
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1666464484
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1666464484
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1666464484
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1666464484
transform 1 0 80864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1666464484
transform 1 0 88816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1666464484
transform 1 0 96768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1666464484
transform 1 0 104720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1666464484
transform 1 0 112672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1666464484
transform 1 0 120624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1666464484
transform 1 0 128576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1666464484
transform 1 0 136528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1666464484
transform 1 0 144480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1666464484
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1666464484
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1666464484
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1666464484
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1666464484
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1666464484
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1666464484
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1666464484
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1666464484
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1666464484
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1666464484
transform 1 0 84784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1666464484
transform 1 0 92736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1666464484
transform 1 0 100688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1666464484
transform 1 0 108640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1666464484
transform 1 0 116592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1666464484
transform 1 0 124544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1666464484
transform 1 0 132496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1666464484
transform 1 0 140448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1666464484
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1666464484
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1666464484
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1666464484
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1666464484
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1666464484
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1666464484
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1666464484
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1666464484
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1666464484
transform 1 0 80864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1666464484
transform 1 0 88816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1666464484
transform 1 0 96768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1666464484
transform 1 0 104720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1666464484
transform 1 0 112672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1666464484
transform 1 0 120624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1666464484
transform 1 0 128576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1666464484
transform 1 0 136528 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1666464484
transform 1 0 144480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1666464484
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1666464484
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1666464484
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1666464484
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1666464484
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1666464484
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1666464484
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1666464484
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1666464484
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1666464484
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1666464484
transform 1 0 84784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1666464484
transform 1 0 92736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1666464484
transform 1 0 100688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1666464484
transform 1 0 108640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1666464484
transform 1 0 116592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1666464484
transform 1 0 124544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1666464484
transform 1 0 132496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1666464484
transform 1 0 140448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1666464484
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1666464484
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1666464484
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1666464484
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1666464484
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1666464484
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1666464484
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1666464484
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1666464484
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1666464484
transform 1 0 80864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1666464484
transform 1 0 88816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1666464484
transform 1 0 96768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1666464484
transform 1 0 104720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1666464484
transform 1 0 112672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1666464484
transform 1 0 120624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1666464484
transform 1 0 128576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1666464484
transform 1 0 136528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1666464484
transform 1 0 144480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1666464484
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1666464484
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1666464484
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1666464484
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1666464484
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1666464484
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1666464484
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1666464484
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1666464484
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1666464484
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1666464484
transform 1 0 84784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1666464484
transform 1 0 92736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1666464484
transform 1 0 100688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1666464484
transform 1 0 108640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1666464484
transform 1 0 116592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1666464484
transform 1 0 124544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1666464484
transform 1 0 132496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1666464484
transform 1 0 140448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1666464484
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1666464484
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1666464484
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1666464484
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1666464484
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1666464484
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1666464484
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1666464484
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1666464484
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1666464484
transform 1 0 80864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1666464484
transform 1 0 88816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1666464484
transform 1 0 96768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1666464484
transform 1 0 104720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1666464484
transform 1 0 112672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1666464484
transform 1 0 120624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1666464484
transform 1 0 128576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1666464484
transform 1 0 136528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1666464484
transform 1 0 144480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1666464484
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1666464484
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1666464484
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1666464484
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1666464484
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1666464484
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1666464484
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1666464484
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1666464484
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1666464484
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1666464484
transform 1 0 84784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1666464484
transform 1 0 92736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1666464484
transform 1 0 100688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1666464484
transform 1 0 108640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1666464484
transform 1 0 116592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1666464484
transform 1 0 124544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1666464484
transform 1 0 132496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1666464484
transform 1 0 140448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1666464484
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1666464484
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1666464484
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1666464484
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1666464484
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1666464484
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1666464484
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1666464484
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1666464484
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1666464484
transform 1 0 80864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1666464484
transform 1 0 88816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1666464484
transform 1 0 96768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1666464484
transform 1 0 104720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1666464484
transform 1 0 112672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1666464484
transform 1 0 120624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1666464484
transform 1 0 128576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1666464484
transform 1 0 136528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1666464484
transform 1 0 144480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1666464484
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1666464484
transform 1 0 9184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1666464484
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1666464484
transform 1 0 17024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1666464484
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1666464484
transform 1 0 24864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1666464484
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1666464484
transform 1 0 32704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1666464484
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1666464484
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1666464484
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1666464484
transform 1 0 48384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1666464484
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1666464484
transform 1 0 56224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1666464484
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1666464484
transform 1 0 64064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1666464484
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1666464484
transform 1 0 71904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1666464484
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1666464484
transform 1 0 79744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1666464484
transform 1 0 83664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1666464484
transform 1 0 87584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1666464484
transform 1 0 91504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1666464484
transform 1 0 95424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1666464484
transform 1 0 99344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1666464484
transform 1 0 103264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1666464484
transform 1 0 107184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1666464484
transform 1 0 111104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1666464484
transform 1 0 115024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1666464484
transform 1 0 118944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1666464484
transform 1 0 122864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1666464484
transform 1 0 126784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1666464484
transform 1 0 130704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1666464484
transform 1 0 134624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1666464484
transform 1 0 138544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1666464484
transform 1 0 142464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1666464484
transform 1 0 146384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _168_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 61824 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _169_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 75712 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _170_
timestamp 1666464484
transform 1 0 39312 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _171_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 140336 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _172_
timestamp 1666464484
transform 1 0 123536 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _173_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 125552 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _174_
timestamp 1666464484
transform -1 0 76048 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _175_
timestamp 1666464484
transform 1 0 122192 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _176_
timestamp 1666464484
transform -1 0 122304 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _177_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 61040 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _178_
timestamp 1666464484
transform 1 0 128912 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _179_
timestamp 1666464484
transform -1 0 141904 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _180_
timestamp 1666464484
transform -1 0 138880 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _181_
timestamp 1666464484
transform -1 0 137648 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _182_
timestamp 1666464484
transform -1 0 140000 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _183_
timestamp 1666464484
transform -1 0 138096 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _184_
timestamp 1666464484
transform -1 0 136192 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _185_
timestamp 1666464484
transform -1 0 140560 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _186_
timestamp 1666464484
transform 1 0 140560 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _187_
timestamp 1666464484
transform -1 0 140000 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _188_
timestamp 1666464484
transform -1 0 137648 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _189_
timestamp 1666464484
transform -1 0 137200 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _190_
timestamp 1666464484
transform 1 0 136528 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _191_
timestamp 1666464484
transform -1 0 136304 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _192_
timestamp 1666464484
transform -1 0 128128 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _193_
timestamp 1666464484
transform -1 0 132272 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _194_
timestamp 1666464484
transform 1 0 131824 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _195_
timestamp 1666464484
transform 1 0 127008 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _196_
timestamp 1666464484
transform -1 0 132720 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _197_
timestamp 1666464484
transform 1 0 132832 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _198_
timestamp 1666464484
transform -1 0 130480 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _199_
timestamp 1666464484
transform 1 0 123312 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _200_
timestamp 1666464484
transform 1 0 110880 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _201_
timestamp 1666464484
transform -1 0 119168 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _202_
timestamp 1666464484
transform -1 0 119504 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _203_
timestamp 1666464484
transform 1 0 123200 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _204_
timestamp 1666464484
transform 1 0 115808 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _205_
timestamp 1666464484
transform -1 0 115248 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _206_
timestamp 1666464484
transform 1 0 62160 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _207_
timestamp 1666464484
transform 1 0 87808 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _208_
timestamp 1666464484
transform -1 0 110656 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _209_
timestamp 1666464484
transform 1 0 107856 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _210_
timestamp 1666464484
transform -1 0 107632 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _211_
timestamp 1666464484
transform -1 0 109984 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _212_
timestamp 1666464484
transform 1 0 108976 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _213_
timestamp 1666464484
transform -1 0 107744 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _214_
timestamp 1666464484
transform -1 0 107632 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _215_
timestamp 1666464484
transform 1 0 50848 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _216_
timestamp 1666464484
transform 1 0 92960 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _217_
timestamp 1666464484
transform 1 0 105168 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _218_
timestamp 1666464484
transform 1 0 103936 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _219_
timestamp 1666464484
transform -1 0 107072 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _220_
timestamp 1666464484
transform 1 0 105168 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _221_
timestamp 1666464484
transform 1 0 104272 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _222_
timestamp 1666464484
transform 1 0 89152 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _223_
timestamp 1666464484
transform -1 0 94976 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _224_
timestamp 1666464484
transform 1 0 94192 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _225_
timestamp 1666464484
transform 1 0 94304 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _226_
timestamp 1666464484
transform -1 0 94976 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _227_
timestamp 1666464484
transform -1 0 95760 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _228_
timestamp 1666464484
transform 1 0 94864 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _229_
timestamp 1666464484
transform -1 0 90832 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _230_
timestamp 1666464484
transform 1 0 85904 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _231_
timestamp 1666464484
transform 1 0 87360 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _232_
timestamp 1666464484
transform 1 0 87360 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _233_
timestamp 1666464484
transform 1 0 88368 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _234_
timestamp 1666464484
transform 1 0 87024 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _235_
timestamp 1666464484
transform 1 0 86128 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _236_
timestamp 1666464484
transform -1 0 75488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _237_
timestamp 1666464484
transform -1 0 78064 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _238_
timestamp 1666464484
transform 1 0 75040 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _239_
timestamp 1666464484
transform 1 0 74816 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _240_
timestamp 1666464484
transform -1 0 78176 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _241_
timestamp 1666464484
transform -1 0 77728 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _242_
timestamp 1666464484
transform 1 0 77168 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _243_
timestamp 1666464484
transform -1 0 67424 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _244_
timestamp 1666464484
transform -1 0 66304 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _245_
timestamp 1666464484
transform -1 0 66976 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _246_
timestamp 1666464484
transform 1 0 66416 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _247_
timestamp 1666464484
transform -1 0 67200 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _248_
timestamp 1666464484
transform -1 0 64848 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _249_
timestamp 1666464484
transform -1 0 64512 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _250_
timestamp 1666464484
transform -1 0 64064 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _251_
timestamp 1666464484
transform -1 0 63952 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _252_
timestamp 1666464484
transform -1 0 65184 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _253_
timestamp 1666464484
transform 1 0 65296 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _254_
timestamp 1666464484
transform -1 0 63840 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _255_
timestamp 1666464484
transform 1 0 60704 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _256_
timestamp 1666464484
transform -1 0 59696 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _257_
timestamp 1666464484
transform -1 0 53312 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _258_
timestamp 1666464484
transform -1 0 54208 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _259_
timestamp 1666464484
transform 1 0 53872 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _260_
timestamp 1666464484
transform 1 0 54208 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _261_
timestamp 1666464484
transform -1 0 54320 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _262_
timestamp 1666464484
transform -1 0 55440 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _263_
timestamp 1666464484
transform 1 0 57456 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _264_
timestamp 1666464484
transform -1 0 60816 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _265_
timestamp 1666464484
transform -1 0 45248 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _266_
timestamp 1666464484
transform 1 0 42784 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _267_
timestamp 1666464484
transform -1 0 42448 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _268_
timestamp 1666464484
transform -1 0 48160 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _269_
timestamp 1666464484
transform 1 0 45360 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _270_
timestamp 1666464484
transform -1 0 44800 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _271_
timestamp 1666464484
transform -1 0 30800 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _272_
timestamp 1666464484
transform 1 0 27776 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _273_
timestamp 1666464484
transform 1 0 28000 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _274_
timestamp 1666464484
transform 1 0 26880 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _275_
timestamp 1666464484
transform 1 0 28784 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _276_
timestamp 1666464484
transform 1 0 26096 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _277_
timestamp 1666464484
transform -1 0 26656 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _278_
timestamp 1666464484
transform -1 0 20384 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _279_
timestamp 1666464484
transform -1 0 20272 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _280_
timestamp 1666464484
transform -1 0 20160 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _281_
timestamp 1666464484
transform -1 0 19264 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _282_
timestamp 1666464484
transform 1 0 17584 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _283_
timestamp 1666464484
transform 1 0 15680 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _284_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 18144 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _285_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 9072 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _286_
timestamp 1666464484
transform 1 0 7280 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _287_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 9184 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _288_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 73696 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _289_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 75712 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _290_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 54208 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _291_
timestamp 1666464484
transform -1 0 52752 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _292_
timestamp 1666464484
transform -1 0 60032 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _293_
timestamp 1666464484
transform -1 0 56896 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _294_
timestamp 1666464484
transform 1 0 26992 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _295_
timestamp 1666464484
transform -1 0 19040 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _296_
timestamp 1666464484
transform -1 0 20832 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _297_
timestamp 1666464484
transform -1 0 28336 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _298_
timestamp 1666464484
transform 1 0 29456 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _299_
timestamp 1666464484
transform 1 0 62272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _300_
timestamp 1666464484
transform -1 0 63840 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _301_
timestamp 1666464484
transform -1 0 47376 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _302_
timestamp 1666464484
transform -1 0 46704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _303_
timestamp 1666464484
transform 1 0 62496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _304_
timestamp 1666464484
transform -1 0 59584 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _305_
timestamp 1666464484
transform -1 0 66864 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _306_
timestamp 1666464484
transform -1 0 62160 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _307_
timestamp 1666464484
transform -1 0 67872 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _308_
timestamp 1666464484
transform 1 0 64400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _309_
timestamp 1666464484
transform -1 0 67984 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _310_
timestamp 1666464484
transform 1 0 85120 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _311_
timestamp 1666464484
transform -1 0 80192 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _312_
timestamp 1666464484
transform 1 0 79744 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _313_
timestamp 1666464484
transform -1 0 89600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _314_
timestamp 1666464484
transform -1 0 90608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _315_
timestamp 1666464484
transform 1 0 89152 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _316_
timestamp 1666464484
transform -1 0 98560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _317_
timestamp 1666464484
transform 1 0 97104 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _318_
timestamp 1666464484
transform 1 0 103488 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _319_
timestamp 1666464484
transform 1 0 104160 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _320_
timestamp 1666464484
transform -1 0 118496 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _321_
timestamp 1666464484
transform -1 0 108416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _322_
timestamp 1666464484
transform -1 0 109536 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _323_
timestamp 1666464484
transform 1 0 115360 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _324_
timestamp 1666464484
transform -1 0 116480 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _325_
timestamp 1666464484
transform 1 0 128912 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _326_
timestamp 1666464484
transform -1 0 131152 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _327_
timestamp 1666464484
transform 1 0 127344 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _328_
timestamp 1666464484
transform -1 0 127568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _329_
timestamp 1666464484
transform -1 0 128352 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _330_
timestamp 1666464484
transform -1 0 129584 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _331_
timestamp 1666464484
transform -1 0 128240 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _332_
timestamp 1666464484
transform -1 0 127120 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _333_
timestamp 1666464484
transform -1 0 126896 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _334_
timestamp 1666464484
transform -1 0 127568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _335_
timestamp 1666464484
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _336_
timestamp 1666464484
transform -1 0 12544 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _337_
timestamp 1666464484
transform 1 0 11984 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _338_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 18368 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _339_
timestamp 1666464484
transform 1 0 17024 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _340_
timestamp 1666464484
transform 1 0 24864 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _341_
timestamp 1666464484
transform 1 0 27664 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _342_
timestamp 1666464484
transform 1 0 43568 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _343_
timestamp 1666464484
transform 1 0 40992 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _344_
timestamp 1666464484
transform 1 0 59808 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _345_
timestamp 1666464484
transform 1 0 55104 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _346_
timestamp 1666464484
transform 1 0 57008 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _347_
timestamp 1666464484
transform -1 0 69104 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _348_
timestamp 1666464484
transform 1 0 62384 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _349_
timestamp 1666464484
transform -1 0 69104 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _350_
timestamp 1666464484
transform -1 0 79520 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _351_
timestamp 1666464484
transform 1 0 77168 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _352_
timestamp 1666464484
transform 1 0 86128 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _353_
timestamp 1666464484
transform 1 0 87024 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _354_
timestamp 1666464484
transform 1 0 95200 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _355_
timestamp 1666464484
transform 1 0 94304 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _356_
timestamp 1666464484
transform -1 0 106848 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _357_
timestamp 1666464484
transform -1 0 106736 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _358_
timestamp 1666464484
transform 1 0 105056 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _359_
timestamp 1666464484
transform 1 0 105056 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _360_
timestamp 1666464484
transform 1 0 113008 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _361_
timestamp 1666464484
transform -1 0 118608 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _362_
timestamp 1666464484
transform 1 0 124880 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _363_
timestamp 1666464484
transform 1 0 128912 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _364_
timestamp 1666464484
transform -1 0 128688 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _365_
timestamp 1666464484
transform 1 0 120624 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _366_
timestamp 1666464484
transform 1 0 122640 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _367_
timestamp 1666464484
transform 1 0 122640 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _368_
timestamp 1666464484
transform 1 0 120624 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _369_
timestamp 1666464484
transform 1 0 122416 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _370_
timestamp 1666464484
transform -1 0 21392 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _371_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 7504 0 1 4704
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _372_
timestamp 1666464484
transform 1 0 9632 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _375_
timestamp 1666464484
transform -1 0 7168 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _376_
timestamp 1666464484
transform 1 0 8512 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _377_
timestamp 1666464484
transform 1 0 12768 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _378_
timestamp 1666464484
transform -1 0 17472 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _379_
timestamp 1666464484
transform -1 0 21504 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _380_
timestamp 1666464484
transform -1 0 24192 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _381_
timestamp 1666464484
transform -1 0 27104 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _382_
timestamp 1666464484
transform -1 0 30128 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _383_
timestamp 1666464484
transform -1 0 32368 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _384_
timestamp 1666464484
transform 1 0 69440 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _385_
timestamp 1666464484
transform 1 0 26096 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _386_
timestamp 1666464484
transform 1 0 34384 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _387_
timestamp 1666464484
transform 1 0 38528 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _388_
timestamp 1666464484
transform 1 0 40320 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _389_
timestamp 1666464484
transform 1 0 52976 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _390_
timestamp 1666464484
transform 1 0 52192 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _391_
timestamp 1666464484
transform 1 0 56336 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _392_
timestamp 1666464484
transform 1 0 86800 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _393_
timestamp 1666464484
transform -1 0 8064 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _394_
timestamp 1666464484
transform 1 0 10080 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _395_
timestamp 1666464484
transform -1 0 14784 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _396_
timestamp 1666464484
transform -1 0 18592 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _397_
timestamp 1666464484
transform -1 0 22400 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _398_
timestamp 1666464484
transform -1 0 25088 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _399_
timestamp 1666464484
transform -1 0 28336 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _400_
timestamp 1666464484
transform 1 0 30352 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _401_
timestamp 1666464484
transform -1 0 34160 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _402_
timestamp 1666464484
transform -1 0 36064 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _403_
timestamp 1666464484
transform -1 0 37968 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _404_
timestamp 1666464484
transform -1 0 39648 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _405_
timestamp 1666464484
transform -1 0 41440 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _406_
timestamp 1666464484
transform -1 0 42896 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _407_
timestamp 1666464484
transform -1 0 58128 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _408_
timestamp 1666464484
transform -1 0 47152 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _409_
timestamp 1666464484
transform 1 0 45920 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _410_
timestamp 1666464484
transform 1 0 48496 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _411_
timestamp 1666464484
transform -1 0 51968 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _412_
timestamp 1666464484
transform -1 0 55104 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _413_
timestamp 1666464484
transform -1 0 84224 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _414_
timestamp 1666464484
transform -1 0 102592 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _415_
timestamp 1666464484
transform -1 0 110880 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _416_
timestamp 1666464484
transform -1 0 113680 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _417_
timestamp 1666464484
transform -1 0 114128 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _418_
timestamp 1666464484
transform -1 0 122080 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _419_
timestamp 1666464484
transform -1 0 126448 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _420_
timestamp 1666464484
transform -1 0 126672 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _421_
timestamp 1666464484
transform -1 0 119280 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _422_
timestamp 1666464484
transform -1 0 85792 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _423_
timestamp 1666464484
transform -1 0 78960 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _424_
timestamp 1666464484
transform -1 0 92624 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _425_
timestamp 1666464484
transform 1 0 73696 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _426_
timestamp 1666464484
transform 1 0 19936 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _427_
timestamp 1666464484
transform 1 0 62048 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _428_
timestamp 1666464484
transform -1 0 90944 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _429_
timestamp 1666464484
transform 1 0 38976 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _430_
timestamp 1666464484
transform 1 0 39424 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _431_
timestamp 1666464484
transform 1 0 47600 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _432_
timestamp 1666464484
transform 1 0 49392 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _433_
timestamp 1666464484
transform 1 0 56672 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _434_
timestamp 1666464484
transform 1 0 79296 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _435_
timestamp 1666464484
transform 1 0 102816 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _436_
timestamp 1666464484
transform 1 0 105056 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _437_
timestamp 1666464484
transform 1 0 106848 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _438_
timestamp 1666464484
transform 1 0 110880 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _439_
timestamp 1666464484
transform 1 0 111776 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _440_
timestamp 1666464484
transform 1 0 113008 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _441_
timestamp 1666464484
transform 1 0 115808 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _442_
timestamp 1666464484
transform 1 0 117600 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _443_
timestamp 1666464484
transform 1 0 119392 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _444_
timestamp 1666464484
transform 1 0 121856 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _445_
timestamp 1666464484
transform 1 0 123200 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _446_
timestamp 1666464484
transform 1 0 107856 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _447_
timestamp 1666464484
transform 1 0 128912 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _448_
timestamp 1666464484
transform 1 0 117712 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _449_
timestamp 1666464484
transform 1 0 132496 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _450_
timestamp 1666464484
transform 1 0 127568 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _451_
timestamp 1666464484
transform 1 0 129136 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _452_
timestamp 1666464484
transform 1 0 129808 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _453_
timestamp 1666464484
transform 1 0 134288 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _454_
timestamp 1666464484
transform 1 0 140784 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _455_
timestamp 1666464484
transform 1 0 142016 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _456_
timestamp 1666464484
transform -1 0 145488 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _457_
timestamp 1666464484
transform 1 0 8288 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _458_
timestamp 1666464484
transform -1 0 13104 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _459_
timestamp 1666464484
transform -1 0 16576 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _460_
timestamp 1666464484
transform 1 0 17808 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _461_
timestamp 1666464484
transform 1 0 22624 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _462_
timestamp 1666464484
transform 1 0 19936 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _463_
timestamp 1666464484
transform 1 0 82992 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _464_
timestamp 1666464484
transform 1 0 59360 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_io_wbs_clk dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 69216 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_io_wbs_clk
timestamp 1666464484
transform 1 0 61264 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_io_wbs_clk
timestamp 1666464484
transform -1 0 64848 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_io_wbs_clk
timestamp 1666464484
transform 1 0 73248 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_io_wbs_clk
timestamp 1666464484
transform 1 0 71120 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1666464484
transform 1 0 8288 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1666464484
transform 1 0 36288 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1666464484
transform 1 0 38080 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1666464484
transform 1 0 39872 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1666464484
transform 1 0 42336 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1666464484
transform 1 0 44128 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1666464484
transform 1 0 45584 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1666464484
transform 1 0 45584 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1666464484
transform 1 0 49504 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1666464484
transform 1 0 50400 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1666464484
transform 1 0 53536 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1666464484
transform 1 0 11536 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1666464484
transform 1 0 54880 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1666464484
transform 1 0 57232 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1666464484
transform 1 0 58464 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1666464484
transform 1 0 58464 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1666464484
transform 1 0 62048 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1666464484
transform 1 0 64064 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1666464484
transform 1 0 64848 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1666464484
transform 1 0 67424 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1666464484
transform 1 0 69216 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1666464484
transform 1 0 70336 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1666464484
transform 1 0 15008 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1666464484
transform 1 0 72800 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1666464484
transform 1 0 73472 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1666464484
transform 1 0 19040 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1666464484
transform 1 0 22624 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1666464484
transform 1 0 25312 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1666464484
transform 1 0 28000 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1666464484
transform 1 0 30688 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1666464484
transform 1 0 32592 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1666464484
transform 1 0 33376 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1666464484
transform -1 0 79744 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1666464484
transform -1 0 108416 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1666464484
transform -1 0 110208 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1666464484
transform -1 0 112000 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1666464484
transform -1 0 114576 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1666464484
transform -1 0 115584 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1666464484
transform -1 0 117376 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1666464484
transform -1 0 120176 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1666464484
transform -1 0 121632 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1666464484
transform -1 0 122976 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1666464484
transform -1 0 125552 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1666464484
transform -1 0 83328 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1666464484
transform -1 0 127344 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1666464484
transform -1 0 129136 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1666464484
transform -1 0 131376 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1666464484
transform -1 0 132272 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1666464484
transform -1 0 133504 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1666464484
transform -1 0 136192 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1666464484
transform -1 0 138096 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1666464484
transform 1 0 137424 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1666464484
transform -1 0 140336 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1666464484
transform -1 0 142464 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1666464484
transform -1 0 86912 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1666464484
transform -1 0 144256 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1666464484
transform -1 0 146384 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1666464484
transform -1 0 92512 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1666464484
transform -1 0 95872 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1666464484
transform -1 0 97664 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1666464484
transform -1 0 100352 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1666464484
transform -1 0 102144 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input63
timestamp 1666464484
transform -1 0 104832 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1666464484
transform -1 0 106624 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input65
timestamp 1666464484
transform 1 0 59136 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input66
timestamp 1666464484
transform -1 0 60816 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input67
timestamp 1666464484
transform 1 0 23296 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input68
timestamp 1666464484
transform -1 0 29792 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input69
timestamp 1666464484
transform 1 0 34048 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input70
timestamp 1666464484
transform -1 0 38640 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input71
timestamp 1666464484
transform -1 0 42560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input72
timestamp 1666464484
transform -1 0 46480 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input73
timestamp 1666464484
transform 1 0 50176 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1666464484
transform -1 0 53536 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1666464484
transform 1 0 6160 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input76
timestamp 1666464484
transform 1 0 15232 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input77
timestamp 1666464484
transform -1 0 59136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input78
timestamp 1666464484
transform -1 0 67760 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input79
timestamp 1666464484
transform 1 0 69328 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input80
timestamp 1666464484
transform -1 0 74704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input81
timestamp 1666464484
transform -1 0 78624 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input82
timestamp 1666464484
transform 1 0 81872 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input83
timestamp 1666464484
transform -1 0 86464 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input84
timestamp 1666464484
transform -1 0 90384 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input85
timestamp 1666464484
transform 1 0 93632 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input86
timestamp 1666464484
transform 1 0 97664 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input87
timestamp 1666464484
transform -1 0 22288 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input88
timestamp 1666464484
transform 1 0 101696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input89
timestamp 1666464484
transform -1 0 106400 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input90
timestamp 1666464484
transform 1 0 109760 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input91
timestamp 1666464484
transform 1 0 113792 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input92
timestamp 1666464484
transform 1 0 117376 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input93
timestamp 1666464484
transform 1 0 121856 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input94
timestamp 1666464484
transform 1 0 125888 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input95
timestamp 1666464484
transform 1 0 129920 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input96
timestamp 1666464484
transform -1 0 134176 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input97
timestamp 1666464484
transform 1 0 137872 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input98
timestamp 1666464484
transform 1 0 25984 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input99
timestamp 1666464484
transform 1 0 141568 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input100
timestamp 1666464484
transform -1 0 146272 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input101
timestamp 1666464484
transform 1 0 31808 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input102
timestamp 1666464484
transform 1 0 36960 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input103
timestamp 1666464484
transform -1 0 41552 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input104
timestamp 1666464484
transform 1 0 44800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input105
timestamp 1666464484
transform 1 0 48832 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input106
timestamp 1666464484
transform -1 0 52192 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input107
timestamp 1666464484
transform 1 0 58352 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input108
timestamp 1666464484
transform 1 0 7056 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input109
timestamp 1666464484
transform 1 0 16240 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input110
timestamp 1666464484
transform -1 0 22624 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input111
timestamp 1666464484
transform 1 0 27328 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input112
timestamp 1666464484
transform 1 0 33040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input113
timestamp 1666464484
transform -1 0 10528 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input114
timestamp 1666464484
transform -1 0 11872 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output115 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 6496 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output116
timestamp 1666464484
transform 1 0 9632 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output117
timestamp 1666464484
transform 1 0 13664 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output118
timestamp 1666464484
transform -1 0 16912 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output119
timestamp 1666464484
transform 1 0 20832 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output120
timestamp 1666464484
transform 1 0 23520 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output121
timestamp 1666464484
transform -1 0 26880 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output122
timestamp 1666464484
transform -1 0 28672 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output123
timestamp 1666464484
transform -1 0 32592 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output124
timestamp 1666464484
transform 1 0 78400 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output125
timestamp 1666464484
transform 1 0 81200 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output126
timestamp 1666464484
transform 1 0 84448 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output127
timestamp 1666464484
transform 1 0 88032 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output128
timestamp 1666464484
transform 1 0 91616 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output129
timestamp 1666464484
transform 1 0 95760 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output130
timestamp 1666464484
transform 1 0 97552 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output131
timestamp 1666464484
transform -1 0 101248 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output132
timestamp 1666464484
transform -1 0 103936 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output133
timestamp 1666464484
transform 1 0 7392 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output134
timestamp 1666464484
transform -1 0 37632 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output135
timestamp 1666464484
transform -1 0 38640 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output136
timestamp 1666464484
transform -1 0 40432 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output137
timestamp 1666464484
transform -1 0 42560 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output138
timestamp 1666464484
transform -1 0 44352 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output139
timestamp 1666464484
transform -1 0 46928 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output140
timestamp 1666464484
transform 1 0 46816 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output141
timestamp 1666464484
transform 1 0 48720 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output142
timestamp 1666464484
transform -1 0 51408 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output143
timestamp 1666464484
transform -1 0 52192 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output144
timestamp 1666464484
transform 1 0 10976 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output145
timestamp 1666464484
transform -1 0 56112 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output146
timestamp 1666464484
transform -1 0 56896 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output147
timestamp 1666464484
transform -1 0 59136 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output148
timestamp 1666464484
transform -1 0 60928 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output149
timestamp 1666464484
transform -1 0 62048 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output150
timestamp 1666464484
transform -1 0 64512 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output151
timestamp 1666464484
transform -1 0 66304 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output152
timestamp 1666464484
transform -1 0 68992 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output153
timestamp 1666464484
transform -1 0 69888 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output154
timestamp 1666464484
transform -1 0 71680 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output155
timestamp 1666464484
transform 1 0 13552 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output156
timestamp 1666464484
transform -1 0 72800 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output157
timestamp 1666464484
transform 1 0 72240 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output158
timestamp 1666464484
transform 1 0 17696 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output159
timestamp 1666464484
transform 1 0 21392 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output160
timestamp 1666464484
transform -1 0 24752 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output161
timestamp 1666464484
transform -1 0 28560 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output162
timestamp 1666464484
transform 1 0 30688 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output163
timestamp 1666464484
transform 1 0 33488 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output164
timestamp 1666464484
transform -1 0 35840 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output165
timestamp 1666464484
transform 1 0 80080 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output166
timestamp 1666464484
transform 1 0 106848 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output167
timestamp 1666464484
transform 1 0 108976 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output168
timestamp 1666464484
transform 1 0 111440 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output169
timestamp 1666464484
transform 1 0 113232 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output170
timestamp 1666464484
transform 1 0 114016 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output171
timestamp 1666464484
transform 1 0 115808 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output172
timestamp 1666464484
transform 1 0 117600 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output173
timestamp 1666464484
transform 1 0 119392 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output174
timestamp 1666464484
transform 1 0 121184 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output175
timestamp 1666464484
transform 1 0 125104 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output176
timestamp 1666464484
transform 1 0 81760 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output177
timestamp 1666464484
transform 1 0 125216 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output178
timestamp 1666464484
transform 1 0 127120 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output179
timestamp 1666464484
transform 1 0 128912 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output180
timestamp 1666464484
transform 1 0 130144 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output181
timestamp 1666464484
transform 1 0 132944 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output182
timestamp 1666464484
transform 1 0 133728 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output183
timestamp 1666464484
transform 1 0 135520 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output184
timestamp 1666464484
transform 1 0 137312 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output185
timestamp 1666464484
transform 1 0 140784 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output186
timestamp 1666464484
transform 1 0 142800 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output187
timestamp 1666464484
transform -1 0 87360 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output188
timestamp 1666464484
transform 1 0 142688 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output189
timestamp 1666464484
transform 1 0 144592 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output190
timestamp 1666464484
transform -1 0 91392 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output191
timestamp 1666464484
transform 1 0 93072 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output192
timestamp 1666464484
transform 1 0 95200 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output193
timestamp 1666464484
transform 1 0 97888 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output194
timestamp 1666464484
transform 1 0 101472 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output195
timestamp 1666464484
transform 1 0 103600 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output196
timestamp 1666464484
transform 1 0 105056 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output197
timestamp 1666464484
transform -1 0 6048 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output198
timestamp 1666464484
transform -1 0 15456 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output199
timestamp 1666464484
transform -1 0 62048 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output200
timestamp 1666464484
transform -1 0 65968 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output201
timestamp 1666464484
transform -1 0 69888 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output202
timestamp 1666464484
transform -1 0 73808 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output203
timestamp 1666464484
transform -1 0 77728 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output204
timestamp 1666464484
transform -1 0 81648 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output205
timestamp 1666464484
transform -1 0 85568 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output206
timestamp 1666464484
transform -1 0 89488 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output207
timestamp 1666464484
transform -1 0 93408 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output208
timestamp 1666464484
transform -1 0 97440 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output209
timestamp 1666464484
transform -1 0 20832 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output210
timestamp 1666464484
transform -1 0 101472 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output211
timestamp 1666464484
transform -1 0 105504 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output212
timestamp 1666464484
transform -1 0 110656 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output213
timestamp 1666464484
transform -1 0 113568 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output214
timestamp 1666464484
transform -1 0 117600 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output215
timestamp 1666464484
transform -1 0 121632 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output216
timestamp 1666464484
transform -1 0 125664 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output217
timestamp 1666464484
transform -1 0 129696 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output218
timestamp 1666464484
transform -1 0 133728 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output219
timestamp 1666464484
transform -1 0 137760 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output220
timestamp 1666464484
transform -1 0 26768 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output221
timestamp 1666464484
transform 1 0 140224 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output222
timestamp 1666464484
transform 1 0 144256 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output223
timestamp 1666464484
transform -1 0 31584 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output224
timestamp 1666464484
transform -1 0 36512 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output225
timestamp 1666464484
transform -1 0 40432 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output226
timestamp 1666464484
transform -1 0 44352 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output227
timestamp 1666464484
transform -1 0 48272 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output228
timestamp 1666464484
transform -1 0 53088 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output229
timestamp 1666464484
transform -1 0 58128 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output230
timestamp 1666464484
transform -1 0 7168 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output231
timestamp 1666464484
transform 1 0 77168 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output232
timestamp 1666464484
transform 1 0 9184 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output233
timestamp 1666464484
transform -1 0 12992 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output234
timestamp 1666464484
transform 1 0 15568 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output235
timestamp 1666464484
transform 1 0 19488 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output236
timestamp 1666464484
transform 1 0 81872 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output237
timestamp 1666464484
transform 1 0 84000 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output238
timestamp 1666464484
transform 1 0 87136 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output239
timestamp 1666464484
transform 1 0 91056 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_memory_240 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 5152 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_memory_241
timestamp 1666464484
transform -1 0 75936 0 -1 34496
box -86 -86 534 870
<< labels >>
flabel metal2 s 6384 39200 6496 40000 0 FreeSans 448 90 0 0 addr_mem0[0]
port 0 nsew signal tristate
flabel metal2 s 9968 39200 10080 40000 0 FreeSans 448 90 0 0 addr_mem0[1]
port 1 nsew signal tristate
flabel metal2 s 13552 39200 13664 40000 0 FreeSans 448 90 0 0 addr_mem0[2]
port 2 nsew signal tristate
flabel metal2 s 17136 39200 17248 40000 0 FreeSans 448 90 0 0 addr_mem0[3]
port 3 nsew signal tristate
flabel metal2 s 20720 39200 20832 40000 0 FreeSans 448 90 0 0 addr_mem0[4]
port 4 nsew signal tristate
flabel metal2 s 23408 39200 23520 40000 0 FreeSans 448 90 0 0 addr_mem0[5]
port 5 nsew signal tristate
flabel metal2 s 26096 39200 26208 40000 0 FreeSans 448 90 0 0 addr_mem0[6]
port 6 nsew signal tristate
flabel metal2 s 28784 39200 28896 40000 0 FreeSans 448 90 0 0 addr_mem0[7]
port 7 nsew signal tristate
flabel metal2 s 31472 39200 31584 40000 0 FreeSans 448 90 0 0 addr_mem0[8]
port 8 nsew signal tristate
flabel metal2 s 77168 39200 77280 40000 0 FreeSans 448 90 0 0 addr_mem1[0]
port 9 nsew signal tristate
flabel metal2 s 80752 39200 80864 40000 0 FreeSans 448 90 0 0 addr_mem1[1]
port 10 nsew signal tristate
flabel metal2 s 84336 39200 84448 40000 0 FreeSans 448 90 0 0 addr_mem1[2]
port 11 nsew signal tristate
flabel metal2 s 87920 39200 88032 40000 0 FreeSans 448 90 0 0 addr_mem1[3]
port 12 nsew signal tristate
flabel metal2 s 91504 39200 91616 40000 0 FreeSans 448 90 0 0 addr_mem1[4]
port 13 nsew signal tristate
flabel metal2 s 94192 39200 94304 40000 0 FreeSans 448 90 0 0 addr_mem1[5]
port 14 nsew signal tristate
flabel metal2 s 96880 39200 96992 40000 0 FreeSans 448 90 0 0 addr_mem1[6]
port 15 nsew signal tristate
flabel metal2 s 99568 39200 99680 40000 0 FreeSans 448 90 0 0 addr_mem1[7]
port 16 nsew signal tristate
flabel metal2 s 102256 39200 102368 40000 0 FreeSans 448 90 0 0 addr_mem1[8]
port 17 nsew signal tristate
flabel metal2 s 4592 39200 4704 40000 0 FreeSans 448 90 0 0 csb_mem0
port 18 nsew signal tristate
flabel metal2 s 75376 39200 75488 40000 0 FreeSans 448 90 0 0 csb_mem1
port 19 nsew signal tristate
flabel metal2 s 7280 39200 7392 40000 0 FreeSans 448 90 0 0 din_mem0[0]
port 20 nsew signal tristate
flabel metal2 s 35952 39200 36064 40000 0 FreeSans 448 90 0 0 din_mem0[10]
port 21 nsew signal tristate
flabel metal2 s 37744 39200 37856 40000 0 FreeSans 448 90 0 0 din_mem0[11]
port 22 nsew signal tristate
flabel metal2 s 39536 39200 39648 40000 0 FreeSans 448 90 0 0 din_mem0[12]
port 23 nsew signal tristate
flabel metal2 s 41328 39200 41440 40000 0 FreeSans 448 90 0 0 din_mem0[13]
port 24 nsew signal tristate
flabel metal2 s 43120 39200 43232 40000 0 FreeSans 448 90 0 0 din_mem0[14]
port 25 nsew signal tristate
flabel metal2 s 44912 39200 45024 40000 0 FreeSans 448 90 0 0 din_mem0[15]
port 26 nsew signal tristate
flabel metal2 s 46704 39200 46816 40000 0 FreeSans 448 90 0 0 din_mem0[16]
port 27 nsew signal tristate
flabel metal2 s 48496 39200 48608 40000 0 FreeSans 448 90 0 0 din_mem0[17]
port 28 nsew signal tristate
flabel metal2 s 50288 39200 50400 40000 0 FreeSans 448 90 0 0 din_mem0[18]
port 29 nsew signal tristate
flabel metal2 s 52080 39200 52192 40000 0 FreeSans 448 90 0 0 din_mem0[19]
port 30 nsew signal tristate
flabel metal2 s 10864 39200 10976 40000 0 FreeSans 448 90 0 0 din_mem0[1]
port 31 nsew signal tristate
flabel metal2 s 53872 39200 53984 40000 0 FreeSans 448 90 0 0 din_mem0[20]
port 32 nsew signal tristate
flabel metal2 s 55664 39200 55776 40000 0 FreeSans 448 90 0 0 din_mem0[21]
port 33 nsew signal tristate
flabel metal2 s 57456 39200 57568 40000 0 FreeSans 448 90 0 0 din_mem0[22]
port 34 nsew signal tristate
flabel metal2 s 59248 39200 59360 40000 0 FreeSans 448 90 0 0 din_mem0[23]
port 35 nsew signal tristate
flabel metal2 s 61040 39200 61152 40000 0 FreeSans 448 90 0 0 din_mem0[24]
port 36 nsew signal tristate
flabel metal2 s 62832 39200 62944 40000 0 FreeSans 448 90 0 0 din_mem0[25]
port 37 nsew signal tristate
flabel metal2 s 64624 39200 64736 40000 0 FreeSans 448 90 0 0 din_mem0[26]
port 38 nsew signal tristate
flabel metal2 s 66416 39200 66528 40000 0 FreeSans 448 90 0 0 din_mem0[27]
port 39 nsew signal tristate
flabel metal2 s 68208 39200 68320 40000 0 FreeSans 448 90 0 0 din_mem0[28]
port 40 nsew signal tristate
flabel metal2 s 70000 39200 70112 40000 0 FreeSans 448 90 0 0 din_mem0[29]
port 41 nsew signal tristate
flabel metal2 s 14448 39200 14560 40000 0 FreeSans 448 90 0 0 din_mem0[2]
port 42 nsew signal tristate
flabel metal2 s 71792 39200 71904 40000 0 FreeSans 448 90 0 0 din_mem0[30]
port 43 nsew signal tristate
flabel metal2 s 73584 39200 73696 40000 0 FreeSans 448 90 0 0 din_mem0[31]
port 44 nsew signal tristate
flabel metal2 s 18032 39200 18144 40000 0 FreeSans 448 90 0 0 din_mem0[3]
port 45 nsew signal tristate
flabel metal2 s 21616 39200 21728 40000 0 FreeSans 448 90 0 0 din_mem0[4]
port 46 nsew signal tristate
flabel metal2 s 24304 39200 24416 40000 0 FreeSans 448 90 0 0 din_mem0[5]
port 47 nsew signal tristate
flabel metal2 s 26992 39200 27104 40000 0 FreeSans 448 90 0 0 din_mem0[6]
port 48 nsew signal tristate
flabel metal2 s 29680 39200 29792 40000 0 FreeSans 448 90 0 0 din_mem0[7]
port 49 nsew signal tristate
flabel metal2 s 32368 39200 32480 40000 0 FreeSans 448 90 0 0 din_mem0[8]
port 50 nsew signal tristate
flabel metal2 s 34160 39200 34272 40000 0 FreeSans 448 90 0 0 din_mem0[9]
port 51 nsew signal tristate
flabel metal2 s 78064 39200 78176 40000 0 FreeSans 448 90 0 0 din_mem1[0]
port 52 nsew signal tristate
flabel metal2 s 106736 39200 106848 40000 0 FreeSans 448 90 0 0 din_mem1[10]
port 53 nsew signal tristate
flabel metal2 s 108528 39200 108640 40000 0 FreeSans 448 90 0 0 din_mem1[11]
port 54 nsew signal tristate
flabel metal2 s 110320 39200 110432 40000 0 FreeSans 448 90 0 0 din_mem1[12]
port 55 nsew signal tristate
flabel metal2 s 112112 39200 112224 40000 0 FreeSans 448 90 0 0 din_mem1[13]
port 56 nsew signal tristate
flabel metal2 s 113904 39200 114016 40000 0 FreeSans 448 90 0 0 din_mem1[14]
port 57 nsew signal tristate
flabel metal2 s 115696 39200 115808 40000 0 FreeSans 448 90 0 0 din_mem1[15]
port 58 nsew signal tristate
flabel metal2 s 117488 39200 117600 40000 0 FreeSans 448 90 0 0 din_mem1[16]
port 59 nsew signal tristate
flabel metal2 s 119280 39200 119392 40000 0 FreeSans 448 90 0 0 din_mem1[17]
port 60 nsew signal tristate
flabel metal2 s 121072 39200 121184 40000 0 FreeSans 448 90 0 0 din_mem1[18]
port 61 nsew signal tristate
flabel metal2 s 122864 39200 122976 40000 0 FreeSans 448 90 0 0 din_mem1[19]
port 62 nsew signal tristate
flabel metal2 s 81648 39200 81760 40000 0 FreeSans 448 90 0 0 din_mem1[1]
port 63 nsew signal tristate
flabel metal2 s 124656 39200 124768 40000 0 FreeSans 448 90 0 0 din_mem1[20]
port 64 nsew signal tristate
flabel metal2 s 126448 39200 126560 40000 0 FreeSans 448 90 0 0 din_mem1[21]
port 65 nsew signal tristate
flabel metal2 s 128240 39200 128352 40000 0 FreeSans 448 90 0 0 din_mem1[22]
port 66 nsew signal tristate
flabel metal2 s 130032 39200 130144 40000 0 FreeSans 448 90 0 0 din_mem1[23]
port 67 nsew signal tristate
flabel metal2 s 131824 39200 131936 40000 0 FreeSans 448 90 0 0 din_mem1[24]
port 68 nsew signal tristate
flabel metal2 s 133616 39200 133728 40000 0 FreeSans 448 90 0 0 din_mem1[25]
port 69 nsew signal tristate
flabel metal2 s 135408 39200 135520 40000 0 FreeSans 448 90 0 0 din_mem1[26]
port 70 nsew signal tristate
flabel metal2 s 137200 39200 137312 40000 0 FreeSans 448 90 0 0 din_mem1[27]
port 71 nsew signal tristate
flabel metal2 s 138992 39200 139104 40000 0 FreeSans 448 90 0 0 din_mem1[28]
port 72 nsew signal tristate
flabel metal2 s 140784 39200 140896 40000 0 FreeSans 448 90 0 0 din_mem1[29]
port 73 nsew signal tristate
flabel metal2 s 85232 39200 85344 40000 0 FreeSans 448 90 0 0 din_mem1[2]
port 74 nsew signal tristate
flabel metal2 s 142576 39200 142688 40000 0 FreeSans 448 90 0 0 din_mem1[30]
port 75 nsew signal tristate
flabel metal2 s 144368 39200 144480 40000 0 FreeSans 448 90 0 0 din_mem1[31]
port 76 nsew signal tristate
flabel metal2 s 88816 39200 88928 40000 0 FreeSans 448 90 0 0 din_mem1[3]
port 77 nsew signal tristate
flabel metal2 s 92400 39200 92512 40000 0 FreeSans 448 90 0 0 din_mem1[4]
port 78 nsew signal tristate
flabel metal2 s 95088 39200 95200 40000 0 FreeSans 448 90 0 0 din_mem1[5]
port 79 nsew signal tristate
flabel metal2 s 97776 39200 97888 40000 0 FreeSans 448 90 0 0 din_mem1[6]
port 80 nsew signal tristate
flabel metal2 s 100464 39200 100576 40000 0 FreeSans 448 90 0 0 din_mem1[7]
port 81 nsew signal tristate
flabel metal2 s 103152 39200 103264 40000 0 FreeSans 448 90 0 0 din_mem1[8]
port 82 nsew signal tristate
flabel metal2 s 104944 39200 105056 40000 0 FreeSans 448 90 0 0 din_mem1[9]
port 83 nsew signal tristate
flabel metal2 s 8176 39200 8288 40000 0 FreeSans 448 90 0 0 dout_mem0[0]
port 84 nsew signal input
flabel metal2 s 36848 39200 36960 40000 0 FreeSans 448 90 0 0 dout_mem0[10]
port 85 nsew signal input
flabel metal2 s 38640 39200 38752 40000 0 FreeSans 448 90 0 0 dout_mem0[11]
port 86 nsew signal input
flabel metal2 s 40432 39200 40544 40000 0 FreeSans 448 90 0 0 dout_mem0[12]
port 87 nsew signal input
flabel metal2 s 42224 39200 42336 40000 0 FreeSans 448 90 0 0 dout_mem0[13]
port 88 nsew signal input
flabel metal2 s 44016 39200 44128 40000 0 FreeSans 448 90 0 0 dout_mem0[14]
port 89 nsew signal input
flabel metal2 s 45808 39200 45920 40000 0 FreeSans 448 90 0 0 dout_mem0[15]
port 90 nsew signal input
flabel metal2 s 47600 39200 47712 40000 0 FreeSans 448 90 0 0 dout_mem0[16]
port 91 nsew signal input
flabel metal2 s 49392 39200 49504 40000 0 FreeSans 448 90 0 0 dout_mem0[17]
port 92 nsew signal input
flabel metal2 s 51184 39200 51296 40000 0 FreeSans 448 90 0 0 dout_mem0[18]
port 93 nsew signal input
flabel metal2 s 52976 39200 53088 40000 0 FreeSans 448 90 0 0 dout_mem0[19]
port 94 nsew signal input
flabel metal2 s 11760 39200 11872 40000 0 FreeSans 448 90 0 0 dout_mem0[1]
port 95 nsew signal input
flabel metal2 s 54768 39200 54880 40000 0 FreeSans 448 90 0 0 dout_mem0[20]
port 96 nsew signal input
flabel metal2 s 56560 39200 56672 40000 0 FreeSans 448 90 0 0 dout_mem0[21]
port 97 nsew signal input
flabel metal2 s 58352 39200 58464 40000 0 FreeSans 448 90 0 0 dout_mem0[22]
port 98 nsew signal input
flabel metal2 s 60144 39200 60256 40000 0 FreeSans 448 90 0 0 dout_mem0[23]
port 99 nsew signal input
flabel metal2 s 61936 39200 62048 40000 0 FreeSans 448 90 0 0 dout_mem0[24]
port 100 nsew signal input
flabel metal2 s 63728 39200 63840 40000 0 FreeSans 448 90 0 0 dout_mem0[25]
port 101 nsew signal input
flabel metal2 s 65520 39200 65632 40000 0 FreeSans 448 90 0 0 dout_mem0[26]
port 102 nsew signal input
flabel metal2 s 67312 39200 67424 40000 0 FreeSans 448 90 0 0 dout_mem0[27]
port 103 nsew signal input
flabel metal2 s 69104 39200 69216 40000 0 FreeSans 448 90 0 0 dout_mem0[28]
port 104 nsew signal input
flabel metal2 s 70896 39200 71008 40000 0 FreeSans 448 90 0 0 dout_mem0[29]
port 105 nsew signal input
flabel metal2 s 15344 39200 15456 40000 0 FreeSans 448 90 0 0 dout_mem0[2]
port 106 nsew signal input
flabel metal2 s 72688 39200 72800 40000 0 FreeSans 448 90 0 0 dout_mem0[30]
port 107 nsew signal input
flabel metal2 s 74480 39200 74592 40000 0 FreeSans 448 90 0 0 dout_mem0[31]
port 108 nsew signal input
flabel metal2 s 18928 39200 19040 40000 0 FreeSans 448 90 0 0 dout_mem0[3]
port 109 nsew signal input
flabel metal2 s 22512 39200 22624 40000 0 FreeSans 448 90 0 0 dout_mem0[4]
port 110 nsew signal input
flabel metal2 s 25200 39200 25312 40000 0 FreeSans 448 90 0 0 dout_mem0[5]
port 111 nsew signal input
flabel metal2 s 27888 39200 28000 40000 0 FreeSans 448 90 0 0 dout_mem0[6]
port 112 nsew signal input
flabel metal2 s 30576 39200 30688 40000 0 FreeSans 448 90 0 0 dout_mem0[7]
port 113 nsew signal input
flabel metal2 s 33264 39200 33376 40000 0 FreeSans 448 90 0 0 dout_mem0[8]
port 114 nsew signal input
flabel metal2 s 35056 39200 35168 40000 0 FreeSans 448 90 0 0 dout_mem0[9]
port 115 nsew signal input
flabel metal2 s 78960 39200 79072 40000 0 FreeSans 448 90 0 0 dout_mem1[0]
port 116 nsew signal input
flabel metal2 s 107632 39200 107744 40000 0 FreeSans 448 90 0 0 dout_mem1[10]
port 117 nsew signal input
flabel metal2 s 109424 39200 109536 40000 0 FreeSans 448 90 0 0 dout_mem1[11]
port 118 nsew signal input
flabel metal2 s 111216 39200 111328 40000 0 FreeSans 448 90 0 0 dout_mem1[12]
port 119 nsew signal input
flabel metal2 s 113008 39200 113120 40000 0 FreeSans 448 90 0 0 dout_mem1[13]
port 120 nsew signal input
flabel metal2 s 114800 39200 114912 40000 0 FreeSans 448 90 0 0 dout_mem1[14]
port 121 nsew signal input
flabel metal2 s 116592 39200 116704 40000 0 FreeSans 448 90 0 0 dout_mem1[15]
port 122 nsew signal input
flabel metal2 s 118384 39200 118496 40000 0 FreeSans 448 90 0 0 dout_mem1[16]
port 123 nsew signal input
flabel metal2 s 120176 39200 120288 40000 0 FreeSans 448 90 0 0 dout_mem1[17]
port 124 nsew signal input
flabel metal2 s 121968 39200 122080 40000 0 FreeSans 448 90 0 0 dout_mem1[18]
port 125 nsew signal input
flabel metal2 s 123760 39200 123872 40000 0 FreeSans 448 90 0 0 dout_mem1[19]
port 126 nsew signal input
flabel metal2 s 82544 39200 82656 40000 0 FreeSans 448 90 0 0 dout_mem1[1]
port 127 nsew signal input
flabel metal2 s 125552 39200 125664 40000 0 FreeSans 448 90 0 0 dout_mem1[20]
port 128 nsew signal input
flabel metal2 s 127344 39200 127456 40000 0 FreeSans 448 90 0 0 dout_mem1[21]
port 129 nsew signal input
flabel metal2 s 129136 39200 129248 40000 0 FreeSans 448 90 0 0 dout_mem1[22]
port 130 nsew signal input
flabel metal2 s 130928 39200 131040 40000 0 FreeSans 448 90 0 0 dout_mem1[23]
port 131 nsew signal input
flabel metal2 s 132720 39200 132832 40000 0 FreeSans 448 90 0 0 dout_mem1[24]
port 132 nsew signal input
flabel metal2 s 134512 39200 134624 40000 0 FreeSans 448 90 0 0 dout_mem1[25]
port 133 nsew signal input
flabel metal2 s 136304 39200 136416 40000 0 FreeSans 448 90 0 0 dout_mem1[26]
port 134 nsew signal input
flabel metal2 s 138096 39200 138208 40000 0 FreeSans 448 90 0 0 dout_mem1[27]
port 135 nsew signal input
flabel metal2 s 139888 39200 140000 40000 0 FreeSans 448 90 0 0 dout_mem1[28]
port 136 nsew signal input
flabel metal2 s 141680 39200 141792 40000 0 FreeSans 448 90 0 0 dout_mem1[29]
port 137 nsew signal input
flabel metal2 s 86128 39200 86240 40000 0 FreeSans 448 90 0 0 dout_mem1[2]
port 138 nsew signal input
flabel metal2 s 143472 39200 143584 40000 0 FreeSans 448 90 0 0 dout_mem1[30]
port 139 nsew signal input
flabel metal2 s 145264 39200 145376 40000 0 FreeSans 448 90 0 0 dout_mem1[31]
port 140 nsew signal input
flabel metal2 s 89712 39200 89824 40000 0 FreeSans 448 90 0 0 dout_mem1[3]
port 141 nsew signal input
flabel metal2 s 93296 39200 93408 40000 0 FreeSans 448 90 0 0 dout_mem1[4]
port 142 nsew signal input
flabel metal2 s 95984 39200 96096 40000 0 FreeSans 448 90 0 0 dout_mem1[5]
port 143 nsew signal input
flabel metal2 s 98672 39200 98784 40000 0 FreeSans 448 90 0 0 dout_mem1[6]
port 144 nsew signal input
flabel metal2 s 101360 39200 101472 40000 0 FreeSans 448 90 0 0 dout_mem1[7]
port 145 nsew signal input
flabel metal2 s 104048 39200 104160 40000 0 FreeSans 448 90 0 0 dout_mem1[8]
port 146 nsew signal input
flabel metal2 s 105840 39200 105952 40000 0 FreeSans 448 90 0 0 dout_mem1[9]
port 147 nsew signal input
flabel metal2 s 4368 0 4480 800 0 FreeSans 448 90 0 0 io_wbs_ack
port 148 nsew signal tristate
flabel metal2 s 12432 0 12544 800 0 FreeSans 448 90 0 0 io_wbs_adr[0]
port 149 nsew signal input
flabel metal2 s 58128 0 58240 800 0 FreeSans 448 90 0 0 io_wbs_adr[10]
port 150 nsew signal input
flabel metal2 s 62160 0 62272 800 0 FreeSans 448 90 0 0 io_wbs_adr[11]
port 151 nsew signal input
flabel metal2 s 66192 0 66304 800 0 FreeSans 448 90 0 0 io_wbs_adr[12]
port 152 nsew signal input
flabel metal2 s 70224 0 70336 800 0 FreeSans 448 90 0 0 io_wbs_adr[13]
port 153 nsew signal input
flabel metal2 s 74256 0 74368 800 0 FreeSans 448 90 0 0 io_wbs_adr[14]
port 154 nsew signal input
flabel metal2 s 78288 0 78400 800 0 FreeSans 448 90 0 0 io_wbs_adr[15]
port 155 nsew signal input
flabel metal2 s 82320 0 82432 800 0 FreeSans 448 90 0 0 io_wbs_adr[16]
port 156 nsew signal input
flabel metal2 s 86352 0 86464 800 0 FreeSans 448 90 0 0 io_wbs_adr[17]
port 157 nsew signal input
flabel metal2 s 90384 0 90496 800 0 FreeSans 448 90 0 0 io_wbs_adr[18]
port 158 nsew signal input
flabel metal2 s 94416 0 94528 800 0 FreeSans 448 90 0 0 io_wbs_adr[19]
port 159 nsew signal input
flabel metal2 s 17808 0 17920 800 0 FreeSans 448 90 0 0 io_wbs_adr[1]
port 160 nsew signal input
flabel metal2 s 98448 0 98560 800 0 FreeSans 448 90 0 0 io_wbs_adr[20]
port 161 nsew signal input
flabel metal2 s 102480 0 102592 800 0 FreeSans 448 90 0 0 io_wbs_adr[21]
port 162 nsew signal input
flabel metal2 s 106512 0 106624 800 0 FreeSans 448 90 0 0 io_wbs_adr[22]
port 163 nsew signal input
flabel metal2 s 110544 0 110656 800 0 FreeSans 448 90 0 0 io_wbs_adr[23]
port 164 nsew signal input
flabel metal2 s 114576 0 114688 800 0 FreeSans 448 90 0 0 io_wbs_adr[24]
port 165 nsew signal input
flabel metal2 s 118608 0 118720 800 0 FreeSans 448 90 0 0 io_wbs_adr[25]
port 166 nsew signal input
flabel metal2 s 122640 0 122752 800 0 FreeSans 448 90 0 0 io_wbs_adr[26]
port 167 nsew signal input
flabel metal2 s 126672 0 126784 800 0 FreeSans 448 90 0 0 io_wbs_adr[27]
port 168 nsew signal input
flabel metal2 s 130704 0 130816 800 0 FreeSans 448 90 0 0 io_wbs_adr[28]
port 169 nsew signal input
flabel metal2 s 134736 0 134848 800 0 FreeSans 448 90 0 0 io_wbs_adr[29]
port 170 nsew signal input
flabel metal2 s 23184 0 23296 800 0 FreeSans 448 90 0 0 io_wbs_adr[2]
port 171 nsew signal input
flabel metal2 s 138768 0 138880 800 0 FreeSans 448 90 0 0 io_wbs_adr[30]
port 172 nsew signal input
flabel metal2 s 142800 0 142912 800 0 FreeSans 448 90 0 0 io_wbs_adr[31]
port 173 nsew signal input
flabel metal2 s 28560 0 28672 800 0 FreeSans 448 90 0 0 io_wbs_adr[3]
port 174 nsew signal input
flabel metal2 s 33936 0 34048 800 0 FreeSans 448 90 0 0 io_wbs_adr[4]
port 175 nsew signal input
flabel metal2 s 37968 0 38080 800 0 FreeSans 448 90 0 0 io_wbs_adr[5]
port 176 nsew signal input
flabel metal2 s 42000 0 42112 800 0 FreeSans 448 90 0 0 io_wbs_adr[6]
port 177 nsew signal input
flabel metal2 s 46032 0 46144 800 0 FreeSans 448 90 0 0 io_wbs_adr[7]
port 178 nsew signal input
flabel metal2 s 50064 0 50176 800 0 FreeSans 448 90 0 0 io_wbs_adr[8]
port 179 nsew signal input
flabel metal2 s 54096 0 54208 800 0 FreeSans 448 90 0 0 io_wbs_adr[9]
port 180 nsew signal input
flabel metal2 s 5712 0 5824 800 0 FreeSans 448 90 0 0 io_wbs_clk
port 181 nsew signal input
flabel metal2 s 7056 0 7168 800 0 FreeSans 448 90 0 0 io_wbs_cyc
port 182 nsew signal input
flabel metal2 s 13776 0 13888 800 0 FreeSans 448 90 0 0 io_wbs_datrd[0]
port 183 nsew signal tristate
flabel metal2 s 59472 0 59584 800 0 FreeSans 448 90 0 0 io_wbs_datrd[10]
port 184 nsew signal tristate
flabel metal2 s 63504 0 63616 800 0 FreeSans 448 90 0 0 io_wbs_datrd[11]
port 185 nsew signal tristate
flabel metal2 s 67536 0 67648 800 0 FreeSans 448 90 0 0 io_wbs_datrd[12]
port 186 nsew signal tristate
flabel metal2 s 71568 0 71680 800 0 FreeSans 448 90 0 0 io_wbs_datrd[13]
port 187 nsew signal tristate
flabel metal2 s 75600 0 75712 800 0 FreeSans 448 90 0 0 io_wbs_datrd[14]
port 188 nsew signal tristate
flabel metal2 s 79632 0 79744 800 0 FreeSans 448 90 0 0 io_wbs_datrd[15]
port 189 nsew signal tristate
flabel metal2 s 83664 0 83776 800 0 FreeSans 448 90 0 0 io_wbs_datrd[16]
port 190 nsew signal tristate
flabel metal2 s 87696 0 87808 800 0 FreeSans 448 90 0 0 io_wbs_datrd[17]
port 191 nsew signal tristate
flabel metal2 s 91728 0 91840 800 0 FreeSans 448 90 0 0 io_wbs_datrd[18]
port 192 nsew signal tristate
flabel metal2 s 95760 0 95872 800 0 FreeSans 448 90 0 0 io_wbs_datrd[19]
port 193 nsew signal tristate
flabel metal2 s 19152 0 19264 800 0 FreeSans 448 90 0 0 io_wbs_datrd[1]
port 194 nsew signal tristate
flabel metal2 s 99792 0 99904 800 0 FreeSans 448 90 0 0 io_wbs_datrd[20]
port 195 nsew signal tristate
flabel metal2 s 103824 0 103936 800 0 FreeSans 448 90 0 0 io_wbs_datrd[21]
port 196 nsew signal tristate
flabel metal2 s 107856 0 107968 800 0 FreeSans 448 90 0 0 io_wbs_datrd[22]
port 197 nsew signal tristate
flabel metal2 s 111888 0 112000 800 0 FreeSans 448 90 0 0 io_wbs_datrd[23]
port 198 nsew signal tristate
flabel metal2 s 115920 0 116032 800 0 FreeSans 448 90 0 0 io_wbs_datrd[24]
port 199 nsew signal tristate
flabel metal2 s 119952 0 120064 800 0 FreeSans 448 90 0 0 io_wbs_datrd[25]
port 200 nsew signal tristate
flabel metal2 s 123984 0 124096 800 0 FreeSans 448 90 0 0 io_wbs_datrd[26]
port 201 nsew signal tristate
flabel metal2 s 128016 0 128128 800 0 FreeSans 448 90 0 0 io_wbs_datrd[27]
port 202 nsew signal tristate
flabel metal2 s 132048 0 132160 800 0 FreeSans 448 90 0 0 io_wbs_datrd[28]
port 203 nsew signal tristate
flabel metal2 s 136080 0 136192 800 0 FreeSans 448 90 0 0 io_wbs_datrd[29]
port 204 nsew signal tristate
flabel metal2 s 24528 0 24640 800 0 FreeSans 448 90 0 0 io_wbs_datrd[2]
port 205 nsew signal tristate
flabel metal2 s 140112 0 140224 800 0 FreeSans 448 90 0 0 io_wbs_datrd[30]
port 206 nsew signal tristate
flabel metal2 s 144144 0 144256 800 0 FreeSans 448 90 0 0 io_wbs_datrd[31]
port 207 nsew signal tristate
flabel metal2 s 29904 0 30016 800 0 FreeSans 448 90 0 0 io_wbs_datrd[3]
port 208 nsew signal tristate
flabel metal2 s 35280 0 35392 800 0 FreeSans 448 90 0 0 io_wbs_datrd[4]
port 209 nsew signal tristate
flabel metal2 s 39312 0 39424 800 0 FreeSans 448 90 0 0 io_wbs_datrd[5]
port 210 nsew signal tristate
flabel metal2 s 43344 0 43456 800 0 FreeSans 448 90 0 0 io_wbs_datrd[6]
port 211 nsew signal tristate
flabel metal2 s 47376 0 47488 800 0 FreeSans 448 90 0 0 io_wbs_datrd[7]
port 212 nsew signal tristate
flabel metal2 s 51408 0 51520 800 0 FreeSans 448 90 0 0 io_wbs_datrd[8]
port 213 nsew signal tristate
flabel metal2 s 55440 0 55552 800 0 FreeSans 448 90 0 0 io_wbs_datrd[9]
port 214 nsew signal tristate
flabel metal2 s 15120 0 15232 800 0 FreeSans 448 90 0 0 io_wbs_datwr[0]
port 215 nsew signal input
flabel metal2 s 60816 0 60928 800 0 FreeSans 448 90 0 0 io_wbs_datwr[10]
port 216 nsew signal input
flabel metal2 s 64848 0 64960 800 0 FreeSans 448 90 0 0 io_wbs_datwr[11]
port 217 nsew signal input
flabel metal2 s 68880 0 68992 800 0 FreeSans 448 90 0 0 io_wbs_datwr[12]
port 218 nsew signal input
flabel metal2 s 72912 0 73024 800 0 FreeSans 448 90 0 0 io_wbs_datwr[13]
port 219 nsew signal input
flabel metal2 s 76944 0 77056 800 0 FreeSans 448 90 0 0 io_wbs_datwr[14]
port 220 nsew signal input
flabel metal2 s 80976 0 81088 800 0 FreeSans 448 90 0 0 io_wbs_datwr[15]
port 221 nsew signal input
flabel metal2 s 85008 0 85120 800 0 FreeSans 448 90 0 0 io_wbs_datwr[16]
port 222 nsew signal input
flabel metal2 s 89040 0 89152 800 0 FreeSans 448 90 0 0 io_wbs_datwr[17]
port 223 nsew signal input
flabel metal2 s 93072 0 93184 800 0 FreeSans 448 90 0 0 io_wbs_datwr[18]
port 224 nsew signal input
flabel metal2 s 97104 0 97216 800 0 FreeSans 448 90 0 0 io_wbs_datwr[19]
port 225 nsew signal input
flabel metal2 s 20496 0 20608 800 0 FreeSans 448 90 0 0 io_wbs_datwr[1]
port 226 nsew signal input
flabel metal2 s 101136 0 101248 800 0 FreeSans 448 90 0 0 io_wbs_datwr[20]
port 227 nsew signal input
flabel metal2 s 105168 0 105280 800 0 FreeSans 448 90 0 0 io_wbs_datwr[21]
port 228 nsew signal input
flabel metal2 s 109200 0 109312 800 0 FreeSans 448 90 0 0 io_wbs_datwr[22]
port 229 nsew signal input
flabel metal2 s 113232 0 113344 800 0 FreeSans 448 90 0 0 io_wbs_datwr[23]
port 230 nsew signal input
flabel metal2 s 117264 0 117376 800 0 FreeSans 448 90 0 0 io_wbs_datwr[24]
port 231 nsew signal input
flabel metal2 s 121296 0 121408 800 0 FreeSans 448 90 0 0 io_wbs_datwr[25]
port 232 nsew signal input
flabel metal2 s 125328 0 125440 800 0 FreeSans 448 90 0 0 io_wbs_datwr[26]
port 233 nsew signal input
flabel metal2 s 129360 0 129472 800 0 FreeSans 448 90 0 0 io_wbs_datwr[27]
port 234 nsew signal input
flabel metal2 s 133392 0 133504 800 0 FreeSans 448 90 0 0 io_wbs_datwr[28]
port 235 nsew signal input
flabel metal2 s 137424 0 137536 800 0 FreeSans 448 90 0 0 io_wbs_datwr[29]
port 236 nsew signal input
flabel metal2 s 25872 0 25984 800 0 FreeSans 448 90 0 0 io_wbs_datwr[2]
port 237 nsew signal input
flabel metal2 s 141456 0 141568 800 0 FreeSans 448 90 0 0 io_wbs_datwr[30]
port 238 nsew signal input
flabel metal2 s 145488 0 145600 800 0 FreeSans 448 90 0 0 io_wbs_datwr[31]
port 239 nsew signal input
flabel metal2 s 31248 0 31360 800 0 FreeSans 448 90 0 0 io_wbs_datwr[3]
port 240 nsew signal input
flabel metal2 s 36624 0 36736 800 0 FreeSans 448 90 0 0 io_wbs_datwr[4]
port 241 nsew signal input
flabel metal2 s 40656 0 40768 800 0 FreeSans 448 90 0 0 io_wbs_datwr[5]
port 242 nsew signal input
flabel metal2 s 44688 0 44800 800 0 FreeSans 448 90 0 0 io_wbs_datwr[6]
port 243 nsew signal input
flabel metal2 s 48720 0 48832 800 0 FreeSans 448 90 0 0 io_wbs_datwr[7]
port 244 nsew signal input
flabel metal2 s 52752 0 52864 800 0 FreeSans 448 90 0 0 io_wbs_datwr[8]
port 245 nsew signal input
flabel metal2 s 56784 0 56896 800 0 FreeSans 448 90 0 0 io_wbs_datwr[9]
port 246 nsew signal input
flabel metal2 s 8400 0 8512 800 0 FreeSans 448 90 0 0 io_wbs_rst
port 247 nsew signal input
flabel metal2 s 16464 0 16576 800 0 FreeSans 448 90 0 0 io_wbs_sel[0]
port 248 nsew signal input
flabel metal2 s 21840 0 21952 800 0 FreeSans 448 90 0 0 io_wbs_sel[1]
port 249 nsew signal input
flabel metal2 s 27216 0 27328 800 0 FreeSans 448 90 0 0 io_wbs_sel[2]
port 250 nsew signal input
flabel metal2 s 32592 0 32704 800 0 FreeSans 448 90 0 0 io_wbs_sel[3]
port 251 nsew signal input
flabel metal2 s 9744 0 9856 800 0 FreeSans 448 90 0 0 io_wbs_stb
port 252 nsew signal input
flabel metal2 s 11088 0 11200 800 0 FreeSans 448 90 0 0 io_wbs_we
port 253 nsew signal input
flabel metal4 s 19594 3076 19914 36908 0 FreeSans 1280 90 0 0 vdd
port 254 nsew power bidirectional
flabel metal4 s 56414 3076 56734 36908 0 FreeSans 1280 90 0 0 vdd
port 254 nsew power bidirectional
flabel metal4 s 93234 3076 93554 36908 0 FreeSans 1280 90 0 0 vdd
port 254 nsew power bidirectional
flabel metal4 s 130054 3076 130374 36908 0 FreeSans 1280 90 0 0 vdd
port 254 nsew power bidirectional
flabel metal4 s 38004 3076 38324 36908 0 FreeSans 1280 90 0 0 vss
port 255 nsew ground bidirectional
flabel metal4 s 74824 3076 75144 36908 0 FreeSans 1280 90 0 0 vss
port 255 nsew ground bidirectional
flabel metal4 s 111644 3076 111964 36908 0 FreeSans 1280 90 0 0 vss
port 255 nsew ground bidirectional
flabel metal4 s 148464 3076 148784 36908 0 FreeSans 1280 90 0 0 vss
port 255 nsew ground bidirectional
flabel metal2 s 5488 39200 5600 40000 0 FreeSans 448 90 0 0 web_mem0
port 256 nsew signal tristate
flabel metal2 s 76272 39200 76384 40000 0 FreeSans 448 90 0 0 web_mem1
port 257 nsew signal tristate
flabel metal2 s 9072 39200 9184 40000 0 FreeSans 448 90 0 0 wmask_mem0[0]
port 258 nsew signal tristate
flabel metal2 s 12656 39200 12768 40000 0 FreeSans 448 90 0 0 wmask_mem0[1]
port 259 nsew signal tristate
flabel metal2 s 16240 39200 16352 40000 0 FreeSans 448 90 0 0 wmask_mem0[2]
port 260 nsew signal tristate
flabel metal2 s 19824 39200 19936 40000 0 FreeSans 448 90 0 0 wmask_mem0[3]
port 261 nsew signal tristate
flabel metal2 s 79856 39200 79968 40000 0 FreeSans 448 90 0 0 wmask_mem1[0]
port 262 nsew signal tristate
flabel metal2 s 83440 39200 83552 40000 0 FreeSans 448 90 0 0 wmask_mem1[1]
port 263 nsew signal tristate
flabel metal2 s 87024 39200 87136 40000 0 FreeSans 448 90 0 0 wmask_mem1[2]
port 264 nsew signal tristate
flabel metal2 s 90608 39200 90720 40000 0 FreeSans 448 90 0 0 wmask_mem1[3]
port 265 nsew signal tristate
rlabel metal1 74984 36848 74984 36848 0 vdd
rlabel via1 75064 36064 75064 36064 0 vss
rlabel metal2 10248 4368 10248 4368 0 _000_
rlabel metal2 8232 4816 8232 4816 0 _001_
rlabel metal2 18760 4144 18760 4144 0 _002_
rlabel metal2 20104 5264 20104 5264 0 _003_
rlabel metal2 28056 4704 28056 4704 0 _004_
rlabel metal3 30184 5320 30184 5320 0 _005_
rlabel metal2 47096 5712 47096 5712 0 _006_
rlabel metal2 44184 5040 44184 5040 0 _007_
rlabel metal2 62776 7056 62776 7056 0 _008_
rlabel metal2 58296 5040 58296 5040 0 _009_
rlabel metal3 60928 6552 60928 6552 0 _010_
rlabel metal2 67592 6272 67592 6272 0 _011_
rlabel metal2 65072 6552 65072 6552 0 _012_
rlabel metal2 67704 5376 67704 5376 0 _013_
rlabel metal3 78232 5992 78232 5992 0 _014_
rlabel metal2 80080 4536 80080 4536 0 _015_
rlabel metal2 89320 5264 89320 5264 0 _016_
rlabel metal2 90272 5320 90272 5320 0 _017_
rlabel metal2 98280 6272 98280 6272 0 _018_
rlabel metal2 97384 5264 97384 5264 0 _019_
rlabel metal2 103768 5264 103768 5264 0 _020_
rlabel metal3 104104 6104 104104 6104 0 _021_
rlabel metal2 108136 4704 108136 4704 0 _022_
rlabel metal3 108752 6104 108752 6104 0 _023_
rlabel metal2 115640 5656 115640 5656 0 _024_
rlabel metal2 115640 4816 115640 4816 0 _025_
rlabel metal2 130872 5656 130872 5656 0 _026_
rlabel metal2 131992 5152 131992 5152 0 _027_
rlabel metal2 125720 4312 125720 4312 0 _028_
rlabel metal2 123816 4704 123816 4704 0 _029_
rlabel metal2 125832 5096 125832 5096 0 _030_
rlabel metal3 126336 7672 126336 7672 0 _031_
rlabel metal2 126616 6272 126616 6272 0 _032_
rlabel metal3 126448 6104 126448 6104 0 _033_
rlabel metal3 17584 4200 17584 4200 0 _034_
rlabel metal3 11368 3752 11368 3752 0 _035_
rlabel metal2 12600 4704 12600 4704 0 _036_
rlabel metal3 16912 6104 16912 6104 0 _037_
rlabel metal2 17752 5544 17752 5544 0 _038_
rlabel metal2 25592 5768 25592 5768 0 _039_
rlabel metal3 27832 6440 27832 6440 0 _040_
rlabel metal2 44296 6720 44296 6720 0 _041_
rlabel metal2 41720 5768 41720 5768 0 _042_
rlabel metal2 57960 4984 57960 4984 0 _043_
rlabel metal2 54712 5096 54712 5096 0 _044_
rlabel metal2 57736 7112 57736 7112 0 _045_
rlabel metal2 68376 7112 68376 7112 0 _046_
rlabel metal3 63560 6104 63560 6104 0 _047_
rlabel metal2 66920 5376 66920 5376 0 _048_
rlabel metal2 77672 6160 77672 6160 0 _049_
rlabel metal2 75320 5544 75320 5544 0 _050_
rlabel metal2 86688 6440 86688 6440 0 _051_
rlabel metal2 87808 6104 87808 6104 0 _052_
rlabel metal2 95368 6272 95368 6272 0 _053_
rlabel metal2 94864 6440 94864 6440 0 _054_
rlabel metal2 104776 7280 104776 7280 0 _055_
rlabel metal2 104440 7112 104440 7112 0 _056_
rlabel metal3 106512 4312 106512 4312 0 _057_
rlabel metal2 105784 6160 105784 6160 0 _058_
rlabel metal2 113736 6160 113736 6160 0 _059_
rlabel metal2 117992 4424 117992 4424 0 _060_
rlabel metal2 125496 5712 125496 5712 0 _061_
rlabel metal3 128520 4424 128520 4424 0 _062_
rlabel metal3 131936 4984 131936 4984 0 _063_
rlabel metal2 123872 3640 123872 3640 0 _064_
rlabel metal2 123368 5712 123368 5712 0 _065_
rlabel metal2 123368 7672 123368 7672 0 _066_
rlabel metal2 121352 7112 121352 7112 0 _067_
rlabel metal2 123144 6944 123144 6944 0 _068_
rlabel metal2 53816 35336 53816 35336 0 _069_
rlabel metal2 75488 36232 75488 36232 0 _070_
rlabel metal3 26040 5936 26040 5936 0 _071_
rlabel metal2 138096 5992 138096 5992 0 _072_
rlabel metal3 124544 8232 124544 8232 0 _073_
rlabel metal3 121352 8344 121352 8344 0 _074_
rlabel metal2 122136 7672 122136 7672 0 _075_
rlabel metal2 20328 32760 20328 32760 0 _076_
rlabel metal2 139216 35000 139216 35000 0 _077_
rlabel metal3 140560 5208 140560 5208 0 _078_
rlabel metal2 137368 6776 137368 6776 0 _079_
rlabel metal3 139440 7672 139440 7672 0 _080_
rlabel metal3 136920 6552 136920 6552 0 _081_
rlabel metal2 140840 6720 140840 6720 0 _082_
rlabel metal2 141288 6216 141288 6216 0 _083_
rlabel metal2 139720 5768 139720 5768 0 _084_
rlabel metal2 138824 4928 138824 4928 0 _085_
rlabel metal2 136472 4984 136472 4984 0 _086_
rlabel metal2 131432 36120 131432 36120 0 _087_
rlabel metal3 133336 6104 133336 6104 0 _088_
rlabel metal2 127288 4760 127288 4760 0 _089_
rlabel metal3 132664 5320 132664 5320 0 _090_
rlabel metal2 130312 5040 130312 5040 0 _091_
rlabel metal3 119056 5320 119056 5320 0 _092_
rlabel metal2 115416 6552 115416 6552 0 _093_
rlabel metal2 119336 4648 119336 4648 0 _094_
rlabel metal3 117096 7448 117096 7448 0 _095_
rlabel metal2 115080 6944 115080 6944 0 _096_
rlabel metal2 74424 34552 74424 34552 0 _097_
rlabel metal2 88536 33768 88536 33768 0 _098_
rlabel metal3 111888 4536 111888 4536 0 _099_
rlabel metal3 107800 3752 107800 3752 0 _100_
rlabel metal3 110488 5208 110488 5208 0 _101_
rlabel metal2 107576 5096 107576 5096 0 _102_
rlabel metal3 106456 8232 106456 8232 0 _103_
rlabel metal2 54040 6384 54040 6384 0 _104_
rlabel metal2 95592 8176 95592 8176 0 _105_
rlabel metal3 104776 7560 104776 7560 0 _106_
rlabel metal3 106680 7448 106680 7448 0 _107_
rlabel metal2 105392 7336 105392 7336 0 _108_
rlabel metal2 93576 35728 93576 35728 0 _109_
rlabel metal3 95480 8232 95480 8232 0 _110_
rlabel metal2 94584 7336 94584 7336 0 _111_
rlabel metal3 95592 7672 95592 7672 0 _112_
rlabel metal2 95200 5880 95200 5880 0 _113_
rlabel metal3 88704 8232 88704 8232 0 _114_
rlabel metal2 78008 7224 78008 7224 0 _115_
rlabel metal2 87528 7000 87528 7000 0 _116_
rlabel metal2 87696 7448 87696 7448 0 _117_
rlabel metal2 86576 6664 86576 6664 0 _118_
rlabel metal3 71624 34888 71624 34888 0 _119_
rlabel metal2 78568 6720 78568 6720 0 _120_
rlabel metal2 75152 5880 75152 5880 0 _121_
rlabel metal3 77784 7448 77784 7448 0 _122_
rlabel metal2 77448 6944 77448 6944 0 _123_
rlabel metal2 66416 7448 66416 7448 0 _124_
rlabel metal3 62776 7448 62776 7448 0 _125_
rlabel metal2 66696 6944 66696 6944 0 _126_
rlabel metal2 64232 7504 64232 7504 0 _127_
rlabel metal2 64344 6608 64344 6608 0 _128_
rlabel metal3 53648 33320 53648 33320 0 _129_
rlabel metal3 65800 8232 65800 8232 0 _130_
rlabel metal2 64904 8736 64904 8736 0 _131_
rlabel metal2 61656 7728 61656 7728 0 _132_
rlabel metal3 60256 7448 60256 7448 0 _133_
rlabel metal2 54488 4760 54488 4760 0 _134_
rlabel metal3 44688 7336 44688 7336 0 _135_
rlabel metal2 54152 4760 54152 4760 0 _136_
rlabel metal2 54824 4928 54824 4928 0 _137_
rlabel metal2 57624 4032 57624 4032 0 _138_
rlabel metal2 29848 36008 29848 36008 0 _139_
rlabel metal2 44912 6664 44912 6664 0 _140_
rlabel metal2 42672 6552 42672 6552 0 _141_
rlabel metal2 47936 6664 47936 6664 0 _142_
rlabel metal3 45136 6664 45136 6664 0 _143_
rlabel metal3 29512 7448 29512 7448 0 _144_
rlabel metal2 26936 7448 26936 7448 0 _145_
rlabel metal2 27160 6944 27160 6944 0 _146_
rlabel metal2 28056 7728 28056 7728 0 _147_
rlabel metal2 26376 6944 26376 6944 0 _148_
rlabel metal2 20552 6776 20552 6776 0 _149_
rlabel metal2 19992 6216 19992 6216 0 _150_
rlabel metal3 19880 5880 19880 5880 0 _151_
rlabel metal3 16912 5880 16912 5880 0 _152_
rlabel metal2 8568 3696 8568 3696 0 _153_
rlabel metal2 8120 3808 8120 3808 0 _154_
rlabel metal3 74984 34328 74984 34328 0 _155_
rlabel metal2 52584 34608 52584 34608 0 _156_
rlabel metal2 119336 3808 119336 3808 0 _157_
rlabel metal2 27160 4480 27160 4480 0 _158_
rlabel metal2 20664 5264 20664 5264 0 _159_
rlabel metal2 70280 4368 70280 4368 0 _160_
rlabel metal2 47712 5208 47712 5208 0 _161_
rlabel metal3 67928 6664 67928 6664 0 _162_
rlabel metal3 90804 4872 90804 4872 0 _163_
rlabel metal2 96600 5712 96600 5712 0 _164_
rlabel metal2 114968 5600 114968 5600 0 _165_
rlabel metal3 128464 6104 128464 6104 0 _166_
rlabel metal2 128072 5656 128072 5656 0 _167_
rlabel metal3 7000 35784 7000 35784 0 addr_mem0[0]
rlabel metal2 10472 36736 10472 36736 0 addr_mem0[1]
rlabel metal2 14448 35560 14448 35560 0 addr_mem0[2]
rlabel metal3 16632 36568 16632 36568 0 addr_mem0[3]
rlabel metal2 21560 35560 21560 35560 0 addr_mem0[4]
rlabel metal3 23912 35560 23912 35560 0 addr_mem0[5]
rlabel metal2 26096 36568 26096 36568 0 addr_mem0[6]
rlabel metal3 28336 36568 28336 36568 0 addr_mem0[7]
rlabel metal2 31528 37898 31528 37898 0 addr_mem0[8]
rlabel metal2 77224 37394 77224 37394 0 addr_mem1[0]
rlabel metal3 81424 35560 81424 35560 0 addr_mem1[1]
rlabel metal2 85176 35560 85176 35560 0 addr_mem1[2]
rlabel metal2 88872 35056 88872 35056 0 addr_mem1[3]
rlabel metal2 92680 34272 92680 34272 0 addr_mem1[4]
rlabel metal3 95424 36568 95424 36568 0 addr_mem1[5]
rlabel metal2 96936 37898 96936 37898 0 addr_mem1[6]
rlabel metal2 100072 37184 100072 37184 0 addr_mem1[7]
rlabel metal3 102592 35784 102592 35784 0 addr_mem1[8]
rlabel metal3 73752 4312 73752 4312 0 clknet_0_io_wbs_clk
rlabel metal2 28728 4816 28728 4816 0 clknet_2_0__leaf_io_wbs_clk
rlabel metal2 27720 6272 27720 6272 0 clknet_2_1__leaf_io_wbs_clk
rlabel metal2 78456 4760 78456 4760 0 clknet_2_2__leaf_io_wbs_clk
rlabel metal2 77448 5152 77448 5152 0 clknet_2_3__leaf_io_wbs_clk
rlabel metal2 8120 36568 8120 36568 0 din_mem0[0]
rlabel metal2 36568 36232 36568 36232 0 din_mem0[10]
rlabel metal2 37800 37898 37800 37898 0 din_mem0[11]
rlabel metal2 39592 37898 39592 37898 0 din_mem0[12]
rlabel metal2 41384 37898 41384 37898 0 din_mem0[13]
rlabel metal2 43176 37898 43176 37898 0 din_mem0[14]
rlabel metal2 45752 35056 45752 35056 0 din_mem0[15]
rlabel metal2 47656 36120 47656 36120 0 din_mem0[16]
rlabel metal3 49056 36568 49056 36568 0 din_mem0[17]
rlabel metal2 50344 37506 50344 37506 0 din_mem0[18]
rlabel metal3 51744 36568 51744 36568 0 din_mem0[19]
rlabel metal2 11816 35784 11816 35784 0 din_mem0[1]
rlabel metal2 54936 37072 54936 37072 0 din_mem0[20]
rlabel metal2 55832 36568 55832 36568 0 din_mem0[21]
rlabel metal2 57960 37184 57960 37184 0 din_mem0[22]
rlabel metal2 59752 36568 59752 36568 0 din_mem0[23]
rlabel metal2 61096 37898 61096 37898 0 din_mem0[24]
rlabel metal3 63168 35000 63168 35000 0 din_mem0[25]
rlabel metal2 65128 36232 65128 36232 0 din_mem0[26]
rlabel metal2 67928 36176 67928 36176 0 din_mem0[27]
rlabel metal2 68936 36736 68936 36736 0 din_mem0[28]
rlabel metal2 70616 36736 70616 36736 0 din_mem0[29]
rlabel metal2 14504 37898 14504 37898 0 din_mem0[2]
rlabel metal2 71848 37394 71848 37394 0 din_mem0[30]
rlabel metal2 73416 37184 73416 37184 0 din_mem0[31]
rlabel metal2 18480 35000 18480 35000 0 din_mem0[3]
rlabel metal3 21952 36568 21952 36568 0 din_mem0[4]
rlabel metal2 23912 37184 23912 37184 0 din_mem0[5]
rlabel metal2 27216 35560 27216 35560 0 din_mem0[6]
rlabel metal3 30632 35560 30632 35560 0 din_mem0[7]
rlabel metal3 33488 35784 33488 35784 0 din_mem0[8]
rlabel metal2 34664 37184 34664 37184 0 din_mem0[9]
rlabel metal2 78120 38010 78120 38010 0 din_mem1[0]
rlabel metal2 107688 35112 107688 35112 0 din_mem1[10]
rlabel metal2 109816 35056 109816 35056 0 din_mem1[11]
rlabel metal2 112280 36624 112280 36624 0 din_mem1[12]
rlabel metal3 113120 36568 113120 36568 0 din_mem1[13]
rlabel metal2 113960 37394 113960 37394 0 din_mem1[14]
rlabel metal3 116200 36568 116200 36568 0 din_mem1[15]
rlabel metal3 117992 35560 117992 35560 0 din_mem1[16]
rlabel metal2 120232 37184 120232 37184 0 din_mem1[17]
rlabel metal2 122024 37184 122024 37184 0 din_mem1[18]
rlabel metal3 124488 36568 124488 36568 0 din_mem1[19]
rlabel metal3 82152 35000 82152 35000 0 din_mem1[1]
rlabel metal3 125496 35784 125496 35784 0 din_mem1[20]
rlabel metal3 127232 36568 127232 36568 0 din_mem1[21]
rlabel metal3 129024 36568 129024 36568 0 din_mem1[22]
rlabel metal2 131096 34944 131096 34944 0 din_mem1[23]
rlabel metal2 133784 36736 133784 36736 0 din_mem1[24]
rlabel metal3 134232 35784 134232 35784 0 din_mem1[25]
rlabel metal2 136360 35056 136360 35056 0 din_mem1[26]
rlabel metal2 138152 35112 138152 35112 0 din_mem1[27]
rlabel metal2 141624 36624 141624 36624 0 din_mem1[28]
rlabel metal3 142240 36568 142240 36568 0 din_mem1[29]
rlabel metal2 86184 36680 86184 36680 0 din_mem1[2]
rlabel metal2 143752 35840 143752 35840 0 din_mem1[30]
rlabel metal3 144928 36568 144928 36568 0 din_mem1[31]
rlabel metal3 89488 35000 89488 35000 0 din_mem1[3]
rlabel metal3 93240 35000 93240 35000 0 din_mem1[4]
rlabel metal2 96040 35056 96040 35056 0 din_mem1[5]
rlabel metal2 98616 35560 98616 35560 0 din_mem1[6]
rlabel metal3 101472 36568 101472 36568 0 din_mem1[7]
rlabel metal3 103824 36568 103824 36568 0 din_mem1[8]
rlabel metal3 105448 35000 105448 35000 0 din_mem1[9]
rlabel metal2 8344 35560 8344 35560 0 dout_mem0[0]
rlabel metal2 36736 34888 36736 34888 0 dout_mem0[10]
rlabel metal2 38472 34888 38472 34888 0 dout_mem0[11]
rlabel metal2 40152 35056 40152 35056 0 dout_mem0[12]
rlabel metal2 42168 35000 42168 35000 0 dout_mem0[13]
rlabel metal2 43960 35000 43960 35000 0 dout_mem0[14]
rlabel metal2 45864 36666 45864 36666 0 dout_mem0[15]
rlabel metal2 45752 36680 45752 36680 0 dout_mem0[16]
rlabel metal2 49672 35000 49672 35000 0 dout_mem0[17]
rlabel metal2 50680 35448 50680 35448 0 dout_mem0[18]
rlabel metal2 53648 35784 53648 35784 0 dout_mem0[19]
rlabel metal2 11872 34888 11872 34888 0 dout_mem0[1]
rlabel metal2 55048 36456 55048 36456 0 dout_mem0[20]
rlabel metal2 56056 36008 56056 36008 0 dout_mem0[21]
rlabel metal2 58520 34888 58520 34888 0 dout_mem0[22]
rlabel metal3 59416 35784 59416 35784 0 dout_mem0[23]
rlabel metal3 61880 33432 61880 33432 0 dout_mem0[24]
rlabel metal2 64232 35896 64232 35896 0 dout_mem0[25]
rlabel metal3 65296 36456 65296 36456 0 dout_mem0[26]
rlabel metal2 67368 37058 67368 37058 0 dout_mem0[27]
rlabel metal2 69272 34888 69272 34888 0 dout_mem0[28]
rlabel metal3 70728 35784 70728 35784 0 dout_mem0[29]
rlabel metal2 15344 34888 15344 34888 0 dout_mem0[2]
rlabel metal2 72856 34888 72856 34888 0 dout_mem0[30]
rlabel metal2 73752 35896 73752 35896 0 dout_mem0[31]
rlabel metal2 19208 35392 19208 35392 0 dout_mem0[3]
rlabel metal2 22680 34888 22680 34888 0 dout_mem0[4]
rlabel metal2 25368 34888 25368 34888 0 dout_mem0[5]
rlabel metal2 27720 35056 27720 35056 0 dout_mem0[6]
rlabel metal2 30408 35056 30408 35056 0 dout_mem0[7]
rlabel metal3 33096 34888 33096 34888 0 dout_mem0[8]
rlabel metal3 35616 36568 35616 36568 0 dout_mem0[9]
rlabel metal2 79016 36778 79016 36778 0 dout_mem1[0]
rlabel metal2 108136 34776 108136 34776 0 dout_mem1[10]
rlabel metal2 109256 34384 109256 34384 0 dout_mem1[11]
rlabel metal2 111720 34944 111720 34944 0 dout_mem1[12]
rlabel metal3 115136 34776 115136 34776 0 dout_mem1[13]
rlabel metal2 115304 35504 115304 35504 0 dout_mem1[14]
rlabel metal2 117096 36232 117096 36232 0 dout_mem1[15]
rlabel metal2 119896 35000 119896 35000 0 dout_mem1[16]
rlabel metal2 120904 37408 120904 37408 0 dout_mem1[17]
rlabel metal3 122416 34888 122416 34888 0 dout_mem1[18]
rlabel metal3 124656 34888 124656 34888 0 dout_mem1[19]
rlabel metal2 82376 35056 82376 35056 0 dout_mem1[1]
rlabel metal3 126336 34888 126336 34888 0 dout_mem1[20]
rlabel metal3 128184 34888 128184 34888 0 dout_mem1[21]
rlabel metal3 130200 34216 130200 34216 0 dout_mem1[22]
rlabel metal2 132104 34720 132104 34720 0 dout_mem1[23]
rlabel metal3 133000 34888 133000 34888 0 dout_mem1[24]
rlabel metal3 135240 35672 135240 35672 0 dout_mem1[25]
rlabel metal2 136360 37842 136360 37842 0 dout_mem1[26]
rlabel metal2 138152 37450 138152 37450 0 dout_mem1[27]
rlabel metal2 140056 35784 140056 35784 0 dout_mem1[28]
rlabel metal2 141512 35056 141512 35056 0 dout_mem1[29]
rlabel metal2 86632 36344 86632 36344 0 dout_mem1[2]
rlabel metal3 143752 34888 143752 34888 0 dout_mem1[30]
rlabel metal2 146216 35840 146216 35840 0 dout_mem1[31]
rlabel metal2 91840 33432 91840 33432 0 dout_mem1[3]
rlabel metal2 95592 35448 95592 35448 0 dout_mem1[4]
rlabel metal2 97384 34944 97384 34944 0 dout_mem1[5]
rlabel metal2 100072 35448 100072 35448 0 dout_mem1[6]
rlabel metal2 101304 35896 101304 35896 0 dout_mem1[7]
rlabel metal2 103992 35000 103992 35000 0 dout_mem1[8]
rlabel metal2 105672 34776 105672 34776 0 dout_mem1[9]
rlabel metal2 4424 2478 4424 2478 0 io_wbs_ack
rlabel metal3 58744 4984 58744 4984 0 io_wbs_adr[10]
rlabel metal3 61432 4984 61432 4984 0 io_wbs_adr[11]
rlabel metal2 23128 3416 23128 3416 0 io_wbs_adr[2]
rlabel metal2 28616 2086 28616 2086 0 io_wbs_adr[3]
rlabel metal2 34104 3416 34104 3416 0 io_wbs_adr[4]
rlabel metal2 38472 2968 38472 2968 0 io_wbs_adr[5]
rlabel metal2 42280 3024 42280 3024 0 io_wbs_adr[6]
rlabel metal2 46144 3528 46144 3528 0 io_wbs_adr[7]
rlabel metal2 50008 3416 50008 3416 0 io_wbs_adr[8]
rlabel metal3 53760 3416 53760 3416 0 io_wbs_adr[9]
rlabel metal2 6440 112 6440 112 0 io_wbs_clk
rlabel metal3 6720 3416 6720 3416 0 io_wbs_cyc
rlabel metal2 13832 2086 13832 2086 0 io_wbs_datrd[0]
rlabel metal2 59528 1246 59528 1246 0 io_wbs_datrd[10]
rlabel metal2 63560 2086 63560 2086 0 io_wbs_datrd[11]
rlabel metal2 67592 1246 67592 1246 0 io_wbs_datrd[12]
rlabel metal2 71624 2086 71624 2086 0 io_wbs_datrd[13]
rlabel metal2 75656 2086 75656 2086 0 io_wbs_datrd[14]
rlabel metal2 79688 2086 79688 2086 0 io_wbs_datrd[15]
rlabel metal2 83720 2086 83720 2086 0 io_wbs_datrd[16]
rlabel metal2 87752 2086 87752 2086 0 io_wbs_datrd[17]
rlabel metal2 91784 2086 91784 2086 0 io_wbs_datrd[18]
rlabel metal2 95816 2086 95816 2086 0 io_wbs_datrd[19]
rlabel metal2 19208 2198 19208 2198 0 io_wbs_datrd[1]
rlabel metal2 99848 2086 99848 2086 0 io_wbs_datrd[20]
rlabel metal2 103880 2086 103880 2086 0 io_wbs_datrd[21]
rlabel metal2 107912 2478 107912 2478 0 io_wbs_datrd[22]
rlabel metal2 111944 854 111944 854 0 io_wbs_datrd[23]
rlabel metal2 115976 2086 115976 2086 0 io_wbs_datrd[24]
rlabel metal2 120008 2086 120008 2086 0 io_wbs_datrd[25]
rlabel metal2 124040 2086 124040 2086 0 io_wbs_datrd[26]
rlabel metal2 128072 2086 128072 2086 0 io_wbs_datrd[27]
rlabel metal2 132104 2086 132104 2086 0 io_wbs_datrd[28]
rlabel metal2 136136 2086 136136 2086 0 io_wbs_datrd[29]
rlabel metal2 24584 2086 24584 2086 0 io_wbs_datrd[2]
rlabel metal2 140168 2086 140168 2086 0 io_wbs_datrd[30]
rlabel metal2 144200 2086 144200 2086 0 io_wbs_datrd[31]
rlabel metal2 29960 2086 29960 2086 0 io_wbs_datrd[3]
rlabel metal2 35336 2198 35336 2198 0 io_wbs_datrd[4]
rlabel metal2 39368 2086 39368 2086 0 io_wbs_datrd[5]
rlabel metal2 43400 2198 43400 2198 0 io_wbs_datrd[6]
rlabel metal2 47432 2198 47432 2198 0 io_wbs_datrd[7]
rlabel metal2 51464 2478 51464 2478 0 io_wbs_datrd[8]
rlabel metal2 55496 2086 55496 2086 0 io_wbs_datrd[9]
rlabel metal2 15288 4312 15288 4312 0 io_wbs_datwr[0]
rlabel metal2 58968 3584 58968 3584 0 io_wbs_datwr[10]
rlabel metal3 69104 3528 69104 3528 0 io_wbs_datwr[11]
rlabel metal2 69496 2520 69496 2520 0 io_wbs_datwr[12]
rlabel metal3 73752 3416 73752 3416 0 io_wbs_datwr[13]
rlabel metal3 77728 3416 77728 3416 0 io_wbs_datwr[14]
rlabel metal3 81536 3416 81536 3416 0 io_wbs_datwr[15]
rlabel metal3 85680 3416 85680 3416 0 io_wbs_datwr[16]
rlabel metal3 89712 3416 89712 3416 0 io_wbs_datwr[17]
rlabel metal3 93464 3416 93464 3416 0 io_wbs_datwr[18]
rlabel metal3 97496 3416 97496 3416 0 io_wbs_datwr[19]
rlabel metal3 21336 4312 21336 4312 0 io_wbs_datwr[1]
rlabel metal3 101528 3416 101528 3416 0 io_wbs_datwr[20]
rlabel metal3 105728 3416 105728 3416 0 io_wbs_datwr[21]
rlabel metal2 109928 2072 109928 2072 0 io_wbs_datwr[22]
rlabel metal2 113960 2072 113960 2072 0 io_wbs_datwr[23]
rlabel metal2 117544 4984 117544 4984 0 io_wbs_datwr[24]
rlabel metal3 121688 3416 121688 3416 0 io_wbs_datwr[25]
rlabel metal2 125384 2142 125384 2142 0 io_wbs_datwr[26]
rlabel metal2 130088 2072 130088 2072 0 io_wbs_datwr[27]
rlabel metal2 133896 3584 133896 3584 0 io_wbs_datwr[28]
rlabel metal2 138040 3976 138040 3976 0 io_wbs_datwr[29]
rlabel metal2 26040 4312 26040 4312 0 io_wbs_datwr[2]
rlabel metal2 141400 4200 141400 4200 0 io_wbs_datwr[30]
rlabel metal2 145432 4200 145432 4200 0 io_wbs_datwr[31]
rlabel metal3 31584 3416 31584 3416 0 io_wbs_datwr[3]
rlabel metal2 36904 3416 36904 3416 0 io_wbs_datwr[4]
rlabel metal3 40992 3528 40992 3528 0 io_wbs_datwr[5]
rlabel metal2 44856 3416 44856 3416 0 io_wbs_datwr[6]
rlabel metal2 48888 3416 48888 3416 0 io_wbs_datwr[7]
rlabel metal3 52416 3528 52416 3528 0 io_wbs_datwr[8]
rlabel metal2 56840 5152 56840 5152 0 io_wbs_datwr[9]
rlabel metal3 6608 3528 6608 3528 0 io_wbs_rst
rlabel metal2 16520 2142 16520 2142 0 io_wbs_sel[0]
rlabel metal2 22344 3136 22344 3136 0 io_wbs_sel[1]
rlabel metal2 27384 3416 27384 3416 0 io_wbs_sel[2]
rlabel metal3 32928 3416 32928 3416 0 io_wbs_sel[3]
rlabel metal3 10080 3416 10080 3416 0 io_wbs_stb
rlabel metal2 11032 3416 11032 3416 0 io_wbs_we
rlabel metal2 17528 33824 17528 33824 0 net1
rlabel metal2 51016 34496 51016 34496 0 net10
rlabel metal2 93464 34440 93464 34440 0 net100
rlabel metal2 25088 4872 25088 4872 0 net101
rlabel metal2 22456 33880 22456 33880 0 net102
rlabel metal2 24920 34440 24920 34440 0 net103
rlabel metal3 46200 26936 46200 26936 0 net104
rlabel metal2 31416 35056 31416 35056 0 net105
rlabel metal2 51688 5320 51688 5320 0 net106
rlabel metal2 58856 4592 58856 4592 0 net107
rlabel metal2 7560 3136 7560 3136 0 net108
rlabel metal2 23352 34384 23352 34384 0 net109
rlabel metal2 54208 35784 54208 35784 0 net11
rlabel metal2 22064 3304 22064 3304 0 net110
rlabel metal2 26936 27944 26936 27944 0 net111
rlabel metal2 18200 20636 18200 20636 0 net112
rlabel metal2 8344 3976 8344 3976 0 net113
rlabel metal3 10136 3304 10136 3304 0 net114
rlabel metal2 6664 35224 6664 35224 0 net115
rlabel metal2 9016 36176 9016 36176 0 net116
rlabel metal3 13552 35784 13552 35784 0 net117
rlabel metal2 16968 35616 16968 35616 0 net118
rlabel metal2 21000 35000 21000 35000 0 net119
rlabel metal2 12040 35224 12040 35224 0 net12
rlabel metal2 23688 35224 23688 35224 0 net120
rlabel metal2 26544 34776 26544 34776 0 net121
rlabel metal2 29624 35616 29624 35616 0 net122
rlabel metal2 31864 35616 31864 35616 0 net123
rlabel metal2 69944 35728 69944 35728 0 net124
rlabel metal2 26600 36736 26600 36736 0 net125
rlabel metal3 59640 29176 59640 29176 0 net126
rlabel metal2 39032 37128 39032 37128 0 net127
rlabel metal2 44520 30380 44520 30380 0 net128
rlabel metal2 96376 35392 96376 35392 0 net129
rlabel metal2 55384 32312 55384 32312 0 net13
rlabel metal2 52472 30772 52472 30772 0 net130
rlabel metal2 92344 37128 92344 37128 0 net131
rlabel metal2 87304 35952 87304 35952 0 net132
rlabel metal2 7616 34776 7616 34776 0 net133
rlabel metal2 37464 35000 37464 35000 0 net134
rlabel metal2 39144 35616 39144 35616 0 net135
rlabel metal2 40936 35616 40936 35616 0 net136
rlabel metal2 42392 36176 42392 36176 0 net137
rlabel metal2 43400 35728 43400 35728 0 net138
rlabel metal2 46648 34608 46648 34608 0 net139
rlabel metal2 57736 33096 57736 33096 0 net14
rlabel metal3 46704 35784 46704 35784 0 net140
rlabel metal2 49000 35616 49000 35616 0 net141
rlabel metal2 51464 35224 51464 35224 0 net142
rlabel metal2 54600 36008 54600 36008 0 net143
rlabel metal2 10584 35728 10584 35728 0 net144
rlabel metal2 55832 33768 55832 33768 0 net145
rlabel metal2 57512 35000 57512 35000 0 net146
rlabel metal3 60144 36456 60144 36456 0 net147
rlabel metal2 60760 36680 60760 36680 0 net148
rlabel metal3 62328 32760 62328 32760 0 net149
rlabel metal2 58968 32368 58968 32368 0 net15
rlabel metal2 64344 36176 64344 36176 0 net150
rlabel metal2 66304 34888 66304 34888 0 net151
rlabel metal2 68936 35672 68936 35672 0 net152
rlabel metal2 69720 37128 69720 37128 0 net153
rlabel metal2 71624 35112 71624 35112 0 net154
rlabel metal2 14280 35616 14280 35616 0 net155
rlabel metal2 72632 35952 72632 35952 0 net156
rlabel metal2 72744 33712 72744 33712 0 net157
rlabel metal2 18088 34608 18088 34608 0 net158
rlabel metal2 21896 35056 21896 35056 0 net159
rlabel metal2 58968 37240 58968 37240 0 net16
rlabel metal2 24528 34776 24528 34776 0 net160
rlabel metal2 27832 35224 27832 35224 0 net161
rlabel metal2 30856 35224 30856 35224 0 net162
rlabel metal2 33656 35224 33656 35224 0 net163
rlabel metal2 35560 35616 35560 35616 0 net164
rlabel metal2 74200 34440 74200 34440 0 net165
rlabel metal3 105168 34776 105168 34776 0 net166
rlabel metal2 109256 35168 109256 35168 0 net167
rlabel metal2 111496 35840 111496 35840 0 net168
rlabel metal3 112392 35896 112392 35896 0 net169
rlabel metal2 62664 32536 62664 32536 0 net17
rlabel metal2 114296 35728 114296 35728 0 net170
rlabel metal2 115976 35560 115976 35560 0 net171
rlabel metal3 117040 35784 117040 35784 0 net172
rlabel metal2 118104 36400 118104 36400 0 net173
rlabel metal2 121352 36176 121352 36176 0 net174
rlabel metal3 123816 35896 123816 35896 0 net175
rlabel metal3 22736 34216 22736 34216 0 net176
rlabel metal2 123704 35224 123704 35224 0 net177
rlabel metal2 108360 35560 108360 35560 0 net178
rlabel metal2 129472 34328 129472 34328 0 net179
rlabel metal2 64624 35896 64624 35896 0 net18
rlabel metal2 118216 33824 118216 33824 0 net180
rlabel metal2 133056 35896 133056 35896 0 net181
rlabel metal2 133896 35392 133896 35392 0 net182
rlabel metal2 135800 34048 135800 34048 0 net183
rlabel metal2 137480 34608 137480 34608 0 net184
rlabel metal2 141064 35504 141064 35504 0 net185
rlabel metal2 141288 35056 141288 35056 0 net186
rlabel metal2 62608 34664 62608 34664 0 net187
rlabel metal2 142520 35224 142520 35224 0 net188
rlabel metal2 144984 36176 144984 36176 0 net189
rlabel metal3 65520 36344 65520 36344 0 net19
rlabel metal2 91000 35168 91000 35168 0 net190
rlabel metal2 93688 34888 93688 34888 0 net191
rlabel metal2 95256 34888 95256 34888 0 net192
rlabel metal3 49224 34664 49224 34664 0 net193
rlabel metal2 49896 31360 49896 31360 0 net194
rlabel metal2 57176 37184 57176 37184 0 net195
rlabel metal2 79800 33656 79800 33656 0 net196
rlabel metal2 6216 4816 6216 4816 0 net197
rlabel metal3 16688 6440 16688 6440 0 net198
rlabel metal2 63560 7392 63560 7392 0 net199
rlabel metal4 52136 33208 52136 33208 0 net2
rlabel metal2 67984 34664 67984 34664 0 net20
rlabel metal2 65352 4760 65352 4760 0 net200
rlabel metal2 70000 3528 70000 3528 0 net201
rlabel metal2 76328 6496 76328 6496 0 net202
rlabel metal2 77560 3584 77560 3584 0 net203
rlabel metal2 90776 7448 90776 7448 0 net204
rlabel metal2 94472 7504 94472 7504 0 net205
rlabel metal2 95368 8064 95368 8064 0 net206
rlabel metal2 93240 3584 93240 3584 0 net207
rlabel metal3 98000 3528 98000 3528 0 net208
rlabel metal2 20720 3528 20720 3528 0 net209
rlabel metal2 69720 33264 69720 33264 0 net21
rlabel metal2 101304 3640 101304 3640 0 net210
rlabel metal2 109032 3472 109032 3472 0 net211
rlabel metal2 116760 5040 116760 5040 0 net212
rlabel metal2 114856 4760 114856 4760 0 net213
rlabel metal2 117208 4928 117208 4928 0 net214
rlabel metal2 121464 3584 121464 3584 0 net215
rlabel metal3 123144 5096 123144 5096 0 net216
rlabel metal2 138712 6048 138712 6048 0 net217
rlabel metal3 129696 4200 129696 4200 0 net218
rlabel metal2 135800 6664 135800 6664 0 net219
rlabel metal2 70840 36008 70840 36008 0 net22
rlabel metal3 27608 5208 27608 5208 0 net220
rlabel metal2 124376 7504 124376 7504 0 net221
rlabel metal3 125384 8344 125384 8344 0 net222
rlabel metal2 31416 6160 31416 6160 0 net223
rlabel metal2 47320 5600 47320 5600 0 net224
rlabel metal2 44744 4984 44744 4984 0 net225
rlabel metal2 45080 3864 45080 3864 0 net226
rlabel metal2 55272 5264 55272 5264 0 net227
rlabel metal2 52920 5152 52920 5152 0 net228
rlabel metal2 58128 7336 58128 7336 0 net229
rlabel metal2 29064 34496 29064 34496 0 net23
rlabel metal2 7000 36176 7000 36176 0 net230
rlabel metal3 76776 34888 76776 34888 0 net231
rlabel metal2 8792 34832 8792 34832 0 net232
rlabel metal2 12600 35616 12600 35616 0 net233
rlabel metal2 16016 34776 16016 34776 0 net234
rlabel metal2 18312 35840 18312 35840 0 net235
rlabel metal2 23128 37184 23128 37184 0 net236
rlabel metal3 60144 29288 60144 29288 0 net237
rlabel metal3 85456 35784 85456 35784 0 net238
rlabel metal2 91056 34328 91056 34328 0 net239
rlabel metal2 73304 35056 73304 35056 0 net24
rlabel metal2 4760 36344 4760 36344 0 net240
rlabel metal2 75656 34608 75656 34608 0 net241
rlabel metal2 73976 36120 73976 36120 0 net25
rlabel metal2 29400 34608 29400 34608 0 net26
rlabel metal2 23128 35000 23128 35000 0 net27
rlabel metal2 25816 35784 25816 35784 0 net28
rlabel metal2 28448 34328 28448 34328 0 net29
rlabel metal2 38584 33096 38584 33096 0 net3
rlabel metal2 31192 33768 31192 33768 0 net30
rlabel metal3 47600 31864 47600 31864 0 net31
rlabel metal2 33880 36680 33880 36680 0 net32
rlabel metal2 28392 30352 28392 30352 0 net33
rlabel metal2 67480 33264 67480 33264 0 net34
rlabel metal2 67816 34328 67816 34328 0 net35
rlabel metal2 77560 35840 77560 35840 0 net36
rlabel metal3 77840 34328 77840 34328 0 net37
rlabel metal3 92792 36344 92792 36344 0 net38
rlabel metal2 93016 36176 93016 36176 0 net39
rlabel metal3 74704 33992 74704 33992 0 net4
rlabel metal2 96040 33600 96040 33600 0 net40
rlabel metal2 97272 36400 97272 36400 0 net41
rlabel metal2 106456 36400 106456 36400 0 net42
rlabel metal2 108808 34720 108808 34720 0 net43
rlabel metal2 24248 35728 24248 35728 0 net44
rlabel metal2 110152 34944 110152 34944 0 net45
rlabel metal2 110824 33712 110824 33712 0 net46
rlabel metal3 128240 34104 128240 34104 0 net47
rlabel metal2 125160 34888 125160 34888 0 net48
rlabel metal2 133000 35224 133000 35224 0 net49
rlabel metal2 76104 32872 76104 32872 0 net5
rlabel metal2 135688 35672 135688 35672 0 net50
rlabel metal2 137592 36176 137592 36176 0 net51
rlabel metal3 138936 35896 138936 35896 0 net52
rlabel metal2 139832 35112 139832 35112 0 net53
rlabel metal2 141960 34944 141960 34944 0 net54
rlabel metal3 59528 26376 59528 26376 0 net55
rlabel metal2 76776 34888 76776 34888 0 net56
rlabel metal2 75096 36792 75096 36792 0 net57
rlabel metal2 30184 37240 30184 37240 0 net58
rlabel metal2 47544 36344 47544 36344 0 net59
rlabel metal2 44632 30408 44632 30408 0 net6
rlabel metal2 44576 35448 44576 35448 0 net60
rlabel metal2 53816 36176 53816 36176 0 net61
rlabel metal2 52696 36176 52696 36176 0 net62
rlabel metal2 64232 32928 64232 32928 0 net63
rlabel metal3 64288 33432 64288 33432 0 net64
rlabel metal2 71400 12880 71400 12880 0 net65
rlabel metal2 60256 4984 60256 4984 0 net66
rlabel metal2 23800 3248 23800 3248 0 net67
rlabel metal3 27776 3304 27776 3304 0 net68
rlabel metal2 13048 34832 13048 34832 0 net69
rlabel metal2 48552 33712 48552 33712 0 net7
rlabel metal2 37968 3304 37968 3304 0 net70
rlabel metal2 21784 33936 21784 33936 0 net71
rlabel metal3 47768 3304 47768 3304 0 net72
rlabel metal2 27160 33768 27160 33768 0 net73
rlabel metal2 29904 34328 29904 34328 0 net74
rlabel metal2 8680 3920 8680 3920 0 net75
rlabel metal2 7896 35000 7896 35000 0 net76
rlabel metal2 58632 3024 58632 3024 0 net77
rlabel metal2 67312 3304 67312 3304 0 net78
rlabel metal3 71456 4984 71456 4984 0 net79
rlabel metal2 46088 36120 46088 36120 0 net8
rlabel metal2 74200 3080 74200 3080 0 net80
rlabel metal2 78176 3304 78176 3304 0 net81
rlabel metal3 47936 33992 47936 33992 0 net82
rlabel metal2 46088 24780 46088 24780 0 net83
rlabel metal2 48720 35560 48720 35560 0 net84
rlabel metal2 94136 3248 94136 3248 0 net85
rlabel metal2 55216 33992 55216 33992 0 net86
rlabel metal2 20664 33544 20664 33544 0 net87
rlabel metal3 98896 3304 98896 3304 0 net88
rlabel metal2 105896 3136 105896 3136 0 net89
rlabel metal2 50008 34720 50008 34720 0 net9
rlabel metal2 110320 3304 110320 3304 0 net90
rlabel metal2 114296 5040 114296 5040 0 net91
rlabel metal2 117880 7252 117880 7252 0 net92
rlabel metal2 122360 4704 122360 4704 0 net93
rlabel metal2 126448 3304 126448 3304 0 net94
rlabel metal2 130480 3304 130480 3304 0 net95
rlabel metal2 119336 33880 119336 33880 0 net96
rlabel metal3 139664 4536 139664 4536 0 net97
rlabel metal2 26488 6888 26488 6888 0 net98
rlabel metal3 96600 34776 96600 34776 0 net99
rlabel metal2 20664 4256 20664 4256 0 operation
rlabel metal2 54040 34664 54040 34664 0 web_mem
rlabel metal2 5992 37184 5992 37184 0 web_mem0
rlabel metal3 77168 35000 77168 35000 0 web_mem1
rlabel metal2 10136 35056 10136 35056 0 wmask_mem0[0]
rlabel metal2 12152 37184 12152 37184 0 wmask_mem0[1]
rlabel metal2 16352 35560 16352 35560 0 wmask_mem0[2]
rlabel metal2 20328 34944 20328 34944 0 wmask_mem0[3]
rlabel metal2 82712 35896 82712 35896 0 wmask_mem1[0]
rlabel metal2 84840 36680 84840 36680 0 wmask_mem1[1]
rlabel metal3 87528 35560 87528 35560 0 wmask_mem1[2]
rlabel metal2 91896 35784 91896 35784 0 wmask_mem1[3]
<< properties >>
string FIXED_BBOX 0 0 150000 40000
<< end >>
