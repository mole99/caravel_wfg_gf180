magic
tech gf180mcuC
magscale 1 10
timestamp 1670096752
<< metal1 >>
rect 82562 37326 82574 37378
rect 82626 37375 82638 37378
rect 83794 37375 83806 37378
rect 82626 37329 83806 37375
rect 82626 37326 82638 37329
rect 83794 37326 83806 37329
rect 83858 37326 83870 37378
rect 1344 36874 148624 36908
rect 1344 36822 19624 36874
rect 19676 36822 19728 36874
rect 19780 36822 19832 36874
rect 19884 36822 56444 36874
rect 56496 36822 56548 36874
rect 56600 36822 56652 36874
rect 56704 36822 93264 36874
rect 93316 36822 93368 36874
rect 93420 36822 93472 36874
rect 93524 36822 130084 36874
rect 130136 36822 130188 36874
rect 130240 36822 130292 36874
rect 130344 36822 148624 36874
rect 1344 36788 148624 36822
rect 77534 36706 77586 36718
rect 40786 36654 40798 36706
rect 40850 36703 40862 36706
rect 41346 36703 41358 36706
rect 40850 36657 41358 36703
rect 40850 36654 40862 36657
rect 41346 36654 41358 36657
rect 41410 36654 41422 36706
rect 77534 36642 77586 36654
rect 13918 36594 13970 36606
rect 27694 36594 27746 36606
rect 67678 36594 67730 36606
rect 8866 36542 8878 36594
rect 8930 36542 8942 36594
rect 12786 36542 12798 36594
rect 12850 36542 12862 36594
rect 16706 36542 16718 36594
rect 16770 36542 16782 36594
rect 20626 36542 20638 36594
rect 20690 36542 20702 36594
rect 24210 36542 24222 36594
rect 24274 36542 24286 36594
rect 26898 36542 26910 36594
rect 26962 36542 26974 36594
rect 32274 36542 32286 36594
rect 32338 36542 32350 36594
rect 36306 36542 36318 36594
rect 36370 36542 36382 36594
rect 40226 36542 40238 36594
rect 40290 36542 40302 36594
rect 43922 36542 43934 36594
rect 43986 36542 43998 36594
rect 48066 36542 48078 36594
rect 48130 36542 48142 36594
rect 51986 36542 51998 36594
rect 52050 36542 52062 36594
rect 55682 36542 55694 36594
rect 55746 36542 55758 36594
rect 59714 36542 59726 36594
rect 59778 36542 59790 36594
rect 63634 36542 63646 36594
rect 63698 36542 63710 36594
rect 64754 36542 64766 36594
rect 64818 36542 64830 36594
rect 67218 36542 67230 36594
rect 67282 36542 67294 36594
rect 13918 36530 13970 36542
rect 27694 36530 27746 36542
rect 67678 36530 67730 36542
rect 68462 36594 68514 36606
rect 71710 36594 71762 36606
rect 77198 36594 77250 36606
rect 92766 36594 92818 36606
rect 122222 36594 122274 36606
rect 70802 36542 70814 36594
rect 70866 36542 70878 36594
rect 75506 36542 75518 36594
rect 75570 36542 75582 36594
rect 78978 36542 78990 36594
rect 79042 36542 79054 36594
rect 80210 36542 80222 36594
rect 80274 36542 80286 36594
rect 85810 36542 85822 36594
rect 85874 36542 85886 36594
rect 89730 36542 89742 36594
rect 89794 36542 89806 36594
rect 93538 36542 93550 36594
rect 93602 36542 93614 36594
rect 96226 36542 96238 36594
rect 96290 36542 96302 36594
rect 99810 36542 99822 36594
rect 99874 36542 99886 36594
rect 104402 36542 104414 36594
rect 104466 36542 104478 36594
rect 107874 36542 107886 36594
rect 107938 36542 107950 36594
rect 111570 36542 111582 36594
rect 111634 36542 111646 36594
rect 115490 36542 115502 36594
rect 115554 36542 115566 36594
rect 119410 36542 119422 36594
rect 119474 36542 119486 36594
rect 123330 36542 123342 36594
rect 123394 36542 123406 36594
rect 129042 36542 129054 36594
rect 129106 36542 129118 36594
rect 132626 36542 132638 36594
rect 132690 36542 132702 36594
rect 135090 36542 135102 36594
rect 135154 36542 135166 36594
rect 139010 36542 139022 36594
rect 139074 36542 139086 36594
rect 144162 36542 144174 36594
rect 144226 36542 144238 36594
rect 147522 36542 147534 36594
rect 147586 36542 147598 36594
rect 68462 36530 68514 36542
rect 71710 36530 71762 36542
rect 77198 36530 77250 36542
rect 92766 36530 92818 36542
rect 122222 36530 122274 36542
rect 33518 36482 33570 36494
rect 6626 36430 6638 36482
rect 6690 36430 6702 36482
rect 33518 36418 33570 36430
rect 37438 36482 37490 36494
rect 49198 36482 49250 36494
rect 45938 36430 45950 36482
rect 46002 36430 46014 36482
rect 37438 36418 37490 36430
rect 49198 36418 49250 36430
rect 53118 36482 53170 36494
rect 73502 36482 73554 36494
rect 89070 36482 89122 36494
rect 102734 36482 102786 36494
rect 53778 36430 53790 36482
rect 53842 36430 53854 36482
rect 65090 36430 65102 36482
rect 65154 36430 65166 36482
rect 78194 36430 78206 36482
rect 78258 36430 78270 36482
rect 88386 36430 88398 36482
rect 88450 36430 88462 36482
rect 98354 36430 98366 36482
rect 98418 36430 98430 36482
rect 53118 36418 53170 36430
rect 73502 36418 73554 36430
rect 89070 36418 89122 36430
rect 102734 36418 102786 36430
rect 103630 36482 103682 36494
rect 103630 36418 103682 36430
rect 106878 36482 106930 36494
rect 141822 36482 141874 36494
rect 129826 36430 129838 36482
rect 129890 36430 129902 36482
rect 106878 36418 106930 36430
rect 141822 36418 141874 36430
rect 145742 36482 145794 36494
rect 146850 36430 146862 36482
rect 146914 36430 146926 36482
rect 145742 36418 145794 36430
rect 4846 36370 4898 36382
rect 10782 36370 10834 36382
rect 14702 36370 14754 36382
rect 18286 36370 18338 36382
rect 21422 36370 21474 36382
rect 7858 36318 7870 36370
rect 7922 36318 7934 36370
rect 11666 36318 11678 36370
rect 11730 36318 11742 36370
rect 15362 36318 15374 36370
rect 15426 36318 15438 36370
rect 19282 36318 19294 36370
rect 19346 36318 19358 36370
rect 4846 36306 4898 36318
rect 10782 36306 10834 36318
rect 14702 36306 14754 36318
rect 18286 36306 18338 36318
rect 21422 36306 21474 36318
rect 22206 36370 22258 36382
rect 28142 36370 28194 36382
rect 22866 36318 22878 36370
rect 22930 36318 22942 36370
rect 25554 36318 25566 36370
rect 25618 36318 25630 36370
rect 22206 36306 22258 36318
rect 28142 36306 28194 36318
rect 29262 36370 29314 36382
rect 29262 36306 29314 36318
rect 29822 36370 29874 36382
rect 34302 36370 34354 36382
rect 38222 36370 38274 36382
rect 41918 36370 41970 36382
rect 45278 36370 45330 36382
rect 49646 36370 49698 36382
rect 57486 36370 57538 36382
rect 60846 36370 60898 36382
rect 30930 36318 30942 36370
rect 30994 36318 31006 36370
rect 35074 36318 35086 36370
rect 35138 36318 35150 36370
rect 38882 36318 38894 36370
rect 38946 36318 38958 36370
rect 42578 36318 42590 36370
rect 42642 36318 42654 36370
rect 46834 36318 46846 36370
rect 46898 36318 46910 36370
rect 50978 36318 50990 36370
rect 51042 36318 51054 36370
rect 54786 36318 54798 36370
rect 54850 36318 54862 36370
rect 58482 36318 58494 36370
rect 58546 36318 58558 36370
rect 29822 36306 29874 36318
rect 34302 36306 34354 36318
rect 38222 36306 38274 36318
rect 41918 36306 41970 36318
rect 45278 36306 45330 36318
rect 49646 36306 49698 36318
rect 57486 36306 57538 36318
rect 60846 36306 60898 36318
rect 61630 36370 61682 36382
rect 68910 36370 68962 36382
rect 72382 36370 72434 36382
rect 62290 36318 62302 36370
rect 62354 36318 62366 36370
rect 65874 36318 65886 36370
rect 65938 36318 65950 36370
rect 69458 36318 69470 36370
rect 69522 36318 69534 36370
rect 61630 36306 61682 36318
rect 68910 36306 68962 36318
rect 72382 36306 72434 36318
rect 73166 36370 73218 36382
rect 82238 36370 82290 36382
rect 74498 36318 74510 36370
rect 74562 36318 74574 36370
rect 76402 36318 76414 36370
rect 76466 36318 76478 36370
rect 76850 36318 76862 36370
rect 76914 36318 76926 36370
rect 81218 36318 81230 36370
rect 81282 36318 81294 36370
rect 73166 36306 73218 36318
rect 82238 36306 82290 36318
rect 82574 36370 82626 36382
rect 82574 36306 82626 36318
rect 83022 36370 83074 36382
rect 83022 36306 83074 36318
rect 84142 36370 84194 36382
rect 91982 36370 92034 36382
rect 99038 36370 99090 36382
rect 109902 36370 109954 36382
rect 86818 36318 86830 36370
rect 86882 36318 86894 36370
rect 90738 36318 90750 36370
rect 90802 36318 90814 36370
rect 94546 36318 94558 36370
rect 94610 36318 94622 36370
rect 97458 36318 97470 36370
rect 97522 36318 97534 36370
rect 100818 36318 100830 36370
rect 100882 36318 100894 36370
rect 105298 36318 105310 36370
rect 105362 36318 105374 36370
rect 108882 36318 108894 36370
rect 108946 36318 108958 36370
rect 84142 36306 84194 36318
rect 91982 36306 92034 36318
rect 99038 36306 99090 36318
rect 109902 36306 109954 36318
rect 110238 36370 110290 36382
rect 113598 36370 113650 36382
rect 112578 36318 112590 36370
rect 112642 36318 112654 36370
rect 110238 36306 110290 36318
rect 113598 36306 113650 36318
rect 114382 36370 114434 36382
rect 117518 36370 117570 36382
rect 116498 36318 116510 36370
rect 116562 36318 116574 36370
rect 114382 36306 114434 36318
rect 117518 36306 117570 36318
rect 118302 36370 118354 36382
rect 121774 36370 121826 36382
rect 125358 36370 125410 36382
rect 120418 36318 120430 36370
rect 120482 36318 120494 36370
rect 124338 36318 124350 36370
rect 124402 36318 124414 36370
rect 118302 36306 118354 36318
rect 121774 36306 121826 36318
rect 125358 36306 125410 36318
rect 125694 36370 125746 36382
rect 125694 36306 125746 36318
rect 126142 36370 126194 36382
rect 130398 36370 130450 36382
rect 133534 36370 133586 36382
rect 137118 36370 137170 36382
rect 142158 36370 142210 36382
rect 145294 36370 145346 36382
rect 127698 36318 127710 36370
rect 127762 36318 127774 36370
rect 131282 36318 131294 36370
rect 131346 36318 131358 36370
rect 136098 36318 136110 36370
rect 136162 36318 136174 36370
rect 140018 36318 140030 36370
rect 140082 36318 140094 36370
rect 143042 36318 143054 36370
rect 143106 36318 143118 36370
rect 126142 36306 126194 36318
rect 130398 36306 130450 36318
rect 133534 36306 133586 36318
rect 137118 36306 137170 36318
rect 142158 36306 142210 36318
rect 145294 36306 145346 36318
rect 6078 36258 6130 36270
rect 6078 36194 6130 36206
rect 6862 36258 6914 36270
rect 6862 36194 6914 36206
rect 9998 36258 10050 36270
rect 9998 36194 10050 36206
rect 10446 36258 10498 36270
rect 10446 36194 10498 36206
rect 14366 36258 14418 36270
rect 14366 36194 14418 36206
rect 17838 36258 17890 36270
rect 17838 36194 17890 36206
rect 18622 36258 18674 36270
rect 18622 36194 18674 36206
rect 21870 36258 21922 36270
rect 21870 36194 21922 36206
rect 28478 36258 28530 36270
rect 28478 36194 28530 36206
rect 30158 36258 30210 36270
rect 30158 36194 30210 36206
rect 33966 36258 34018 36270
rect 33966 36194 34018 36206
rect 37886 36258 37938 36270
rect 37886 36194 37938 36206
rect 41134 36258 41186 36270
rect 41134 36194 41186 36206
rect 41582 36258 41634 36270
rect 41582 36194 41634 36206
rect 45726 36258 45778 36270
rect 45726 36194 45778 36206
rect 49982 36258 50034 36270
rect 49982 36194 50034 36206
rect 53566 36258 53618 36270
rect 53566 36194 53618 36206
rect 57038 36258 57090 36270
rect 57038 36194 57090 36206
rect 57822 36258 57874 36270
rect 57822 36194 57874 36206
rect 61294 36258 61346 36270
rect 61294 36194 61346 36206
rect 72494 36258 72546 36270
rect 72494 36194 72546 36206
rect 72718 36258 72770 36270
rect 72718 36194 72770 36206
rect 84478 36258 84530 36270
rect 84478 36194 84530 36206
rect 84926 36258 84978 36270
rect 84926 36194 84978 36206
rect 88622 36258 88674 36270
rect 88622 36194 88674 36206
rect 92318 36258 92370 36270
rect 92318 36194 92370 36206
rect 98590 36258 98642 36270
rect 98590 36194 98642 36206
rect 102174 36258 102226 36270
rect 102174 36194 102226 36206
rect 106318 36258 106370 36270
rect 106318 36194 106370 36206
rect 110686 36258 110738 36270
rect 110686 36194 110738 36206
rect 113934 36258 113986 36270
rect 113934 36194 113986 36206
rect 117854 36258 117906 36270
rect 117854 36194 117906 36206
rect 121438 36258 121490 36270
rect 121438 36194 121490 36206
rect 129614 36258 129666 36270
rect 129614 36194 129666 36206
rect 133198 36258 133250 36270
rect 133198 36194 133250 36206
rect 133982 36258 134034 36270
rect 133982 36194 134034 36206
rect 137454 36258 137506 36270
rect 137454 36194 137506 36206
rect 138014 36258 138066 36270
rect 138014 36194 138066 36206
rect 140926 36258 140978 36270
rect 140926 36194 140978 36206
rect 144958 36258 145010 36270
rect 144958 36194 145010 36206
rect 1344 36090 148784 36124
rect 1344 36038 38034 36090
rect 38086 36038 38138 36090
rect 38190 36038 38242 36090
rect 38294 36038 74854 36090
rect 74906 36038 74958 36090
rect 75010 36038 75062 36090
rect 75114 36038 111674 36090
rect 111726 36038 111778 36090
rect 111830 36038 111882 36090
rect 111934 36038 148494 36090
rect 148546 36038 148598 36090
rect 148650 36038 148702 36090
rect 148754 36038 148784 36090
rect 1344 36004 148784 36038
rect 9662 35922 9714 35934
rect 9662 35858 9714 35870
rect 21422 35922 21474 35934
rect 21422 35858 21474 35870
rect 35758 35922 35810 35934
rect 35758 35858 35810 35870
rect 43598 35922 43650 35934
rect 43598 35858 43650 35870
rect 48414 35922 48466 35934
rect 48414 35858 48466 35870
rect 59502 35922 59554 35934
rect 59502 35858 59554 35870
rect 69694 35922 69746 35934
rect 69694 35858 69746 35870
rect 100382 35922 100434 35934
rect 100382 35858 100434 35870
rect 105086 35922 105138 35934
rect 105086 35858 105138 35870
rect 132190 35922 132242 35934
rect 132190 35858 132242 35870
rect 146862 35922 146914 35934
rect 146862 35858 146914 35870
rect 32510 35810 32562 35822
rect 36542 35810 36594 35822
rect 52222 35810 52274 35822
rect 70254 35810 70306 35822
rect 81678 35810 81730 35822
rect 97918 35810 97970 35822
rect 104078 35810 104130 35822
rect 108446 35810 108498 35822
rect 17826 35758 17838 35810
rect 17890 35758 17902 35810
rect 19730 35758 19742 35810
rect 19794 35758 19806 35810
rect 21970 35758 21982 35810
rect 22034 35758 22046 35810
rect 28242 35758 28254 35810
rect 28306 35758 28318 35810
rect 30594 35758 30606 35810
rect 30658 35758 30670 35810
rect 33730 35758 33742 35810
rect 33794 35758 33806 35810
rect 37202 35758 37214 35810
rect 37266 35758 37278 35810
rect 39330 35758 39342 35810
rect 39394 35758 39406 35810
rect 41682 35758 41694 35810
rect 41746 35758 41758 35810
rect 44146 35758 44158 35810
rect 44210 35758 44222 35810
rect 46162 35758 46174 35810
rect 46226 35758 46238 35810
rect 49746 35758 49758 35810
rect 49810 35758 49822 35810
rect 53330 35758 53342 35810
rect 53394 35758 53406 35810
rect 55570 35758 55582 35810
rect 55634 35758 55646 35810
rect 57586 35758 57598 35810
rect 57650 35758 57662 35810
rect 60498 35758 60510 35810
rect 60562 35758 60574 35810
rect 63634 35758 63646 35810
rect 63698 35758 63710 35810
rect 65650 35758 65662 35810
rect 65714 35758 65726 35810
rect 67666 35758 67678 35810
rect 67730 35758 67742 35810
rect 71250 35758 71262 35810
rect 71314 35758 71326 35810
rect 73490 35758 73502 35810
rect 73554 35758 73566 35810
rect 75618 35758 75630 35810
rect 75682 35758 75694 35810
rect 76066 35758 76078 35810
rect 76130 35758 76142 35810
rect 83794 35758 83806 35810
rect 83858 35758 83870 35810
rect 84914 35758 84926 35810
rect 84978 35758 84990 35810
rect 86706 35758 86718 35810
rect 86770 35758 86782 35810
rect 89506 35758 89518 35810
rect 89570 35758 89582 35810
rect 89954 35758 89966 35810
rect 90018 35758 90030 35810
rect 91410 35758 91422 35810
rect 91474 35758 91486 35810
rect 93314 35758 93326 35810
rect 93378 35758 93390 35810
rect 93762 35758 93774 35810
rect 93826 35758 93838 35810
rect 98690 35758 98702 35810
rect 98754 35758 98766 35810
rect 102610 35758 102622 35810
rect 102674 35758 102686 35810
rect 107090 35758 107102 35810
rect 107154 35758 107166 35810
rect 32510 35746 32562 35758
rect 36542 35746 36594 35758
rect 52222 35746 52274 35758
rect 70254 35746 70306 35758
rect 81678 35746 81730 35758
rect 97918 35746 97970 35758
rect 104078 35746 104130 35758
rect 108446 35746 108498 35758
rect 108894 35810 108946 35822
rect 111694 35810 111746 35822
rect 110898 35758 110910 35810
rect 110962 35758 110974 35810
rect 108894 35746 108946 35758
rect 111694 35746 111746 35758
rect 112030 35810 112082 35822
rect 115614 35810 115666 35822
rect 114258 35758 114270 35810
rect 114322 35758 114334 35810
rect 112030 35746 112082 35758
rect 115614 35746 115666 35758
rect 116062 35810 116114 35822
rect 123118 35810 123170 35822
rect 131406 35810 131458 35822
rect 139358 35810 139410 35822
rect 117842 35758 117854 35810
rect 117906 35758 117918 35810
rect 119186 35758 119198 35810
rect 119250 35758 119262 35810
rect 122098 35758 122110 35810
rect 122162 35758 122174 35810
rect 125010 35758 125022 35810
rect 125074 35758 125086 35810
rect 126130 35758 126142 35810
rect 126194 35758 126206 35810
rect 129490 35758 129502 35810
rect 129554 35758 129566 35810
rect 133970 35758 133982 35810
rect 134034 35758 134046 35810
rect 138002 35758 138014 35810
rect 138066 35758 138078 35810
rect 140242 35758 140254 35810
rect 140306 35758 140318 35810
rect 142930 35758 142942 35810
rect 142994 35758 143006 35810
rect 143154 35758 143166 35810
rect 143218 35758 143230 35810
rect 146178 35758 146190 35810
rect 146242 35758 146254 35810
rect 116062 35746 116114 35758
rect 123118 35746 123170 35758
rect 131406 35746 131458 35758
rect 139358 35746 139410 35758
rect 20414 35698 20466 35710
rect 32846 35698 32898 35710
rect 7186 35646 7198 35698
rect 7250 35646 7262 35698
rect 8978 35646 8990 35698
rect 9042 35646 9054 35698
rect 10434 35646 10446 35698
rect 10498 35646 10510 35698
rect 13346 35646 13358 35698
rect 13410 35646 13422 35698
rect 14130 35646 14142 35698
rect 14194 35646 14206 35698
rect 16930 35646 16942 35698
rect 16994 35646 17006 35698
rect 18946 35646 18958 35698
rect 19010 35646 19022 35698
rect 19618 35646 19630 35698
rect 19682 35646 19694 35698
rect 23090 35646 23102 35698
rect 23154 35646 23166 35698
rect 24770 35646 24782 35698
rect 24834 35646 24846 35698
rect 27570 35646 27582 35698
rect 27634 35646 27646 35698
rect 30818 35646 30830 35698
rect 30882 35646 30894 35698
rect 20414 35634 20466 35646
rect 32846 35634 32898 35646
rect 36206 35698 36258 35710
rect 48750 35698 48802 35710
rect 59838 35698 59890 35710
rect 70590 35698 70642 35710
rect 81342 35698 81394 35710
rect 88286 35698 88338 35710
rect 39218 35646 39230 35698
rect 39282 35646 39294 35698
rect 56466 35646 56478 35698
rect 56530 35646 56542 35698
rect 65538 35646 65550 35698
rect 65602 35646 65614 35698
rect 77298 35646 77310 35698
rect 77362 35646 77374 35698
rect 79090 35646 79102 35698
rect 79154 35646 79166 35698
rect 85810 35646 85822 35698
rect 85874 35646 85886 35698
rect 87602 35646 87614 35698
rect 87666 35646 87678 35698
rect 36206 35634 36258 35646
rect 48750 35634 48802 35646
rect 59838 35634 59890 35646
rect 70590 35634 70642 35646
rect 81342 35634 81394 35646
rect 88286 35634 88338 35646
rect 90190 35698 90242 35710
rect 97582 35698 97634 35710
rect 100942 35698 100994 35710
rect 91298 35646 91310 35698
rect 91362 35646 91374 35698
rect 94994 35646 95006 35698
rect 95058 35646 95070 35698
rect 98578 35646 98590 35698
rect 98642 35646 98654 35698
rect 90190 35634 90242 35646
rect 97582 35634 97634 35646
rect 100942 35634 100994 35646
rect 103742 35698 103794 35710
rect 103742 35634 103794 35646
rect 105534 35698 105586 35710
rect 105534 35634 105586 35646
rect 108110 35698 108162 35710
rect 108110 35634 108162 35646
rect 115278 35698 115330 35710
rect 123454 35698 123506 35710
rect 139022 35698 139074 35710
rect 119074 35646 119086 35698
rect 119138 35646 119150 35698
rect 131618 35646 131630 35698
rect 131682 35646 131694 35698
rect 134978 35646 134990 35698
rect 135042 35646 135054 35698
rect 115278 35634 115330 35646
rect 123454 35634 123506 35646
rect 139022 35634 139074 35646
rect 142606 35698 142658 35710
rect 142606 35634 142658 35646
rect 25566 35586 25618 35598
rect 52670 35586 52722 35598
rect 62638 35586 62690 35598
rect 82126 35586 82178 35598
rect 92094 35586 92146 35598
rect 127934 35586 127986 35598
rect 143950 35586 144002 35598
rect 6402 35534 6414 35586
rect 6466 35534 6478 35586
rect 8306 35534 8318 35586
rect 8370 35534 8382 35586
rect 10994 35534 11006 35586
rect 11058 35534 11070 35586
rect 12674 35534 12686 35586
rect 12738 35534 12750 35586
rect 14578 35534 14590 35586
rect 14642 35534 14654 35586
rect 16258 35534 16270 35586
rect 16322 35534 16334 35586
rect 24210 35534 24222 35586
rect 24274 35534 24286 35586
rect 26786 35534 26798 35586
rect 26850 35534 26862 35586
rect 29586 35534 29598 35586
rect 29650 35534 29662 35586
rect 34850 35534 34862 35586
rect 34914 35534 34926 35586
rect 38546 35534 38558 35586
rect 38610 35534 38622 35586
rect 43026 35534 43038 35586
rect 43090 35534 43102 35586
rect 45490 35534 45502 35586
rect 45554 35534 45566 35586
rect 47282 35534 47294 35586
rect 47346 35534 47358 35586
rect 51090 35534 51102 35586
rect 51154 35534 51166 35586
rect 54450 35534 54462 35586
rect 54514 35534 54526 35586
rect 58930 35534 58942 35586
rect 58994 35534 59006 35586
rect 61618 35534 61630 35586
rect 61682 35534 61694 35586
rect 64642 35534 64654 35586
rect 64706 35534 64718 35586
rect 69010 35534 69022 35586
rect 69074 35534 69086 35586
rect 72370 35534 72382 35586
rect 72434 35534 72446 35586
rect 74834 35534 74846 35586
rect 74898 35534 74910 35586
rect 78082 35534 78094 35586
rect 78146 35534 78158 35586
rect 79762 35534 79774 35586
rect 79826 35534 79838 35586
rect 82786 35534 82798 35586
rect 82850 35534 82862 35586
rect 87826 35534 87838 35586
rect 87890 35583 87902 35586
rect 88162 35583 88174 35586
rect 87890 35537 88174 35583
rect 87890 35534 87902 35537
rect 88162 35534 88174 35537
rect 88226 35534 88238 35586
rect 95890 35534 95902 35586
rect 95954 35534 95966 35586
rect 101602 35534 101614 35586
rect 101666 35534 101678 35586
rect 106082 35534 106094 35586
rect 106146 35534 106158 35586
rect 109666 35534 109678 35586
rect 109730 35534 109742 35586
rect 113250 35534 113262 35586
rect 113314 35534 113326 35586
rect 116834 35534 116846 35586
rect 116898 35534 116910 35586
rect 121090 35534 121102 35586
rect 121154 35534 121166 35586
rect 124002 35534 124014 35586
rect 124066 35534 124078 35586
rect 127474 35534 127486 35586
rect 127538 35534 127550 35586
rect 130610 35534 130622 35586
rect 130674 35534 130686 35586
rect 132962 35534 132974 35586
rect 133026 35534 133038 35586
rect 135650 35534 135662 35586
rect 135714 35534 135726 35586
rect 136994 35534 137006 35586
rect 137058 35534 137070 35586
rect 141586 35534 141598 35586
rect 141650 35534 141662 35586
rect 144946 35534 144958 35586
rect 145010 35534 145022 35586
rect 25566 35522 25618 35534
rect 52670 35522 52722 35534
rect 62638 35522 62690 35534
rect 82126 35522 82178 35534
rect 92094 35522 92146 35534
rect 127934 35522 127986 35534
rect 143950 35522 144002 35534
rect 20750 35474 20802 35486
rect 20750 35410 20802 35422
rect 31278 35474 31330 35486
rect 31278 35410 31330 35422
rect 31614 35474 31666 35486
rect 31614 35410 31666 35422
rect 40014 35474 40066 35486
rect 40014 35410 40066 35422
rect 40350 35474 40402 35486
rect 40350 35410 40402 35422
rect 51662 35474 51714 35486
rect 51662 35410 51714 35422
rect 51998 35474 52050 35486
rect 51998 35410 52050 35422
rect 66334 35474 66386 35486
rect 66334 35410 66386 35422
rect 66670 35474 66722 35486
rect 66670 35410 66722 35422
rect 76302 35474 76354 35486
rect 76302 35410 76354 35422
rect 76638 35474 76690 35486
rect 76638 35410 76690 35422
rect 90526 35474 90578 35486
rect 90526 35410 90578 35422
rect 92430 35474 92482 35486
rect 92430 35410 92482 35422
rect 93998 35474 94050 35486
rect 93998 35410 94050 35422
rect 94334 35474 94386 35486
rect 94334 35410 94386 35422
rect 99374 35474 99426 35486
rect 99374 35410 99426 35422
rect 99710 35474 99762 35486
rect 99710 35410 99762 35422
rect 119870 35474 119922 35486
rect 119870 35410 119922 35422
rect 120206 35474 120258 35486
rect 120206 35410 120258 35422
rect 142270 35474 142322 35486
rect 142270 35410 142322 35422
rect 1344 35306 148624 35340
rect 1344 35254 19624 35306
rect 19676 35254 19728 35306
rect 19780 35254 19832 35306
rect 19884 35254 56444 35306
rect 56496 35254 56548 35306
rect 56600 35254 56652 35306
rect 56704 35254 93264 35306
rect 93316 35254 93368 35306
rect 93420 35254 93472 35306
rect 93524 35254 130084 35306
rect 130136 35254 130188 35306
rect 130240 35254 130292 35306
rect 130344 35254 148624 35306
rect 1344 35220 148624 35254
rect 30046 35138 30098 35150
rect 30046 35074 30098 35086
rect 49758 35138 49810 35150
rect 49758 35074 49810 35086
rect 52670 35138 52722 35150
rect 52670 35074 52722 35086
rect 68126 35138 68178 35150
rect 68126 35074 68178 35086
rect 120654 35138 120706 35150
rect 120654 35074 120706 35086
rect 123118 35138 123170 35150
rect 123118 35074 123170 35086
rect 130734 35138 130786 35150
rect 130734 35074 130786 35086
rect 138798 35138 138850 35150
rect 138798 35074 138850 35086
rect 12910 35026 12962 35038
rect 38446 35026 38498 35038
rect 88958 35026 89010 35038
rect 100270 35026 100322 35038
rect 121550 35026 121602 35038
rect 5842 34974 5854 35026
rect 5906 34974 5918 35026
rect 6962 34974 6974 35026
rect 7026 35023 7038 35026
rect 7522 35023 7534 35026
rect 7026 34977 7534 35023
rect 7026 34974 7038 34977
rect 7522 34974 7534 34977
rect 7586 34974 7598 35026
rect 8418 34974 8430 35026
rect 8482 34974 8494 35026
rect 10322 34974 10334 35026
rect 10386 34974 10398 35026
rect 13906 34974 13918 35026
rect 13970 34974 13982 35026
rect 17154 34974 17166 35026
rect 17218 34974 17230 35026
rect 21858 34974 21870 35026
rect 21922 34974 21934 35026
rect 23762 34974 23774 35026
rect 23826 34974 23838 35026
rect 26114 34974 26126 35026
rect 26178 34974 26190 35026
rect 28130 34974 28142 35026
rect 28194 34974 28206 35026
rect 32386 34974 32398 35026
rect 32450 34974 32462 35026
rect 34178 34974 34190 35026
rect 34242 34974 34254 35026
rect 35970 34974 35982 35026
rect 36034 34974 36046 35026
rect 39890 34974 39902 35026
rect 39954 34974 39966 35026
rect 41794 34974 41806 35026
rect 41858 34974 41870 35026
rect 43474 34974 43486 35026
rect 43538 34974 43550 35026
rect 50866 34974 50878 35026
rect 50930 34974 50942 35026
rect 54226 34974 54238 35026
rect 54290 34974 54302 35026
rect 57698 34974 57710 35026
rect 57762 34974 57774 35026
rect 59490 34974 59502 35026
rect 59554 34974 59566 35026
rect 62962 34974 62974 35026
rect 63026 34974 63038 35026
rect 70354 34974 70366 35026
rect 70418 34974 70430 35026
rect 72258 34974 72270 35026
rect 72322 34974 72334 35026
rect 74498 34974 74510 35026
rect 74562 34974 74574 35026
rect 80770 34974 80782 35026
rect 80834 34974 80846 35026
rect 82562 34974 82574 35026
rect 82626 34974 82638 35026
rect 85922 34974 85934 35026
rect 85986 34974 85998 35026
rect 87938 34974 87950 35026
rect 88002 34974 88014 35026
rect 93314 34974 93326 35026
rect 93378 34974 93390 35026
rect 95778 34974 95790 35026
rect 95842 34974 95854 35026
rect 97570 34974 97582 35026
rect 97634 34974 97646 35026
rect 99250 34974 99262 35026
rect 99314 34974 99326 35026
rect 101826 34974 101838 35026
rect 101890 34974 101902 35026
rect 103618 34974 103630 35026
rect 103682 34974 103694 35026
rect 109778 34974 109790 35026
rect 109842 34974 109854 35026
rect 111570 34974 111582 35026
rect 111634 34974 111646 35026
rect 115490 34974 115502 35026
rect 115554 34974 115566 35026
rect 118402 34974 118414 35026
rect 118466 34974 118478 35026
rect 12910 34962 12962 34974
rect 38446 34962 38498 34974
rect 88958 34962 89010 34974
rect 100270 34962 100322 34974
rect 121550 34962 121602 34974
rect 124014 35026 124066 35038
rect 140142 35026 140194 35038
rect 142830 35026 142882 35038
rect 125122 34974 125134 35026
rect 125186 34974 125198 35026
rect 127698 34974 127710 35026
rect 127762 34974 127774 35026
rect 133634 34974 133646 35026
rect 133698 34974 133710 35026
rect 136322 34974 136334 35026
rect 136386 34974 136398 35026
rect 141698 34974 141710 35026
rect 141762 34974 141774 35026
rect 124014 34962 124066 34974
rect 140142 34962 140194 34974
rect 142830 34962 142882 34974
rect 143278 35026 143330 35038
rect 143714 34974 143726 35026
rect 143778 34974 143790 35026
rect 143278 34962 143330 34974
rect 19742 34914 19794 34926
rect 45614 34914 45666 34926
rect 6738 34862 6750 34914
rect 6802 34862 6814 34914
rect 7522 34862 7534 34914
rect 7586 34862 7598 34914
rect 11218 34862 11230 34914
rect 11282 34862 11294 34914
rect 15026 34862 15038 34914
rect 15090 34862 15102 34914
rect 18274 34862 18286 34914
rect 18338 34862 18350 34914
rect 19058 34862 19070 34914
rect 19122 34862 19134 34914
rect 22866 34862 22878 34914
rect 22930 34862 22942 34914
rect 24882 34862 24894 34914
rect 24946 34862 24958 34914
rect 27010 34862 27022 34914
rect 27074 34862 27086 34914
rect 28802 34862 28814 34914
rect 28866 34862 28878 34914
rect 30818 34862 30830 34914
rect 30882 34862 30894 34914
rect 33170 34862 33182 34914
rect 33234 34862 33246 34914
rect 34962 34862 34974 34914
rect 35026 34862 35038 34914
rect 36754 34862 36766 34914
rect 36818 34862 36830 34914
rect 41010 34862 41022 34914
rect 41074 34862 41086 34914
rect 42802 34862 42814 34914
rect 42866 34862 42878 34914
rect 44594 34862 44606 34914
rect 44658 34862 44670 34914
rect 19742 34850 19794 34862
rect 45614 34850 45666 34862
rect 46398 34914 46450 34926
rect 46398 34850 46450 34862
rect 47854 34914 47906 34926
rect 61742 34914 61794 34926
rect 65550 34914 65602 34926
rect 76190 34914 76242 34926
rect 89966 34914 90018 34926
rect 104862 34914 104914 34926
rect 51986 34862 51998 34914
rect 52050 34862 52062 34914
rect 55346 34862 55358 34914
rect 55410 34862 55422 34914
rect 58706 34862 58718 34914
rect 58770 34862 58782 34914
rect 60610 34862 60622 34914
rect 60674 34862 60686 34914
rect 62178 34862 62190 34914
rect 62242 34862 62254 34914
rect 64082 34862 64094 34914
rect 64146 34862 64158 34914
rect 64866 34862 64878 34914
rect 64930 34862 64942 34914
rect 71474 34862 71486 34914
rect 71538 34862 71550 34914
rect 73266 34862 73278 34914
rect 73330 34862 73342 34914
rect 73826 34862 73838 34914
rect 73890 34862 73902 34914
rect 75730 34862 75742 34914
rect 75794 34862 75806 34914
rect 77410 34862 77422 34914
rect 77474 34862 77486 34914
rect 80098 34862 80110 34914
rect 80162 34862 80174 34914
rect 82002 34862 82014 34914
rect 82066 34862 82078 34914
rect 85250 34862 85262 34914
rect 85314 34862 85326 34914
rect 87266 34862 87278 34914
rect 87330 34862 87342 34914
rect 90402 34862 90414 34914
rect 90466 34862 90478 34914
rect 94210 34862 94222 34914
rect 94274 34862 94286 34914
rect 95106 34862 95118 34914
rect 95170 34862 95182 34914
rect 96786 34862 96798 34914
rect 96850 34862 96862 34914
rect 98578 34862 98590 34914
rect 98642 34862 98654 34914
rect 101154 34862 101166 34914
rect 101218 34862 101230 34914
rect 102946 34862 102958 34914
rect 103010 34862 103022 34914
rect 47854 34850 47906 34862
rect 61742 34850 61794 34862
rect 65550 34850 65602 34862
rect 76190 34850 76242 34862
rect 89966 34850 90018 34862
rect 104862 34850 104914 34862
rect 105422 34914 105474 34926
rect 105422 34850 105474 34862
rect 106878 34914 106930 34926
rect 113822 34914 113874 34926
rect 128830 34914 128882 34926
rect 109218 34862 109230 34914
rect 109282 34862 109294 34914
rect 110898 34862 110910 34914
rect 110962 34862 110974 34914
rect 114818 34862 114830 34914
rect 114882 34862 114894 34914
rect 117730 34862 117742 34914
rect 117794 34862 117806 34914
rect 119970 34862 119982 34914
rect 120034 34862 120046 34914
rect 122658 34862 122670 34914
rect 122722 34862 122734 34914
rect 126018 34862 126030 34914
rect 126082 34862 126094 34914
rect 126802 34862 126814 34914
rect 126866 34862 126878 34914
rect 130050 34862 130062 34914
rect 130114 34862 130126 34914
rect 132962 34862 132974 34914
rect 133026 34862 133038 34914
rect 135650 34862 135662 34914
rect 135714 34862 135726 34914
rect 141138 34862 141150 34914
rect 141202 34862 141214 34914
rect 106878 34850 106930 34862
rect 113822 34850 113874 34862
rect 128830 34850 128882 34862
rect 9326 34802 9378 34814
rect 9326 34738 9378 34750
rect 9662 34802 9714 34814
rect 9662 34738 9714 34750
rect 16158 34802 16210 34814
rect 52558 34802 52610 34814
rect 18946 34750 18958 34802
rect 19010 34750 19022 34802
rect 30594 34750 30606 34802
rect 30658 34750 30670 34802
rect 37650 34750 37662 34802
rect 37714 34750 37726 34802
rect 38210 34750 38222 34802
rect 38274 34750 38286 34802
rect 47058 34750 47070 34802
rect 47122 34750 47134 34802
rect 47506 34750 47518 34802
rect 47570 34750 47582 34802
rect 48962 34750 48974 34802
rect 49026 34750 49038 34802
rect 49522 34750 49534 34802
rect 49586 34750 49598 34802
rect 16158 34738 16210 34750
rect 52558 34738 52610 34750
rect 56702 34802 56754 34814
rect 56702 34738 56754 34750
rect 57038 34802 57090 34814
rect 78206 34802 78258 34814
rect 64754 34750 64766 34802
rect 64818 34750 64830 34802
rect 67330 34750 67342 34802
rect 67394 34750 67406 34802
rect 67890 34750 67902 34802
rect 67954 34750 67966 34802
rect 57038 34738 57090 34750
rect 78206 34738 78258 34750
rect 78542 34802 78594 34814
rect 78542 34738 78594 34750
rect 79438 34802 79490 34814
rect 79438 34738 79490 34750
rect 84030 34802 84082 34814
rect 84030 34738 84082 34750
rect 84366 34802 84418 34814
rect 92094 34802 92146 34814
rect 107886 34802 107938 34814
rect 131742 34802 131794 34814
rect 90514 34750 90526 34802
rect 90578 34750 90590 34802
rect 106082 34750 106094 34802
rect 106146 34750 106158 34802
rect 106642 34750 106654 34802
rect 106706 34750 106718 34802
rect 113138 34750 113150 34802
rect 113202 34750 113214 34802
rect 113474 34750 113486 34802
rect 113538 34750 113550 34802
rect 119858 34750 119870 34802
rect 119922 34750 119934 34802
rect 122322 34750 122334 34802
rect 122386 34750 122398 34802
rect 129938 34750 129950 34802
rect 130002 34750 130014 34802
rect 84366 34738 84418 34750
rect 92094 34738 92146 34750
rect 107886 34738 107938 34750
rect 131742 34738 131794 34750
rect 132078 34802 132130 34814
rect 132078 34738 132130 34750
rect 134766 34802 134818 34814
rect 139694 34802 139746 34814
rect 138002 34750 138014 34802
rect 138066 34750 138078 34802
rect 138562 34750 138574 34802
rect 138626 34750 138638 34802
rect 144722 34750 144734 34802
rect 144786 34750 144798 34802
rect 134766 34738 134818 34750
rect 139694 34738 139746 34750
rect 15598 34690 15650 34702
rect 15598 34626 15650 34638
rect 16494 34690 16546 34702
rect 16494 34626 16546 34638
rect 20078 34690 20130 34702
rect 20078 34626 20130 34638
rect 20750 34690 20802 34702
rect 20750 34626 20802 34638
rect 29710 34690 29762 34702
rect 29710 34626 29762 34638
rect 31502 34690 31554 34702
rect 31502 34626 31554 34638
rect 38782 34690 38834 34702
rect 38782 34626 38834 34638
rect 46062 34690 46114 34702
rect 46062 34626 46114 34638
rect 48190 34690 48242 34702
rect 48190 34626 48242 34638
rect 50094 34690 50146 34702
rect 50094 34626 50146 34638
rect 53678 34690 53730 34702
rect 53678 34626 53730 34638
rect 56254 34690 56306 34702
rect 56254 34626 56306 34638
rect 65886 34690 65938 34702
rect 65886 34626 65938 34638
rect 66782 34690 66834 34702
rect 66782 34626 66834 34638
rect 68462 34690 68514 34702
rect 68462 34626 68514 34638
rect 69470 34690 69522 34702
rect 69470 34626 69522 34638
rect 77646 34690 77698 34702
rect 77646 34626 77698 34638
rect 78990 34690 79042 34702
rect 78990 34626 79042 34638
rect 89630 34690 89682 34702
rect 89630 34626 89682 34638
rect 91310 34690 91362 34702
rect 91310 34626 91362 34638
rect 92430 34690 92482 34702
rect 92430 34626 92482 34638
rect 107214 34690 107266 34702
rect 107214 34626 107266 34638
rect 108222 34690 108274 34702
rect 108222 34626 108274 34638
rect 114158 34690 114210 34702
rect 114158 34626 114210 34638
rect 116958 34690 117010 34702
rect 116958 34626 117010 34638
rect 120990 34690 121042 34702
rect 120990 34626 121042 34638
rect 123454 34690 123506 34702
rect 123454 34626 123506 34638
rect 129278 34690 129330 34702
rect 129278 34626 129330 34638
rect 131070 34690 131122 34702
rect 131070 34626 131122 34638
rect 135102 34690 135154 34702
rect 135102 34626 135154 34638
rect 137342 34690 137394 34702
rect 137342 34626 137394 34638
rect 139134 34690 139186 34702
rect 139134 34626 139186 34638
rect 145630 34690 145682 34702
rect 145630 34626 145682 34638
rect 1344 34522 148784 34556
rect 1344 34470 38034 34522
rect 38086 34470 38138 34522
rect 38190 34470 38242 34522
rect 38294 34470 74854 34522
rect 74906 34470 74958 34522
rect 75010 34470 75062 34522
rect 75114 34470 111674 34522
rect 111726 34470 111778 34522
rect 111830 34470 111882 34522
rect 111934 34470 148494 34522
rect 148546 34470 148598 34522
rect 148650 34470 148702 34522
rect 148754 34470 148784 34522
rect 1344 34436 148784 34470
rect 7758 34354 7810 34366
rect 7758 34290 7810 34302
rect 10894 34354 10946 34366
rect 10894 34290 10946 34302
rect 11678 34354 11730 34366
rect 11678 34290 11730 34302
rect 14254 34354 14306 34366
rect 14254 34290 14306 34302
rect 15934 34354 15986 34366
rect 15934 34290 15986 34302
rect 16718 34354 16770 34366
rect 16718 34290 16770 34302
rect 17838 34354 17890 34366
rect 17838 34290 17890 34302
rect 18286 34354 18338 34366
rect 18286 34290 18338 34302
rect 19182 34354 19234 34366
rect 19182 34290 19234 34302
rect 22766 34354 22818 34366
rect 22766 34290 22818 34302
rect 23662 34354 23714 34366
rect 23662 34290 23714 34302
rect 24446 34354 24498 34366
rect 24446 34290 24498 34302
rect 27358 34354 27410 34366
rect 27358 34290 27410 34302
rect 27918 34354 27970 34366
rect 27918 34290 27970 34302
rect 28366 34354 28418 34366
rect 28366 34290 28418 34302
rect 29374 34354 29426 34366
rect 29374 34290 29426 34302
rect 33518 34354 33570 34366
rect 33518 34290 33570 34302
rect 33966 34354 34018 34366
rect 33966 34290 34018 34302
rect 35646 34354 35698 34366
rect 35646 34290 35698 34302
rect 36654 34354 36706 34366
rect 36654 34290 36706 34302
rect 37102 34354 37154 34366
rect 37102 34290 37154 34302
rect 39902 34354 39954 34366
rect 39902 34290 39954 34302
rect 43150 34354 43202 34366
rect 43150 34290 43202 34302
rect 44270 34354 44322 34366
rect 44270 34290 44322 34302
rect 44718 34354 44770 34366
rect 44718 34290 44770 34302
rect 48750 34354 48802 34366
rect 48750 34290 48802 34302
rect 56366 34354 56418 34366
rect 56366 34290 56418 34302
rect 56814 34354 56866 34366
rect 56814 34290 56866 34302
rect 57486 34354 57538 34366
rect 57486 34290 57538 34302
rect 72718 34354 72770 34366
rect 72718 34290 72770 34302
rect 73726 34354 73778 34366
rect 73726 34290 73778 34302
rect 74174 34354 74226 34366
rect 74174 34290 74226 34302
rect 74734 34354 74786 34366
rect 74734 34290 74786 34302
rect 75630 34354 75682 34366
rect 75630 34290 75682 34302
rect 76302 34354 76354 34366
rect 76302 34290 76354 34302
rect 78654 34354 78706 34366
rect 78654 34290 78706 34302
rect 85486 34354 85538 34366
rect 85486 34290 85538 34302
rect 87614 34354 87666 34366
rect 87614 34290 87666 34302
rect 93774 34354 93826 34366
rect 93774 34290 93826 34302
rect 95566 34354 95618 34366
rect 95566 34290 95618 34302
rect 96462 34354 96514 34366
rect 96462 34290 96514 34302
rect 98926 34354 98978 34366
rect 98926 34290 98978 34302
rect 101502 34354 101554 34366
rect 101502 34290 101554 34302
rect 102062 34354 102114 34366
rect 102062 34290 102114 34302
rect 109230 34354 109282 34366
rect 109230 34290 109282 34302
rect 109566 34354 109618 34366
rect 109566 34290 109618 34302
rect 110126 34354 110178 34366
rect 110126 34290 110178 34302
rect 110910 34354 110962 34366
rect 110910 34290 110962 34302
rect 111358 34354 111410 34366
rect 111358 34290 111410 34302
rect 115054 34354 115106 34366
rect 115054 34290 115106 34302
rect 117742 34354 117794 34366
rect 117742 34290 117794 34302
rect 125246 34354 125298 34366
rect 125246 34290 125298 34302
rect 125694 34354 125746 34366
rect 125694 34290 125746 34302
rect 126254 34354 126306 34366
rect 126254 34290 126306 34302
rect 129390 34354 129442 34366
rect 129390 34290 129442 34302
rect 132638 34354 132690 34366
rect 132638 34290 132690 34302
rect 133870 34354 133922 34366
rect 133870 34290 133922 34302
rect 134318 34354 134370 34366
rect 134318 34290 134370 34302
rect 134766 34354 134818 34366
rect 134766 34290 134818 34302
rect 135326 34354 135378 34366
rect 135326 34290 135378 34302
rect 136334 34354 136386 34366
rect 136334 34290 136386 34302
rect 11230 34242 11282 34254
rect 11230 34178 11282 34190
rect 16270 34242 16322 34254
rect 16270 34178 16322 34190
rect 18622 34242 18674 34254
rect 18622 34178 18674 34190
rect 21870 34242 21922 34254
rect 21870 34178 21922 34190
rect 22206 34242 22258 34254
rect 22206 34178 22258 34190
rect 23214 34242 23266 34254
rect 23214 34178 23266 34190
rect 26126 34242 26178 34254
rect 40462 34242 40514 34254
rect 29922 34190 29934 34242
rect 29986 34190 29998 34242
rect 31714 34190 31726 34242
rect 31778 34190 31790 34242
rect 38098 34190 38110 34242
rect 38162 34190 38174 34242
rect 26126 34178 26178 34190
rect 40462 34178 40514 34190
rect 40798 34242 40850 34254
rect 40798 34178 40850 34190
rect 42478 34242 42530 34254
rect 51438 34242 51490 34254
rect 54126 34242 54178 34254
rect 45266 34190 45278 34242
rect 45330 34190 45342 34242
rect 47058 34190 47070 34242
rect 47122 34190 47134 34242
rect 49634 34190 49646 34242
rect 49698 34190 49710 34242
rect 52434 34190 52446 34242
rect 52498 34190 52510 34242
rect 42478 34178 42530 34190
rect 51438 34178 51490 34190
rect 54126 34178 54178 34190
rect 58942 34242 58994 34254
rect 58942 34178 58994 34190
rect 60734 34242 60786 34254
rect 63646 34242 63698 34254
rect 61394 34190 61406 34242
rect 61458 34190 61470 34242
rect 60734 34178 60786 34190
rect 63646 34178 63698 34190
rect 64542 34242 64594 34254
rect 76862 34242 76914 34254
rect 68114 34190 68126 34242
rect 68178 34190 68190 34242
rect 68562 34190 68574 34242
rect 68626 34190 68638 34242
rect 69906 34190 69918 34242
rect 69970 34190 69982 34242
rect 64542 34178 64594 34190
rect 76862 34178 76914 34190
rect 77198 34242 77250 34254
rect 77198 34178 77250 34190
rect 88622 34242 88674 34254
rect 88622 34178 88674 34190
rect 89294 34242 89346 34254
rect 102622 34242 102674 34254
rect 137006 34242 137058 34254
rect 90402 34190 90414 34242
rect 90466 34190 90478 34242
rect 113362 34190 113374 34242
rect 113426 34190 113438 34242
rect 113810 34190 113822 34242
rect 113874 34190 113886 34242
rect 121426 34190 121438 34242
rect 121490 34190 121502 34242
rect 130610 34190 130622 34242
rect 130674 34190 130686 34242
rect 138338 34190 138350 34242
rect 138402 34190 138414 34242
rect 143042 34190 143054 34242
rect 143106 34190 143118 34242
rect 89294 34178 89346 34190
rect 102622 34178 102674 34190
rect 137006 34178 137058 34190
rect 8094 34130 8146 34142
rect 8094 34066 8146 34078
rect 14590 34130 14642 34142
rect 25790 34130 25842 34142
rect 37438 34130 37490 34142
rect 42142 34130 42194 34142
rect 51774 34130 51826 34142
rect 54462 34130 54514 34142
rect 19394 34078 19406 34130
rect 19458 34078 19470 34130
rect 20178 34078 20190 34130
rect 20242 34078 20254 34130
rect 31042 34078 31054 34130
rect 31106 34078 31118 34130
rect 32834 34078 32846 34130
rect 32898 34078 32910 34130
rect 39106 34078 39118 34130
rect 39170 34078 39182 34130
rect 46274 34078 46286 34130
rect 46338 34078 46350 34130
rect 48178 34078 48190 34130
rect 48242 34078 48254 34130
rect 50754 34078 50766 34130
rect 50818 34078 50830 34130
rect 53554 34078 53566 34130
rect 53618 34078 53630 34130
rect 14590 34066 14642 34078
rect 25790 34066 25842 34078
rect 37438 34066 37490 34078
rect 42142 34066 42194 34078
rect 51774 34066 51826 34078
rect 54462 34066 54514 34078
rect 57822 34130 57874 34142
rect 57822 34066 57874 34078
rect 58606 34130 58658 34142
rect 58606 34066 58658 34078
rect 60398 34130 60450 34142
rect 63310 34130 63362 34142
rect 68798 34130 68850 34142
rect 83806 34130 83858 34142
rect 62514 34078 62526 34130
rect 62578 34078 62590 34130
rect 64306 34078 64318 34130
rect 64370 34078 64382 34130
rect 67330 34078 67342 34130
rect 67394 34078 67406 34130
rect 71026 34078 71038 34130
rect 71090 34078 71102 34130
rect 73490 34078 73502 34130
rect 73554 34078 73566 34130
rect 81890 34078 81902 34130
rect 81954 34078 81966 34130
rect 60398 34066 60450 34078
rect 63310 34066 63362 34078
rect 68798 34066 68850 34078
rect 83806 34066 83858 34078
rect 89630 34130 89682 34142
rect 110462 34130 110514 34142
rect 90290 34078 90302 34130
rect 90354 34078 90366 34130
rect 92194 34078 92206 34130
rect 92258 34078 92270 34130
rect 97234 34078 97246 34130
rect 97298 34078 97310 34130
rect 100034 34078 100046 34130
rect 100098 34078 100110 34130
rect 103170 34078 103182 34130
rect 103234 34078 103246 34130
rect 105186 34078 105198 34130
rect 105250 34078 105262 34130
rect 106978 34078 106990 34130
rect 107042 34078 107054 34130
rect 89630 34066 89682 34078
rect 110462 34066 110514 34078
rect 111918 34130 111970 34142
rect 111918 34066 111970 34078
rect 114158 34130 114210 34142
rect 118078 34130 118130 34142
rect 131294 34130 131346 34142
rect 115938 34078 115950 34130
rect 116002 34078 116014 34130
rect 120082 34078 120094 34130
rect 120146 34078 120158 34130
rect 122546 34078 122558 34130
rect 122610 34078 122622 34130
rect 123106 34078 123118 34130
rect 123170 34078 123182 34130
rect 130498 34078 130510 34130
rect 130562 34078 130574 34130
rect 114158 34066 114210 34078
rect 118078 34066 118130 34078
rect 131294 34066 131346 34078
rect 132302 34130 132354 34142
rect 132302 34066 132354 34078
rect 133534 34130 133586 34142
rect 139022 34130 139074 34142
rect 143726 34130 143778 34142
rect 138562 34078 138574 34130
rect 138626 34078 138638 34130
rect 140018 34078 140030 34130
rect 140082 34078 140094 34130
rect 142930 34078 142942 34130
rect 142994 34078 143006 34130
rect 145058 34078 145070 34130
rect 145122 34078 145134 34130
rect 133534 34066 133586 34078
rect 139022 34066 139074 34078
rect 143726 34066 143778 34078
rect 7198 34018 7250 34030
rect 7198 33954 7250 33966
rect 8542 34018 8594 34030
rect 8542 33954 8594 33966
rect 9886 34018 9938 34030
rect 9886 33954 9938 33966
rect 15038 34018 15090 34030
rect 24894 34018 24946 34030
rect 20738 33966 20750 34018
rect 20802 33966 20814 34018
rect 15038 33954 15090 33966
rect 24894 33954 24946 33966
rect 28814 34018 28866 34030
rect 34526 34018 34578 34030
rect 31042 33966 31054 34018
rect 31106 34015 31118 34018
rect 31378 34015 31390 34018
rect 31106 33969 31390 34015
rect 31106 33966 31118 33969
rect 31378 33966 31390 33969
rect 31442 33966 31454 34018
rect 28814 33954 28866 33966
rect 34526 33954 34578 33966
rect 35198 34018 35250 34030
rect 35198 33954 35250 33966
rect 36094 34018 36146 34030
rect 36094 33954 36146 33966
rect 41582 34018 41634 34030
rect 41582 33954 41634 33966
rect 54910 34018 54962 34030
rect 54910 33954 54962 33966
rect 59502 34018 59554 34030
rect 59502 33954 59554 33966
rect 59838 34018 59890 34030
rect 59838 33954 59890 33966
rect 65662 34018 65714 34030
rect 71486 34018 71538 34030
rect 66434 33966 66446 34018
rect 66498 33966 66510 34018
rect 71026 33966 71038 34018
rect 71090 34015 71102 34018
rect 71090 33969 71311 34015
rect 71090 33966 71102 33969
rect 65662 33954 65714 33966
rect 69134 33906 69186 33918
rect 71265 33903 71311 33969
rect 71486 33954 71538 33966
rect 71934 34018 71986 34030
rect 71934 33954 71986 33966
rect 75070 34018 75122 34030
rect 75070 33954 75122 33966
rect 77646 34018 77698 34030
rect 77646 33954 77698 33966
rect 78206 34018 78258 34030
rect 78206 33954 78258 33966
rect 79102 34018 79154 34030
rect 79102 33954 79154 33966
rect 79774 34018 79826 34030
rect 79774 33954 79826 33966
rect 80558 34018 80610 34030
rect 80558 33954 80610 33966
rect 81454 34018 81506 34030
rect 84590 34018 84642 34030
rect 82674 33966 82686 34018
rect 82738 33966 82750 34018
rect 81454 33954 81506 33966
rect 84590 33954 84642 33966
rect 85150 34018 85202 34030
rect 85150 33954 85202 33966
rect 87054 34018 87106 34030
rect 87054 33954 87106 33966
rect 88174 34018 88226 34030
rect 88174 33954 88226 33966
rect 91086 34018 91138 34030
rect 94222 34018 94274 34030
rect 92754 33966 92766 34018
rect 92818 33966 92830 34018
rect 91086 33954 91138 33966
rect 94222 33954 94274 33966
rect 94782 34018 94834 34030
rect 94782 33954 94834 33966
rect 95118 34018 95170 34030
rect 95118 33954 95170 33966
rect 96014 34018 96066 34030
rect 108670 34018 108722 34030
rect 97906 33966 97918 34018
rect 97970 33966 97982 34018
rect 100482 33966 100494 34018
rect 100546 33966 100558 34018
rect 103842 33966 103854 34018
rect 103906 33966 103918 34018
rect 105858 33966 105870 34018
rect 105922 33966 105934 34018
rect 107650 33966 107662 34018
rect 107714 33966 107726 34018
rect 96014 33954 96066 33966
rect 108670 33954 108722 33966
rect 112478 34018 112530 34030
rect 118526 34018 118578 34030
rect 124798 34018 124850 34030
rect 116610 33966 116622 34018
rect 116674 33966 116686 34018
rect 119298 33966 119310 34018
rect 119362 33966 119374 34018
rect 123778 33966 123790 34018
rect 123842 33966 123854 34018
rect 112478 33954 112530 33966
rect 118526 33954 118578 33966
rect 124798 33954 124850 33966
rect 126590 34018 126642 34030
rect 126590 33954 126642 33966
rect 128942 34018 128994 34030
rect 128942 33954 128994 33966
rect 129950 34018 130002 34030
rect 129950 33954 130002 33966
rect 137342 34018 137394 34030
rect 141822 34018 141874 34030
rect 140690 33966 140702 34018
rect 140754 33966 140766 34018
rect 137342 33954 137394 33966
rect 141822 33954 141874 33966
rect 142382 34018 142434 34030
rect 145618 33966 145630 34018
rect 145682 33966 145694 34018
rect 142382 33954 142434 33966
rect 91422 33906 91474 33918
rect 114494 33906 114546 33918
rect 71474 33903 71486 33906
rect 71265 33857 71486 33903
rect 71474 33854 71486 33857
rect 71538 33854 71550 33906
rect 78194 33854 78206 33906
rect 78258 33903 78270 33906
rect 78754 33903 78766 33906
rect 78258 33857 78766 33903
rect 78258 33854 78270 33857
rect 78754 33854 78766 33857
rect 78818 33854 78830 33906
rect 96002 33854 96014 33906
rect 96066 33903 96078 33906
rect 96674 33903 96686 33906
rect 96066 33857 96686 33903
rect 96066 33854 96078 33857
rect 96674 33854 96686 33857
rect 96738 33854 96750 33906
rect 69134 33842 69186 33854
rect 91422 33842 91474 33854
rect 114494 33842 114546 33854
rect 131630 33906 131682 33918
rect 131630 33842 131682 33854
rect 139358 33906 139410 33918
rect 139358 33842 139410 33854
rect 144062 33906 144114 33918
rect 144062 33842 144114 33854
rect 1344 33738 148624 33772
rect 1344 33686 19624 33738
rect 19676 33686 19728 33738
rect 19780 33686 19832 33738
rect 19884 33686 56444 33738
rect 56496 33686 56548 33738
rect 56600 33686 56652 33738
rect 56704 33686 93264 33738
rect 93316 33686 93368 33738
rect 93420 33686 93472 33738
rect 93524 33686 130084 33738
rect 130136 33686 130188 33738
rect 130240 33686 130292 33738
rect 130344 33686 148624 33738
rect 1344 33652 148624 33686
rect 45490 33518 45502 33570
rect 45554 33567 45566 33570
rect 46162 33567 46174 33570
rect 45554 33521 46174 33567
rect 45554 33518 45566 33521
rect 46162 33518 46174 33521
rect 46226 33518 46238 33570
rect 69234 33518 69246 33570
rect 69298 33567 69310 33570
rect 69794 33567 69806 33570
rect 69298 33521 69806 33567
rect 69298 33518 69310 33521
rect 69794 33518 69806 33521
rect 69858 33518 69870 33570
rect 104850 33518 104862 33570
rect 104914 33567 104926 33570
rect 105410 33567 105422 33570
rect 104914 33521 105422 33567
rect 104914 33518 104926 33521
rect 105410 33518 105422 33521
rect 105474 33518 105486 33570
rect 121762 33518 121774 33570
rect 121826 33567 121838 33570
rect 122210 33567 122222 33570
rect 121826 33521 122222 33567
rect 121826 33518 121838 33521
rect 122210 33518 122222 33521
rect 122274 33518 122286 33570
rect 14926 33458 14978 33470
rect 14926 33394 14978 33406
rect 18846 33458 18898 33470
rect 18846 33394 18898 33406
rect 19742 33458 19794 33470
rect 19742 33394 19794 33406
rect 21534 33458 21586 33470
rect 21534 33394 21586 33406
rect 25230 33458 25282 33470
rect 25230 33394 25282 33406
rect 29486 33458 29538 33470
rect 29486 33394 29538 33406
rect 31838 33458 31890 33470
rect 31838 33394 31890 33406
rect 32622 33458 32674 33470
rect 32622 33394 32674 33406
rect 33406 33458 33458 33470
rect 33406 33394 33458 33406
rect 36878 33458 36930 33470
rect 36878 33394 36930 33406
rect 41806 33458 41858 33470
rect 41806 33394 41858 33406
rect 42142 33458 42194 33470
rect 42142 33394 42194 33406
rect 42702 33458 42754 33470
rect 42702 33394 42754 33406
rect 45502 33458 45554 33470
rect 45502 33394 45554 33406
rect 47518 33458 47570 33470
rect 47518 33394 47570 33406
rect 50766 33458 50818 33470
rect 50766 33394 50818 33406
rect 52446 33458 52498 33470
rect 52446 33394 52498 33406
rect 53454 33458 53506 33470
rect 53454 33394 53506 33406
rect 53902 33458 53954 33470
rect 53902 33394 53954 33406
rect 57150 33458 57202 33470
rect 57150 33394 57202 33406
rect 58270 33458 58322 33470
rect 58270 33394 58322 33406
rect 59166 33458 59218 33470
rect 59166 33394 59218 33406
rect 59614 33458 59666 33470
rect 59614 33394 59666 33406
rect 60174 33458 60226 33470
rect 60174 33394 60226 33406
rect 60734 33458 60786 33470
rect 67118 33458 67170 33470
rect 64978 33406 64990 33458
rect 65042 33406 65054 33458
rect 60734 33394 60786 33406
rect 67118 33394 67170 33406
rect 67678 33458 67730 33470
rect 67678 33394 67730 33406
rect 68126 33458 68178 33470
rect 68126 33394 68178 33406
rect 69358 33458 69410 33470
rect 69358 33394 69410 33406
rect 69806 33458 69858 33470
rect 69806 33394 69858 33406
rect 71374 33458 71426 33470
rect 71374 33394 71426 33406
rect 73726 33458 73778 33470
rect 73726 33394 73778 33406
rect 76078 33458 76130 33470
rect 76078 33394 76130 33406
rect 76526 33458 76578 33470
rect 76526 33394 76578 33406
rect 77982 33458 78034 33470
rect 77982 33394 78034 33406
rect 82574 33458 82626 33470
rect 91870 33458 91922 33470
rect 89058 33406 89070 33458
rect 89122 33406 89134 33458
rect 90738 33406 90750 33458
rect 90802 33406 90814 33458
rect 82574 33394 82626 33406
rect 91870 33394 91922 33406
rect 93214 33458 93266 33470
rect 93214 33394 93266 33406
rect 94110 33458 94162 33470
rect 94110 33394 94162 33406
rect 95230 33458 95282 33470
rect 95230 33394 95282 33406
rect 98254 33458 98306 33470
rect 98254 33394 98306 33406
rect 98590 33458 98642 33470
rect 98590 33394 98642 33406
rect 101054 33458 101106 33470
rect 101054 33394 101106 33406
rect 101614 33458 101666 33470
rect 101614 33394 101666 33406
rect 102734 33458 102786 33470
rect 102734 33394 102786 33406
rect 104078 33458 104130 33470
rect 104078 33394 104130 33406
rect 104974 33458 105026 33470
rect 104974 33394 105026 33406
rect 105422 33458 105474 33470
rect 105422 33394 105474 33406
rect 105870 33458 105922 33470
rect 105870 33394 105922 33406
rect 106318 33458 106370 33470
rect 106318 33394 106370 33406
rect 107662 33458 107714 33470
rect 107662 33394 107714 33406
rect 107998 33458 108050 33470
rect 107998 33394 108050 33406
rect 111918 33458 111970 33470
rect 114606 33458 114658 33470
rect 113026 33406 113038 33458
rect 113090 33406 113102 33458
rect 111918 33394 111970 33406
rect 114606 33394 114658 33406
rect 117070 33458 117122 33470
rect 117070 33394 117122 33406
rect 120654 33458 120706 33470
rect 120654 33394 120706 33406
rect 121102 33458 121154 33470
rect 121102 33394 121154 33406
rect 122894 33458 122946 33470
rect 133198 33458 133250 33470
rect 128594 33406 128606 33458
rect 128658 33406 128670 33458
rect 130498 33406 130510 33458
rect 130562 33406 130574 33458
rect 122894 33394 122946 33406
rect 133198 33394 133250 33406
rect 136782 33458 136834 33470
rect 139582 33458 139634 33470
rect 138114 33406 138126 33458
rect 138178 33406 138190 33458
rect 136782 33394 136834 33406
rect 139582 33394 139634 33406
rect 140142 33458 140194 33470
rect 140142 33394 140194 33406
rect 142718 33458 142770 33470
rect 142718 33394 142770 33406
rect 45950 33346 46002 33358
rect 45950 33282 46002 33294
rect 50206 33346 50258 33358
rect 50206 33282 50258 33294
rect 61518 33346 61570 33358
rect 61518 33282 61570 33294
rect 62078 33346 62130 33358
rect 62078 33282 62130 33294
rect 62638 33346 62690 33358
rect 106766 33346 106818 33358
rect 131966 33346 132018 33358
rect 65874 33294 65886 33346
rect 65938 33294 65950 33346
rect 88162 33294 88174 33346
rect 88226 33294 88238 33346
rect 89954 33294 89966 33346
rect 90018 33294 90030 33346
rect 112354 33294 112366 33346
rect 112418 33294 112430 33346
rect 129602 33294 129614 33346
rect 129666 33294 129678 33346
rect 131394 33294 131406 33346
rect 131458 33294 131470 33346
rect 137442 33294 137454 33346
rect 137506 33294 137518 33346
rect 62638 33282 62690 33294
rect 106766 33282 106818 33294
rect 131966 33282 132018 33294
rect 19406 33234 19458 33246
rect 19406 33170 19458 33182
rect 38670 33234 38722 33246
rect 38670 33170 38722 33182
rect 39902 33234 39954 33246
rect 39902 33170 39954 33182
rect 40462 33234 40514 33246
rect 40462 33170 40514 33182
rect 46398 33234 46450 33246
rect 46398 33170 46450 33182
rect 46734 33234 46786 33246
rect 46734 33170 46786 33182
rect 47966 33234 48018 33246
rect 47966 33170 48018 33182
rect 48302 33234 48354 33246
rect 48302 33170 48354 33182
rect 48862 33234 48914 33246
rect 48862 33170 48914 33182
rect 49198 33234 49250 33246
rect 49198 33170 49250 33182
rect 51214 33234 51266 33246
rect 51214 33170 51266 33182
rect 51550 33234 51602 33246
rect 99822 33234 99874 33246
rect 62962 33182 62974 33234
rect 63026 33182 63038 33234
rect 51550 33170 51602 33182
rect 99822 33170 99874 33182
rect 100270 33234 100322 33246
rect 100270 33170 100322 33182
rect 118414 33234 118466 33246
rect 118414 33170 118466 33182
rect 118750 33234 118802 33246
rect 118750 33170 118802 33182
rect 119646 33234 119698 33246
rect 119646 33170 119698 33182
rect 123902 33234 123954 33246
rect 123902 33170 123954 33182
rect 20526 33122 20578 33134
rect 20526 33058 20578 33070
rect 22094 33122 22146 33134
rect 22094 33058 22146 33070
rect 30830 33122 30882 33134
rect 30830 33058 30882 33070
rect 31390 33122 31442 33134
rect 31390 33058 31442 33070
rect 32286 33122 32338 33134
rect 32286 33058 32338 33070
rect 37662 33122 37714 33134
rect 37662 33058 37714 33070
rect 38110 33122 38162 33134
rect 38110 33058 38162 33070
rect 39006 33122 39058 33134
rect 39006 33058 39058 33070
rect 39566 33122 39618 33134
rect 39566 33058 39618 33070
rect 40798 33122 40850 33134
rect 40798 33058 40850 33070
rect 41246 33122 41298 33134
rect 41246 33058 41298 33070
rect 49870 33122 49922 33134
rect 49870 33058 49922 33070
rect 51998 33122 52050 33134
rect 51998 33058 52050 33070
rect 57822 33122 57874 33134
rect 57822 33058 57874 33070
rect 63422 33122 63474 33134
rect 63422 33058 63474 33070
rect 63870 33122 63922 33134
rect 63870 33058 63922 33070
rect 64318 33122 64370 33134
rect 64318 33058 64370 33070
rect 66670 33122 66722 33134
rect 66670 33058 66722 33070
rect 70814 33122 70866 33134
rect 70814 33058 70866 33070
rect 87726 33122 87778 33134
rect 87726 33058 87778 33070
rect 92206 33122 92258 33134
rect 92206 33058 92258 33070
rect 93550 33122 93602 33134
rect 93550 33058 93602 33070
rect 94782 33122 94834 33134
rect 94782 33058 94834 33070
rect 97246 33122 97298 33134
rect 97246 33058 97298 33070
rect 99486 33122 99538 33134
rect 99486 33058 99538 33070
rect 114046 33122 114098 33134
rect 114046 33058 114098 33070
rect 117406 33122 117458 33134
rect 117406 33058 117458 33070
rect 117854 33122 117906 33134
rect 117854 33058 117906 33070
rect 119310 33122 119362 33134
rect 119310 33058 119362 33070
rect 120094 33122 120146 33134
rect 120094 33058 120146 33070
rect 121774 33122 121826 33134
rect 121774 33058 121826 33070
rect 122110 33122 122162 33134
rect 122110 33058 122162 33070
rect 123566 33122 123618 33134
rect 123566 33058 123618 33070
rect 124910 33122 124962 33134
rect 124910 33058 124962 33070
rect 1344 32954 148784 32988
rect 1344 32902 38034 32954
rect 38086 32902 38138 32954
rect 38190 32902 38242 32954
rect 38294 32902 74854 32954
rect 74906 32902 74958 32954
rect 75010 32902 75062 32954
rect 75114 32902 111674 32954
rect 111726 32902 111778 32954
rect 111830 32902 111882 32954
rect 111934 32902 148494 32954
rect 148546 32902 148598 32954
rect 148650 32902 148702 32954
rect 148754 32902 148784 32954
rect 1344 32868 148784 32902
rect 39454 32786 39506 32798
rect 39454 32722 39506 32734
rect 40126 32786 40178 32798
rect 40126 32722 40178 32734
rect 41582 32786 41634 32798
rect 41582 32722 41634 32734
rect 42030 32786 42082 32798
rect 42030 32722 42082 32734
rect 46510 32786 46562 32798
rect 46510 32722 46562 32734
rect 46958 32786 47010 32798
rect 46958 32722 47010 32734
rect 47630 32786 47682 32798
rect 47630 32722 47682 32734
rect 48190 32786 48242 32798
rect 48190 32722 48242 32734
rect 49422 32786 49474 32798
rect 49422 32722 49474 32734
rect 49870 32786 49922 32798
rect 49870 32722 49922 32734
rect 50542 32786 50594 32798
rect 50542 32722 50594 32734
rect 62302 32786 62354 32798
rect 62302 32722 62354 32734
rect 62862 32786 62914 32798
rect 62862 32722 62914 32734
rect 63198 32786 63250 32798
rect 63198 32722 63250 32734
rect 63982 32786 64034 32798
rect 63982 32722 64034 32734
rect 65438 32786 65490 32798
rect 65438 32722 65490 32734
rect 65774 32786 65826 32798
rect 65774 32722 65826 32734
rect 66222 32786 66274 32798
rect 66222 32722 66274 32734
rect 67118 32786 67170 32798
rect 67118 32722 67170 32734
rect 89294 32786 89346 32798
rect 89294 32722 89346 32734
rect 90750 32786 90802 32798
rect 90750 32722 90802 32734
rect 91198 32786 91250 32798
rect 91198 32722 91250 32734
rect 92430 32786 92482 32798
rect 92430 32722 92482 32734
rect 119758 32786 119810 32798
rect 119758 32722 119810 32734
rect 130958 32786 131010 32798
rect 130958 32722 131010 32734
rect 131406 32786 131458 32798
rect 131406 32722 131458 32734
rect 38446 32674 38498 32686
rect 38446 32610 38498 32622
rect 91646 32674 91698 32686
rect 91646 32610 91698 32622
rect 39006 32562 39058 32574
rect 39006 32498 39058 32510
rect 40798 32562 40850 32574
rect 40798 32498 40850 32510
rect 48526 32562 48578 32574
rect 48526 32498 48578 32510
rect 91982 32562 92034 32574
rect 91982 32498 92034 32510
rect 51326 32450 51378 32462
rect 51326 32386 51378 32398
rect 52558 32450 52610 32462
rect 52558 32386 52610 32398
rect 61854 32450 61906 32462
rect 61854 32386 61906 32398
rect 64430 32450 64482 32462
rect 64430 32386 64482 32398
rect 89742 32450 89794 32462
rect 89742 32386 89794 32398
rect 92990 32450 93042 32462
rect 92990 32386 93042 32398
rect 118750 32450 118802 32462
rect 118750 32386 118802 32398
rect 119310 32450 119362 32462
rect 119310 32386 119362 32398
rect 1344 32170 148624 32204
rect 1344 32118 19624 32170
rect 19676 32118 19728 32170
rect 19780 32118 19832 32170
rect 19884 32118 56444 32170
rect 56496 32118 56548 32170
rect 56600 32118 56652 32170
rect 56704 32118 93264 32170
rect 93316 32118 93368 32170
rect 93420 32118 93472 32170
rect 93524 32118 130084 32170
rect 130136 32118 130188 32170
rect 130240 32118 130292 32170
rect 130344 32118 148624 32170
rect 1344 32084 148624 32118
rect 64878 31890 64930 31902
rect 64878 31826 64930 31838
rect 48974 31554 49026 31566
rect 48974 31490 49026 31502
rect 1344 31386 148784 31420
rect 1344 31334 38034 31386
rect 38086 31334 38138 31386
rect 38190 31334 38242 31386
rect 38294 31334 74854 31386
rect 74906 31334 74958 31386
rect 75010 31334 75062 31386
rect 75114 31334 111674 31386
rect 111726 31334 111778 31386
rect 111830 31334 111882 31386
rect 111934 31334 148494 31386
rect 148546 31334 148598 31386
rect 148650 31334 148702 31386
rect 148754 31334 148784 31386
rect 1344 31300 148784 31334
rect 1344 30602 148624 30636
rect 1344 30550 19624 30602
rect 19676 30550 19728 30602
rect 19780 30550 19832 30602
rect 19884 30550 56444 30602
rect 56496 30550 56548 30602
rect 56600 30550 56652 30602
rect 56704 30550 93264 30602
rect 93316 30550 93368 30602
rect 93420 30550 93472 30602
rect 93524 30550 130084 30602
rect 130136 30550 130188 30602
rect 130240 30550 130292 30602
rect 130344 30550 148624 30602
rect 1344 30516 148624 30550
rect 1344 29818 148784 29852
rect 1344 29766 38034 29818
rect 38086 29766 38138 29818
rect 38190 29766 38242 29818
rect 38294 29766 74854 29818
rect 74906 29766 74958 29818
rect 75010 29766 75062 29818
rect 75114 29766 111674 29818
rect 111726 29766 111778 29818
rect 111830 29766 111882 29818
rect 111934 29766 148494 29818
rect 148546 29766 148598 29818
rect 148650 29766 148702 29818
rect 148754 29766 148784 29818
rect 1344 29732 148784 29766
rect 1344 29034 148624 29068
rect 1344 28982 19624 29034
rect 19676 28982 19728 29034
rect 19780 28982 19832 29034
rect 19884 28982 56444 29034
rect 56496 28982 56548 29034
rect 56600 28982 56652 29034
rect 56704 28982 93264 29034
rect 93316 28982 93368 29034
rect 93420 28982 93472 29034
rect 93524 28982 130084 29034
rect 130136 28982 130188 29034
rect 130240 28982 130292 29034
rect 130344 28982 148624 29034
rect 1344 28948 148624 28982
rect 1344 28250 148784 28284
rect 1344 28198 38034 28250
rect 38086 28198 38138 28250
rect 38190 28198 38242 28250
rect 38294 28198 74854 28250
rect 74906 28198 74958 28250
rect 75010 28198 75062 28250
rect 75114 28198 111674 28250
rect 111726 28198 111778 28250
rect 111830 28198 111882 28250
rect 111934 28198 148494 28250
rect 148546 28198 148598 28250
rect 148650 28198 148702 28250
rect 148754 28198 148784 28250
rect 1344 28164 148784 28198
rect 1344 27466 148624 27500
rect 1344 27414 19624 27466
rect 19676 27414 19728 27466
rect 19780 27414 19832 27466
rect 19884 27414 56444 27466
rect 56496 27414 56548 27466
rect 56600 27414 56652 27466
rect 56704 27414 93264 27466
rect 93316 27414 93368 27466
rect 93420 27414 93472 27466
rect 93524 27414 130084 27466
rect 130136 27414 130188 27466
rect 130240 27414 130292 27466
rect 130344 27414 148624 27466
rect 1344 27380 148624 27414
rect 1344 26682 148784 26716
rect 1344 26630 38034 26682
rect 38086 26630 38138 26682
rect 38190 26630 38242 26682
rect 38294 26630 74854 26682
rect 74906 26630 74958 26682
rect 75010 26630 75062 26682
rect 75114 26630 111674 26682
rect 111726 26630 111778 26682
rect 111830 26630 111882 26682
rect 111934 26630 148494 26682
rect 148546 26630 148598 26682
rect 148650 26630 148702 26682
rect 148754 26630 148784 26682
rect 1344 26596 148784 26630
rect 1344 25898 148624 25932
rect 1344 25846 19624 25898
rect 19676 25846 19728 25898
rect 19780 25846 19832 25898
rect 19884 25846 56444 25898
rect 56496 25846 56548 25898
rect 56600 25846 56652 25898
rect 56704 25846 93264 25898
rect 93316 25846 93368 25898
rect 93420 25846 93472 25898
rect 93524 25846 130084 25898
rect 130136 25846 130188 25898
rect 130240 25846 130292 25898
rect 130344 25846 148624 25898
rect 1344 25812 148624 25846
rect 1344 25114 148784 25148
rect 1344 25062 38034 25114
rect 38086 25062 38138 25114
rect 38190 25062 38242 25114
rect 38294 25062 74854 25114
rect 74906 25062 74958 25114
rect 75010 25062 75062 25114
rect 75114 25062 111674 25114
rect 111726 25062 111778 25114
rect 111830 25062 111882 25114
rect 111934 25062 148494 25114
rect 148546 25062 148598 25114
rect 148650 25062 148702 25114
rect 148754 25062 148784 25114
rect 1344 25028 148784 25062
rect 1344 24330 148624 24364
rect 1344 24278 19624 24330
rect 19676 24278 19728 24330
rect 19780 24278 19832 24330
rect 19884 24278 56444 24330
rect 56496 24278 56548 24330
rect 56600 24278 56652 24330
rect 56704 24278 93264 24330
rect 93316 24278 93368 24330
rect 93420 24278 93472 24330
rect 93524 24278 130084 24330
rect 130136 24278 130188 24330
rect 130240 24278 130292 24330
rect 130344 24278 148624 24330
rect 1344 24244 148624 24278
rect 1344 23546 148784 23580
rect 1344 23494 38034 23546
rect 38086 23494 38138 23546
rect 38190 23494 38242 23546
rect 38294 23494 74854 23546
rect 74906 23494 74958 23546
rect 75010 23494 75062 23546
rect 75114 23494 111674 23546
rect 111726 23494 111778 23546
rect 111830 23494 111882 23546
rect 111934 23494 148494 23546
rect 148546 23494 148598 23546
rect 148650 23494 148702 23546
rect 148754 23494 148784 23546
rect 1344 23460 148784 23494
rect 1344 22762 148624 22796
rect 1344 22710 19624 22762
rect 19676 22710 19728 22762
rect 19780 22710 19832 22762
rect 19884 22710 56444 22762
rect 56496 22710 56548 22762
rect 56600 22710 56652 22762
rect 56704 22710 93264 22762
rect 93316 22710 93368 22762
rect 93420 22710 93472 22762
rect 93524 22710 130084 22762
rect 130136 22710 130188 22762
rect 130240 22710 130292 22762
rect 130344 22710 148624 22762
rect 1344 22676 148624 22710
rect 1344 21978 148784 22012
rect 1344 21926 38034 21978
rect 38086 21926 38138 21978
rect 38190 21926 38242 21978
rect 38294 21926 74854 21978
rect 74906 21926 74958 21978
rect 75010 21926 75062 21978
rect 75114 21926 111674 21978
rect 111726 21926 111778 21978
rect 111830 21926 111882 21978
rect 111934 21926 148494 21978
rect 148546 21926 148598 21978
rect 148650 21926 148702 21978
rect 148754 21926 148784 21978
rect 1344 21892 148784 21926
rect 1344 21194 148624 21228
rect 1344 21142 19624 21194
rect 19676 21142 19728 21194
rect 19780 21142 19832 21194
rect 19884 21142 56444 21194
rect 56496 21142 56548 21194
rect 56600 21142 56652 21194
rect 56704 21142 93264 21194
rect 93316 21142 93368 21194
rect 93420 21142 93472 21194
rect 93524 21142 130084 21194
rect 130136 21142 130188 21194
rect 130240 21142 130292 21194
rect 130344 21142 148624 21194
rect 1344 21108 148624 21142
rect 1344 20410 148784 20444
rect 1344 20358 38034 20410
rect 38086 20358 38138 20410
rect 38190 20358 38242 20410
rect 38294 20358 74854 20410
rect 74906 20358 74958 20410
rect 75010 20358 75062 20410
rect 75114 20358 111674 20410
rect 111726 20358 111778 20410
rect 111830 20358 111882 20410
rect 111934 20358 148494 20410
rect 148546 20358 148598 20410
rect 148650 20358 148702 20410
rect 148754 20358 148784 20410
rect 1344 20324 148784 20358
rect 1344 19626 148624 19660
rect 1344 19574 19624 19626
rect 19676 19574 19728 19626
rect 19780 19574 19832 19626
rect 19884 19574 56444 19626
rect 56496 19574 56548 19626
rect 56600 19574 56652 19626
rect 56704 19574 93264 19626
rect 93316 19574 93368 19626
rect 93420 19574 93472 19626
rect 93524 19574 130084 19626
rect 130136 19574 130188 19626
rect 130240 19574 130292 19626
rect 130344 19574 148624 19626
rect 1344 19540 148624 19574
rect 1344 18842 148784 18876
rect 1344 18790 38034 18842
rect 38086 18790 38138 18842
rect 38190 18790 38242 18842
rect 38294 18790 74854 18842
rect 74906 18790 74958 18842
rect 75010 18790 75062 18842
rect 75114 18790 111674 18842
rect 111726 18790 111778 18842
rect 111830 18790 111882 18842
rect 111934 18790 148494 18842
rect 148546 18790 148598 18842
rect 148650 18790 148702 18842
rect 148754 18790 148784 18842
rect 1344 18756 148784 18790
rect 1344 18058 148624 18092
rect 1344 18006 19624 18058
rect 19676 18006 19728 18058
rect 19780 18006 19832 18058
rect 19884 18006 56444 18058
rect 56496 18006 56548 18058
rect 56600 18006 56652 18058
rect 56704 18006 93264 18058
rect 93316 18006 93368 18058
rect 93420 18006 93472 18058
rect 93524 18006 130084 18058
rect 130136 18006 130188 18058
rect 130240 18006 130292 18058
rect 130344 18006 148624 18058
rect 1344 17972 148624 18006
rect 1344 17274 148784 17308
rect 1344 17222 38034 17274
rect 38086 17222 38138 17274
rect 38190 17222 38242 17274
rect 38294 17222 74854 17274
rect 74906 17222 74958 17274
rect 75010 17222 75062 17274
rect 75114 17222 111674 17274
rect 111726 17222 111778 17274
rect 111830 17222 111882 17274
rect 111934 17222 148494 17274
rect 148546 17222 148598 17274
rect 148650 17222 148702 17274
rect 148754 17222 148784 17274
rect 1344 17188 148784 17222
rect 1344 16490 148624 16524
rect 1344 16438 19624 16490
rect 19676 16438 19728 16490
rect 19780 16438 19832 16490
rect 19884 16438 56444 16490
rect 56496 16438 56548 16490
rect 56600 16438 56652 16490
rect 56704 16438 93264 16490
rect 93316 16438 93368 16490
rect 93420 16438 93472 16490
rect 93524 16438 130084 16490
rect 130136 16438 130188 16490
rect 130240 16438 130292 16490
rect 130344 16438 148624 16490
rect 1344 16404 148624 16438
rect 1344 15706 148784 15740
rect 1344 15654 38034 15706
rect 38086 15654 38138 15706
rect 38190 15654 38242 15706
rect 38294 15654 74854 15706
rect 74906 15654 74958 15706
rect 75010 15654 75062 15706
rect 75114 15654 111674 15706
rect 111726 15654 111778 15706
rect 111830 15654 111882 15706
rect 111934 15654 148494 15706
rect 148546 15654 148598 15706
rect 148650 15654 148702 15706
rect 148754 15654 148784 15706
rect 1344 15620 148784 15654
rect 1344 14922 148624 14956
rect 1344 14870 19624 14922
rect 19676 14870 19728 14922
rect 19780 14870 19832 14922
rect 19884 14870 56444 14922
rect 56496 14870 56548 14922
rect 56600 14870 56652 14922
rect 56704 14870 93264 14922
rect 93316 14870 93368 14922
rect 93420 14870 93472 14922
rect 93524 14870 130084 14922
rect 130136 14870 130188 14922
rect 130240 14870 130292 14922
rect 130344 14870 148624 14922
rect 1344 14836 148624 14870
rect 1344 14138 148784 14172
rect 1344 14086 38034 14138
rect 38086 14086 38138 14138
rect 38190 14086 38242 14138
rect 38294 14086 74854 14138
rect 74906 14086 74958 14138
rect 75010 14086 75062 14138
rect 75114 14086 111674 14138
rect 111726 14086 111778 14138
rect 111830 14086 111882 14138
rect 111934 14086 148494 14138
rect 148546 14086 148598 14138
rect 148650 14086 148702 14138
rect 148754 14086 148784 14138
rect 1344 14052 148784 14086
rect 1344 13354 148624 13388
rect 1344 13302 19624 13354
rect 19676 13302 19728 13354
rect 19780 13302 19832 13354
rect 19884 13302 56444 13354
rect 56496 13302 56548 13354
rect 56600 13302 56652 13354
rect 56704 13302 93264 13354
rect 93316 13302 93368 13354
rect 93420 13302 93472 13354
rect 93524 13302 130084 13354
rect 130136 13302 130188 13354
rect 130240 13302 130292 13354
rect 130344 13302 148624 13354
rect 1344 13268 148624 13302
rect 1344 12570 148784 12604
rect 1344 12518 38034 12570
rect 38086 12518 38138 12570
rect 38190 12518 38242 12570
rect 38294 12518 74854 12570
rect 74906 12518 74958 12570
rect 75010 12518 75062 12570
rect 75114 12518 111674 12570
rect 111726 12518 111778 12570
rect 111830 12518 111882 12570
rect 111934 12518 148494 12570
rect 148546 12518 148598 12570
rect 148650 12518 148702 12570
rect 148754 12518 148784 12570
rect 1344 12484 148784 12518
rect 1344 11786 148624 11820
rect 1344 11734 19624 11786
rect 19676 11734 19728 11786
rect 19780 11734 19832 11786
rect 19884 11734 56444 11786
rect 56496 11734 56548 11786
rect 56600 11734 56652 11786
rect 56704 11734 93264 11786
rect 93316 11734 93368 11786
rect 93420 11734 93472 11786
rect 93524 11734 130084 11786
rect 130136 11734 130188 11786
rect 130240 11734 130292 11786
rect 130344 11734 148624 11786
rect 1344 11700 148624 11734
rect 1344 11002 148784 11036
rect 1344 10950 38034 11002
rect 38086 10950 38138 11002
rect 38190 10950 38242 11002
rect 38294 10950 74854 11002
rect 74906 10950 74958 11002
rect 75010 10950 75062 11002
rect 75114 10950 111674 11002
rect 111726 10950 111778 11002
rect 111830 10950 111882 11002
rect 111934 10950 148494 11002
rect 148546 10950 148598 11002
rect 148650 10950 148702 11002
rect 148754 10950 148784 11002
rect 1344 10916 148784 10950
rect 1344 10218 148624 10252
rect 1344 10166 19624 10218
rect 19676 10166 19728 10218
rect 19780 10166 19832 10218
rect 19884 10166 56444 10218
rect 56496 10166 56548 10218
rect 56600 10166 56652 10218
rect 56704 10166 93264 10218
rect 93316 10166 93368 10218
rect 93420 10166 93472 10218
rect 93524 10166 130084 10218
rect 130136 10166 130188 10218
rect 130240 10166 130292 10218
rect 130344 10166 148624 10218
rect 1344 10132 148624 10166
rect 128718 9938 128770 9950
rect 128718 9874 128770 9886
rect 129278 9602 129330 9614
rect 129278 9538 129330 9550
rect 1344 9434 148784 9468
rect 1344 9382 38034 9434
rect 38086 9382 38138 9434
rect 38190 9382 38242 9434
rect 38294 9382 74854 9434
rect 74906 9382 74958 9434
rect 75010 9382 75062 9434
rect 75114 9382 111674 9434
rect 111726 9382 111778 9434
rect 111830 9382 111882 9434
rect 111934 9382 148494 9434
rect 148546 9382 148598 9434
rect 148650 9382 148702 9434
rect 148754 9382 148784 9434
rect 1344 9348 148784 9382
rect 67230 9266 67282 9278
rect 67230 9202 67282 9214
rect 64654 9154 64706 9166
rect 128270 9154 128322 9166
rect 131294 9154 131346 9166
rect 66098 9102 66110 9154
rect 66162 9102 66174 9154
rect 66434 9102 66446 9154
rect 66498 9102 66510 9154
rect 130162 9102 130174 9154
rect 130226 9102 130238 9154
rect 64654 9090 64706 9102
rect 128270 9090 128322 9102
rect 131294 9090 131346 9102
rect 65886 9042 65938 9054
rect 129166 9042 129218 9054
rect 128034 8990 128046 9042
rect 128098 8990 128110 9042
rect 65886 8978 65938 8990
rect 129166 8978 129218 8990
rect 129502 9042 129554 9054
rect 130846 9042 130898 9054
rect 130274 8990 130286 9042
rect 130338 8990 130350 9042
rect 129502 8978 129554 8990
rect 130846 8978 130898 8990
rect 64318 8930 64370 8942
rect 64318 8866 64370 8878
rect 65550 8818 65602 8830
rect 65550 8754 65602 8766
rect 1344 8650 148624 8684
rect 1344 8598 19624 8650
rect 19676 8598 19728 8650
rect 19780 8598 19832 8650
rect 19884 8598 56444 8650
rect 56496 8598 56548 8650
rect 56600 8598 56652 8650
rect 56704 8598 93264 8650
rect 93316 8598 93368 8650
rect 93420 8598 93472 8650
rect 93524 8598 130084 8650
rect 130136 8598 130188 8650
rect 130240 8598 130292 8650
rect 130344 8598 148624 8650
rect 1344 8564 148624 8598
rect 67678 8370 67730 8382
rect 67678 8306 67730 8318
rect 63646 8258 63698 8270
rect 119198 8258 119250 8270
rect 64194 8206 64206 8258
rect 64258 8206 64270 8258
rect 63646 8194 63698 8206
rect 119198 8194 119250 8206
rect 120542 8258 120594 8270
rect 131854 8258 131906 8270
rect 131282 8206 131294 8258
rect 131346 8206 131358 8258
rect 120542 8194 120594 8206
rect 131854 8194 131906 8206
rect 118302 8146 118354 8158
rect 127374 8146 127426 8158
rect 119410 8094 119422 8146
rect 119474 8094 119486 8146
rect 119858 8094 119870 8146
rect 119922 8094 119934 8146
rect 118302 8082 118354 8094
rect 127374 8082 127426 8094
rect 63198 8034 63250 8046
rect 67342 8034 67394 8046
rect 66770 7982 66782 8034
rect 66834 7982 66846 8034
rect 63198 7970 63250 7982
rect 67342 7970 67394 7982
rect 68238 8034 68290 8046
rect 68238 7970 68290 7982
rect 88958 8034 89010 8046
rect 88958 7970 89010 7982
rect 118862 8034 118914 8046
rect 118862 7970 118914 7982
rect 121102 8034 121154 8046
rect 121102 7970 121154 7982
rect 121438 8034 121490 8046
rect 121438 7970 121490 7982
rect 126814 8034 126866 8046
rect 126814 7970 126866 7982
rect 127710 8034 127762 8046
rect 127710 7970 127762 7982
rect 128158 8034 128210 8046
rect 132302 8034 132354 8046
rect 128930 7982 128942 8034
rect 128994 7982 129006 8034
rect 128158 7970 128210 7982
rect 132302 7970 132354 7982
rect 132862 8034 132914 8046
rect 132862 7970 132914 7982
rect 1344 7866 148784 7900
rect 1344 7814 38034 7866
rect 38086 7814 38138 7866
rect 38190 7814 38242 7866
rect 38294 7814 74854 7866
rect 74906 7814 74958 7866
rect 75010 7814 75062 7866
rect 75114 7814 111674 7866
rect 111726 7814 111778 7866
rect 111830 7814 111882 7866
rect 111934 7814 148494 7866
rect 148546 7814 148598 7866
rect 148650 7814 148702 7866
rect 148754 7814 148784 7866
rect 1344 7780 148784 7814
rect 19966 7698 20018 7710
rect 19966 7634 20018 7646
rect 78318 7698 78370 7710
rect 78318 7634 78370 7646
rect 90862 7698 90914 7710
rect 90862 7634 90914 7646
rect 113598 7698 113650 7710
rect 113598 7634 113650 7646
rect 123342 7698 123394 7710
rect 123342 7634 123394 7646
rect 126366 7698 126418 7710
rect 126366 7634 126418 7646
rect 127038 7698 127090 7710
rect 127038 7634 127090 7646
rect 28366 7586 28418 7598
rect 62526 7586 62578 7598
rect 19058 7534 19070 7586
rect 19122 7534 19134 7586
rect 50306 7534 50318 7586
rect 50370 7534 50382 7586
rect 28366 7522 28418 7534
rect 62526 7522 62578 7534
rect 62862 7586 62914 7598
rect 63534 7586 63586 7598
rect 67790 7586 67842 7598
rect 99598 7586 99650 7598
rect 63074 7534 63086 7586
rect 63138 7583 63150 7586
rect 63298 7583 63310 7586
rect 63138 7537 63310 7583
rect 63138 7534 63150 7537
rect 63298 7534 63310 7537
rect 63362 7534 63374 7586
rect 66098 7534 66110 7586
rect 66162 7534 66174 7586
rect 66434 7534 66446 7586
rect 66498 7534 66510 7586
rect 76290 7534 76302 7586
rect 76354 7534 76366 7586
rect 76738 7534 76750 7586
rect 76802 7534 76814 7586
rect 62862 7522 62914 7534
rect 63534 7522 63586 7534
rect 67790 7522 67842 7534
rect 99598 7522 99650 7534
rect 118078 7586 118130 7598
rect 126030 7586 126082 7598
rect 129726 7586 129778 7598
rect 119634 7534 119646 7586
rect 119698 7534 119710 7586
rect 120194 7534 120206 7586
rect 120258 7534 120270 7586
rect 121314 7534 121326 7586
rect 121378 7534 121390 7586
rect 128034 7534 128046 7586
rect 128098 7534 128110 7586
rect 118078 7522 118130 7534
rect 126030 7522 126082 7534
rect 129726 7522 129778 7534
rect 141486 7586 141538 7598
rect 141486 7522 141538 7534
rect 142382 7586 142434 7598
rect 142382 7522 142434 7534
rect 18510 7474 18562 7486
rect 28702 7474 28754 7486
rect 18946 7422 18958 7474
rect 19010 7422 19022 7474
rect 18510 7410 18562 7422
rect 28702 7410 28754 7422
rect 48750 7474 48802 7486
rect 51550 7474 51602 7486
rect 50530 7422 50542 7474
rect 50594 7422 50606 7474
rect 48750 7410 48802 7422
rect 51550 7410 51602 7422
rect 63870 7474 63922 7486
rect 63870 7410 63922 7422
rect 65550 7474 65602 7486
rect 65550 7410 65602 7422
rect 65886 7474 65938 7486
rect 65886 7410 65938 7422
rect 68126 7474 68178 7486
rect 68126 7410 68178 7422
rect 76974 7474 77026 7486
rect 76974 7410 77026 7422
rect 88510 7474 88562 7486
rect 88510 7410 88562 7422
rect 99262 7474 99314 7486
rect 99262 7410 99314 7422
rect 118414 7474 118466 7486
rect 118414 7410 118466 7422
rect 119086 7474 119138 7486
rect 119086 7410 119138 7422
rect 119422 7474 119474 7486
rect 121998 7474 122050 7486
rect 132638 7474 132690 7486
rect 121202 7422 121214 7474
rect 121266 7422 121278 7474
rect 128146 7422 128158 7474
rect 128210 7422 128222 7474
rect 132066 7422 132078 7474
rect 132130 7422 132142 7474
rect 119422 7410 119474 7422
rect 121998 7410 122050 7422
rect 132638 7410 132690 7422
rect 141822 7474 141874 7486
rect 142594 7422 142606 7474
rect 142658 7422 142670 7474
rect 141822 7410 141874 7422
rect 20302 7362 20354 7374
rect 20302 7298 20354 7310
rect 20750 7362 20802 7374
rect 20750 7298 20802 7310
rect 26350 7362 26402 7374
rect 26350 7298 26402 7310
rect 29150 7362 29202 7374
rect 29150 7298 29202 7310
rect 39230 7362 39282 7374
rect 39230 7298 39282 7310
rect 39790 7362 39842 7374
rect 39790 7298 39842 7310
rect 48414 7362 48466 7374
rect 48414 7298 48466 7310
rect 49758 7362 49810 7374
rect 49758 7298 49810 7310
rect 51102 7362 51154 7374
rect 51102 7298 51154 7310
rect 64654 7362 64706 7374
rect 64654 7298 64706 7310
rect 67230 7362 67282 7374
rect 67230 7298 67282 7310
rect 68686 7362 68738 7374
rect 68686 7298 68738 7310
rect 69134 7362 69186 7374
rect 69134 7298 69186 7310
rect 69470 7362 69522 7374
rect 69470 7298 69522 7310
rect 69918 7362 69970 7374
rect 69918 7298 69970 7310
rect 75070 7362 75122 7374
rect 75070 7298 75122 7310
rect 75518 7362 75570 7374
rect 75518 7298 75570 7310
rect 77870 7362 77922 7374
rect 77870 7298 77922 7310
rect 89182 7362 89234 7374
rect 89182 7298 89234 7310
rect 89630 7362 89682 7374
rect 89630 7298 89682 7310
rect 90414 7362 90466 7374
rect 90414 7298 90466 7310
rect 91422 7362 91474 7374
rect 91422 7298 91474 7310
rect 113038 7362 113090 7374
rect 113038 7298 113090 7310
rect 114158 7362 114210 7374
rect 114158 7298 114210 7310
rect 115950 7362 116002 7374
rect 115950 7298 116002 7310
rect 116734 7362 116786 7374
rect 116734 7298 116786 7310
rect 117518 7362 117570 7374
rect 117518 7298 117570 7310
rect 122894 7362 122946 7374
rect 122894 7298 122946 7310
rect 133086 7362 133138 7374
rect 133086 7298 133138 7310
rect 133534 7362 133586 7374
rect 133534 7298 133586 7310
rect 18174 7250 18226 7262
rect 18174 7186 18226 7198
rect 64542 7250 64594 7262
rect 64542 7186 64594 7198
rect 77310 7250 77362 7262
rect 122334 7250 122386 7262
rect 77634 7198 77646 7250
rect 77698 7247 77710 7250
rect 78194 7247 78206 7250
rect 77698 7201 78206 7247
rect 77698 7198 77710 7201
rect 78194 7198 78206 7201
rect 78258 7198 78270 7250
rect 113362 7198 113374 7250
rect 113426 7247 113438 7250
rect 114146 7247 114158 7250
rect 113426 7201 114158 7247
rect 113426 7198 113438 7201
rect 114146 7198 114158 7201
rect 114210 7198 114222 7250
rect 77310 7186 77362 7198
rect 122334 7186 122386 7198
rect 127374 7250 127426 7262
rect 127374 7186 127426 7198
rect 128942 7250 128994 7262
rect 128942 7186 128994 7198
rect 1344 7082 148624 7116
rect 1344 7030 19624 7082
rect 19676 7030 19728 7082
rect 19780 7030 19832 7082
rect 19884 7030 56444 7082
rect 56496 7030 56548 7082
rect 56600 7030 56652 7082
rect 56704 7030 93264 7082
rect 93316 7030 93368 7082
rect 93420 7030 93472 7082
rect 93524 7030 130084 7082
rect 130136 7030 130188 7082
rect 130240 7030 130292 7082
rect 130344 7030 148624 7082
rect 1344 6996 148624 7030
rect 27134 6914 27186 6926
rect 27134 6850 27186 6862
rect 29710 6914 29762 6926
rect 29710 6850 29762 6862
rect 30046 6914 30098 6926
rect 30046 6850 30098 6862
rect 47854 6914 47906 6926
rect 47854 6850 47906 6862
rect 50206 6914 50258 6926
rect 50206 6850 50258 6862
rect 68126 6914 68178 6926
rect 68126 6850 68178 6862
rect 68462 6914 68514 6926
rect 68462 6850 68514 6862
rect 87390 6914 87442 6926
rect 87390 6850 87442 6862
rect 89742 6914 89794 6926
rect 89742 6850 89794 6862
rect 91198 6914 91250 6926
rect 91198 6850 91250 6862
rect 99150 6914 99202 6926
rect 99150 6850 99202 6862
rect 99486 6914 99538 6926
rect 141822 6914 141874 6926
rect 126578 6862 126590 6914
rect 126642 6911 126654 6914
rect 127362 6911 127374 6914
rect 126642 6865 127374 6911
rect 126642 6862 126654 6865
rect 127362 6862 127374 6865
rect 127426 6862 127438 6914
rect 99486 6850 99538 6862
rect 141822 6850 141874 6862
rect 142158 6914 142210 6926
rect 142158 6850 142210 6862
rect 39118 6802 39170 6814
rect 39118 6738 39170 6750
rect 40126 6802 40178 6814
rect 40126 6738 40178 6750
rect 114382 6802 114434 6814
rect 114382 6738 114434 6750
rect 115726 6802 115778 6814
rect 115726 6738 115778 6750
rect 7422 6690 7474 6702
rect 16158 6690 16210 6702
rect 20862 6690 20914 6702
rect 31502 6690 31554 6702
rect 51214 6690 51266 6702
rect 78206 6690 78258 6702
rect 93102 6690 93154 6702
rect 7858 6638 7870 6690
rect 7922 6638 7934 6690
rect 16706 6638 16718 6690
rect 16770 6638 16782 6690
rect 20402 6638 20414 6690
rect 20466 6638 20478 6690
rect 27794 6638 27806 6690
rect 27858 6638 27870 6690
rect 49522 6638 49534 6690
rect 49586 6638 49598 6690
rect 62290 6638 62302 6690
rect 62354 6638 62366 6690
rect 62850 6638 62862 6690
rect 62914 6638 62926 6690
rect 71250 6638 71262 6690
rect 71314 6638 71326 6690
rect 81106 6638 81118 6690
rect 81170 6638 81182 6690
rect 89170 6638 89182 6690
rect 89234 6638 89246 6690
rect 91970 6638 91982 6690
rect 92034 6638 92046 6690
rect 7422 6626 7474 6638
rect 16158 6626 16210 6638
rect 20862 6626 20914 6638
rect 31502 6626 31554 6638
rect 51214 6626 51266 6638
rect 78206 6626 78258 6638
rect 93102 6626 93154 6638
rect 98478 6690 98530 6702
rect 101054 6690 101106 6702
rect 100258 6638 100270 6690
rect 100322 6638 100334 6690
rect 98478 6626 98530 6638
rect 101054 6626 101106 6638
rect 111582 6690 111634 6702
rect 117630 6690 117682 6702
rect 122110 6690 122162 6702
rect 113362 6638 113374 6690
rect 113426 6638 113438 6690
rect 115154 6638 115166 6690
rect 115218 6638 115230 6690
rect 118290 6638 118302 6690
rect 118354 6638 118366 6690
rect 111582 6626 111634 6638
rect 117630 6626 117682 6638
rect 122110 6626 122162 6638
rect 127038 6690 127090 6702
rect 127038 6626 127090 6638
rect 128046 6690 128098 6702
rect 133646 6690 133698 6702
rect 128370 6638 128382 6690
rect 128434 6638 128446 6690
rect 128046 6626 128098 6638
rect 133646 6626 133698 6638
rect 143950 6690 144002 6702
rect 143950 6626 144002 6638
rect 10894 6578 10946 6590
rect 10894 6514 10946 6526
rect 26126 6578 26178 6590
rect 26126 6514 26178 6526
rect 26798 6578 26850 6590
rect 28814 6578 28866 6590
rect 50542 6578 50594 6590
rect 27906 6526 27918 6578
rect 27970 6526 27982 6578
rect 30258 6526 30270 6578
rect 30322 6526 30334 6578
rect 30818 6526 30830 6578
rect 30882 6526 30894 6578
rect 38322 6526 38334 6578
rect 38386 6526 38398 6578
rect 38882 6526 38894 6578
rect 38946 6526 38958 6578
rect 48066 6526 48078 6578
rect 48130 6526 48142 6578
rect 48402 6526 48414 6578
rect 48466 6526 48478 6578
rect 49410 6526 49422 6578
rect 49474 6526 49486 6578
rect 26798 6514 26850 6526
rect 28814 6514 28866 6526
rect 50542 6514 50594 6526
rect 52110 6578 52162 6590
rect 52110 6514 52162 6526
rect 66334 6578 66386 6590
rect 66334 6514 66386 6526
rect 66670 6578 66722 6590
rect 69470 6578 69522 6590
rect 77646 6578 77698 6590
rect 81566 6578 81618 6590
rect 131966 6578 132018 6590
rect 67554 6526 67566 6578
rect 67618 6526 67630 6578
rect 67890 6526 67902 6578
rect 67954 6526 67966 6578
rect 73266 6526 73278 6578
rect 73330 6526 73342 6578
rect 79986 6526 79998 6578
rect 80050 6526 80062 6578
rect 87602 6526 87614 6578
rect 87666 6526 87678 6578
rect 88162 6526 88174 6578
rect 88226 6526 88238 6578
rect 89058 6526 89070 6578
rect 89122 6526 89134 6578
rect 91858 6526 91870 6578
rect 91922 6526 91934 6578
rect 100034 6526 100046 6578
rect 100098 6526 100110 6578
rect 112242 6526 112254 6578
rect 112306 6526 112318 6578
rect 115042 6526 115054 6578
rect 115106 6526 115118 6578
rect 66670 6514 66722 6526
rect 69470 6514 69522 6526
rect 77646 6514 77698 6526
rect 81566 6514 81618 6526
rect 131966 6514 132018 6526
rect 132078 6578 132130 6590
rect 132078 6514 132130 6526
rect 133086 6578 133138 6590
rect 133086 6514 133138 6526
rect 133758 6578 133810 6590
rect 142482 6526 142494 6578
rect 142546 6526 142558 6578
rect 142706 6526 142718 6578
rect 142770 6526 142782 6578
rect 133758 6514 133810 6526
rect 11230 6466 11282 6478
rect 19854 6466 19906 6478
rect 10322 6414 10334 6466
rect 10386 6414 10398 6466
rect 19170 6414 19182 6466
rect 19234 6414 19246 6466
rect 11230 6402 11282 6414
rect 19854 6402 19906 6414
rect 21534 6466 21586 6478
rect 21534 6402 21586 6414
rect 25790 6466 25842 6478
rect 25790 6402 25842 6414
rect 39454 6466 39506 6478
rect 39454 6402 39506 6414
rect 40462 6466 40514 6478
rect 40462 6402 40514 6414
rect 47518 6466 47570 6478
rect 47518 6402 47570 6414
rect 51550 6466 51602 6478
rect 51550 6402 51602 6414
rect 52446 6466 52498 6478
rect 52446 6402 52498 6414
rect 61854 6466 61906 6478
rect 65886 6466 65938 6478
rect 65314 6414 65326 6466
rect 65378 6414 65390 6466
rect 61854 6402 61906 6414
rect 65886 6402 65938 6414
rect 69358 6466 69410 6478
rect 69358 6402 69410 6414
rect 69918 6466 69970 6478
rect 69918 6402 69970 6414
rect 70702 6466 70754 6478
rect 70702 6402 70754 6414
rect 77310 6466 77362 6478
rect 77310 6402 77362 6414
rect 78542 6466 78594 6478
rect 78542 6402 78594 6414
rect 87054 6466 87106 6478
rect 87054 6402 87106 6414
rect 90078 6466 90130 6478
rect 90078 6402 90130 6414
rect 90862 6466 90914 6478
rect 90862 6402 90914 6414
rect 93662 6466 93714 6478
rect 93662 6402 93714 6414
rect 101614 6466 101666 6478
rect 101614 6402 101666 6414
rect 110462 6466 110514 6478
rect 110462 6402 110514 6414
rect 111022 6466 111074 6478
rect 111022 6402 111074 6414
rect 114046 6466 114098 6478
rect 114046 6402 114098 6414
rect 116286 6466 116338 6478
rect 116286 6402 116338 6414
rect 117182 6466 117234 6478
rect 121326 6466 121378 6478
rect 120530 6414 120542 6466
rect 120594 6414 120606 6466
rect 117182 6402 117234 6414
rect 121326 6402 121378 6414
rect 121774 6466 121826 6478
rect 121774 6402 121826 6414
rect 127374 6466 127426 6478
rect 131518 6466 131570 6478
rect 130946 6414 130958 6466
rect 131010 6414 131022 6466
rect 127374 6402 127426 6414
rect 131518 6402 131570 6414
rect 132974 6466 133026 6478
rect 132974 6402 133026 6414
rect 134206 6466 134258 6478
rect 134206 6402 134258 6414
rect 141262 6466 141314 6478
rect 141262 6402 141314 6414
rect 143502 6466 143554 6478
rect 143502 6402 143554 6414
rect 1344 6298 148784 6332
rect 1344 6246 38034 6298
rect 38086 6246 38138 6298
rect 38190 6246 38242 6298
rect 38294 6246 74854 6298
rect 74906 6246 74958 6298
rect 75010 6246 75062 6298
rect 75114 6246 111674 6298
rect 111726 6246 111778 6298
rect 111830 6246 111882 6298
rect 111934 6246 148494 6298
rect 148546 6246 148598 6298
rect 148650 6246 148702 6298
rect 148754 6246 148784 6298
rect 1344 6212 148784 6246
rect 8094 6130 8146 6142
rect 8094 6066 8146 6078
rect 11342 6130 11394 6142
rect 11342 6066 11394 6078
rect 14926 6130 14978 6142
rect 14926 6066 14978 6078
rect 16046 6130 16098 6142
rect 16046 6066 16098 6078
rect 17838 6130 17890 6142
rect 17838 6066 17890 6078
rect 20526 6130 20578 6142
rect 31502 6130 31554 6142
rect 30930 6078 30942 6130
rect 30994 6078 31006 6130
rect 20526 6066 20578 6078
rect 31502 6066 31554 6078
rect 50318 6130 50370 6142
rect 50318 6066 50370 6078
rect 51102 6130 51154 6142
rect 51102 6066 51154 6078
rect 59950 6130 60002 6142
rect 59950 6066 60002 6078
rect 60846 6130 60898 6142
rect 60846 6066 60898 6078
rect 65550 6130 65602 6142
rect 72158 6130 72210 6142
rect 70130 6078 70142 6130
rect 70194 6078 70206 6130
rect 65550 6066 65602 6078
rect 72158 6066 72210 6078
rect 73502 6130 73554 6142
rect 73502 6066 73554 6078
rect 74062 6130 74114 6142
rect 74062 6066 74114 6078
rect 75742 6130 75794 6142
rect 75742 6066 75794 6078
rect 87390 6130 87442 6142
rect 87390 6066 87442 6078
rect 88510 6130 88562 6142
rect 88510 6066 88562 6078
rect 90414 6130 90466 6142
rect 90414 6066 90466 6078
rect 101726 6130 101778 6142
rect 101726 6066 101778 6078
rect 107886 6130 107938 6142
rect 107886 6066 107938 6078
rect 110350 6130 110402 6142
rect 110350 6066 110402 6078
rect 113374 6130 113426 6142
rect 126478 6130 126530 6142
rect 140254 6130 140306 6142
rect 117058 6078 117070 6130
rect 117122 6078 117134 6130
rect 132066 6078 132078 6130
rect 132130 6078 132142 6130
rect 113374 6066 113426 6078
rect 126478 6066 126530 6078
rect 140254 6066 140306 6078
rect 143726 6130 143778 6142
rect 143726 6066 143778 6078
rect 145294 6130 145346 6142
rect 145294 6066 145346 6078
rect 16606 6018 16658 6030
rect 16606 5954 16658 5966
rect 16942 6018 16994 6030
rect 21982 6018 22034 6030
rect 39678 6018 39730 6030
rect 18946 5966 18958 6018
rect 19010 5966 19022 6018
rect 19506 5966 19518 6018
rect 19570 5966 19582 6018
rect 38434 5966 38446 6018
rect 38498 5966 38510 6018
rect 16942 5954 16994 5966
rect 21982 5954 22034 5966
rect 39678 5954 39730 5966
rect 46622 6018 46674 6030
rect 46622 5954 46674 5966
rect 46958 6018 47010 6030
rect 71150 6018 71202 6030
rect 77086 6018 77138 6030
rect 61506 5966 61518 6018
rect 61570 5966 61582 6018
rect 74722 5966 74734 6018
rect 74786 5966 74798 6018
rect 75170 5966 75182 6018
rect 75234 5966 75246 6018
rect 46958 5954 47010 5966
rect 71150 5954 71202 5966
rect 77086 5954 77138 5966
rect 86158 6018 86210 6030
rect 86158 5954 86210 5966
rect 86494 6018 86546 6030
rect 86494 5954 86546 5966
rect 89630 6018 89682 6030
rect 89630 5954 89682 5966
rect 91534 6018 91586 6030
rect 91534 5954 91586 5966
rect 91870 6018 91922 6030
rect 91870 5954 91922 5966
rect 108558 6018 108610 6030
rect 112030 6018 112082 6030
rect 109666 5966 109678 6018
rect 109730 5966 109742 6018
rect 108558 5954 108610 5966
rect 112030 5954 112082 5966
rect 112366 6018 112418 6030
rect 115614 6018 115666 6030
rect 115042 5966 115054 6018
rect 115106 5966 115118 6018
rect 112366 5954 112418 5966
rect 115614 5954 115666 5966
rect 133086 6018 133138 6030
rect 133086 5954 133138 5966
rect 134094 6018 134146 6030
rect 134094 5954 134146 5966
rect 137902 6018 137954 6030
rect 144846 6018 144898 6030
rect 138674 5966 138686 6018
rect 138738 5966 138750 6018
rect 139122 5966 139134 6018
rect 139186 5966 139198 6018
rect 142706 5966 142718 6018
rect 142770 5966 142782 6018
rect 137902 5954 137954 5966
rect 144846 5954 144898 5966
rect 8430 5906 8482 5918
rect 18398 5906 18450 5918
rect 15810 5854 15822 5906
rect 15874 5854 15886 5906
rect 8430 5842 8482 5854
rect 18398 5842 18450 5854
rect 18734 5906 18786 5918
rect 28030 5906 28082 5918
rect 31838 5906 31890 5918
rect 37886 5906 37938 5918
rect 41470 5906 41522 5918
rect 49758 5906 49810 5918
rect 53342 5906 53394 5918
rect 66110 5906 66162 5918
rect 26898 5854 26910 5906
rect 26962 5854 26974 5906
rect 28354 5854 28366 5906
rect 28418 5854 28430 5906
rect 36754 5854 36766 5906
rect 36818 5854 36830 5906
rect 38658 5854 38670 5906
rect 38722 5854 38734 5906
rect 39442 5854 39454 5906
rect 39506 5854 39518 5906
rect 48738 5854 48750 5906
rect 48802 5854 48814 5906
rect 52882 5854 52894 5906
rect 52946 5854 52958 5906
rect 64642 5854 64654 5906
rect 64706 5854 64718 5906
rect 18734 5842 18786 5854
rect 28030 5842 28082 5854
rect 31838 5842 31890 5854
rect 37886 5842 37938 5854
rect 41470 5842 41522 5854
rect 49758 5842 49810 5854
rect 53342 5842 53394 5854
rect 66110 5842 66162 5854
rect 67006 5906 67058 5918
rect 70702 5906 70754 5918
rect 67666 5854 67678 5906
rect 67730 5854 67742 5906
rect 67006 5842 67058 5854
rect 70702 5842 70754 5854
rect 75406 5906 75458 5918
rect 79998 5906 80050 5918
rect 79314 5854 79326 5906
rect 79378 5854 79390 5906
rect 75406 5842 75458 5854
rect 79998 5842 80050 5854
rect 87950 5906 88002 5918
rect 90974 5906 91026 5918
rect 108894 5906 108946 5918
rect 114270 5906 114322 5918
rect 116510 5906 116562 5918
rect 119982 5906 120034 5918
rect 129166 5906 129218 5918
rect 139358 5906 139410 5918
rect 89394 5854 89406 5906
rect 89458 5854 89470 5906
rect 101266 5854 101278 5906
rect 101330 5854 101342 5906
rect 109554 5854 109566 5906
rect 109618 5854 109630 5906
rect 114930 5854 114942 5906
rect 114994 5854 115006 5906
rect 119634 5854 119646 5906
rect 119698 5854 119710 5906
rect 127138 5854 127150 5906
rect 127202 5854 127214 5906
rect 129602 5854 129614 5906
rect 129666 5854 129678 5906
rect 133298 5854 133310 5906
rect 133362 5854 133374 5906
rect 87950 5842 88002 5854
rect 90974 5842 91026 5854
rect 108894 5842 108946 5854
rect 114270 5842 114322 5854
rect 116510 5842 116562 5854
rect 119982 5842 120034 5854
rect 129166 5842 129218 5854
rect 139358 5842 139410 5854
rect 140814 5906 140866 5918
rect 140814 5842 140866 5854
rect 141374 5906 141426 5918
rect 143390 5906 143442 5918
rect 142594 5854 142606 5906
rect 142658 5854 142670 5906
rect 141374 5842 141426 5854
rect 143390 5842 143442 5854
rect 9774 5794 9826 5806
rect 9774 5730 9826 5742
rect 10110 5794 10162 5806
rect 10110 5730 10162 5742
rect 11902 5794 11954 5806
rect 11902 5730 11954 5742
rect 12462 5794 12514 5806
rect 12462 5730 12514 5742
rect 20638 5794 20690 5806
rect 20638 5730 20690 5742
rect 21198 5794 21250 5806
rect 21198 5730 21250 5742
rect 21534 5794 21586 5806
rect 27470 5794 27522 5806
rect 40238 5794 40290 5806
rect 25778 5742 25790 5794
rect 25842 5742 25854 5794
rect 35634 5742 35646 5794
rect 35698 5742 35710 5794
rect 21534 5730 21586 5742
rect 27470 5730 27522 5742
rect 40238 5730 40290 5742
rect 40910 5794 40962 5806
rect 40910 5730 40962 5742
rect 45278 5794 45330 5806
rect 56478 5794 56530 5806
rect 47618 5742 47630 5794
rect 47682 5742 47694 5794
rect 51762 5742 51774 5794
rect 51826 5742 51838 5794
rect 45278 5730 45330 5742
rect 56478 5730 56530 5742
rect 57486 5794 57538 5806
rect 57486 5730 57538 5742
rect 60510 5794 60562 5806
rect 66670 5794 66722 5806
rect 62626 5742 62638 5794
rect 62690 5742 62702 5794
rect 63522 5742 63534 5794
rect 63586 5742 63598 5794
rect 60510 5730 60562 5742
rect 66670 5730 66722 5742
rect 71262 5794 71314 5806
rect 71262 5730 71314 5742
rect 71710 5794 71762 5806
rect 71710 5730 71762 5742
rect 72606 5794 72658 5806
rect 72606 5730 72658 5742
rect 80446 5794 80498 5806
rect 80446 5730 80498 5742
rect 92430 5794 92482 5806
rect 92430 5730 92482 5742
rect 94894 5794 94946 5806
rect 110686 5794 110738 5806
rect 100146 5742 100158 5794
rect 100210 5742 100222 5794
rect 94894 5730 94946 5742
rect 110686 5730 110738 5742
rect 111134 5794 111186 5806
rect 111134 5730 111186 5742
rect 116174 5794 116226 5806
rect 116174 5730 116226 5742
rect 120990 5794 121042 5806
rect 134542 5794 134594 5806
rect 128146 5742 128158 5794
rect 128210 5742 128222 5794
rect 120990 5730 121042 5742
rect 134542 5730 134594 5742
rect 134990 5794 135042 5806
rect 134990 5730 135042 5742
rect 135438 5794 135490 5806
rect 135438 5730 135490 5742
rect 137454 5794 137506 5806
rect 137454 5730 137506 5742
rect 141934 5794 141986 5806
rect 141934 5730 141986 5742
rect 37550 5682 37602 5694
rect 37550 5618 37602 5630
rect 40350 5682 40402 5694
rect 76302 5682 76354 5694
rect 60498 5630 60510 5682
rect 60562 5679 60574 5682
rect 61170 5679 61182 5682
rect 60562 5633 61182 5679
rect 60562 5630 60574 5633
rect 61170 5630 61182 5633
rect 61234 5630 61246 5682
rect 40350 5618 40402 5630
rect 76302 5618 76354 5630
rect 113934 5682 113986 5694
rect 113934 5618 113986 5630
rect 132638 5682 132690 5694
rect 132638 5618 132690 5630
rect 133982 5682 134034 5694
rect 133982 5618 134034 5630
rect 139694 5682 139746 5694
rect 139694 5618 139746 5630
rect 1344 5514 148624 5548
rect 1344 5462 19624 5514
rect 19676 5462 19728 5514
rect 19780 5462 19832 5514
rect 19884 5462 56444 5514
rect 56496 5462 56548 5514
rect 56600 5462 56652 5514
rect 56704 5462 93264 5514
rect 93316 5462 93368 5514
rect 93420 5462 93472 5514
rect 93524 5462 130084 5514
rect 130136 5462 130188 5514
rect 130240 5462 130292 5514
rect 130344 5462 148624 5514
rect 1344 5428 148624 5462
rect 20862 5346 20914 5358
rect 20862 5282 20914 5294
rect 28702 5346 28754 5358
rect 28702 5282 28754 5294
rect 31950 5346 32002 5358
rect 31950 5282 32002 5294
rect 37438 5346 37490 5358
rect 37438 5282 37490 5294
rect 49086 5346 49138 5358
rect 49086 5282 49138 5294
rect 67342 5346 67394 5358
rect 67342 5282 67394 5294
rect 67678 5346 67730 5358
rect 67678 5282 67730 5294
rect 72942 5346 72994 5358
rect 72942 5282 72994 5294
rect 88958 5346 89010 5358
rect 88958 5282 89010 5294
rect 98702 5346 98754 5358
rect 98702 5282 98754 5294
rect 115502 5346 115554 5358
rect 115502 5282 115554 5294
rect 116286 5346 116338 5358
rect 116286 5282 116338 5294
rect 131518 5346 131570 5358
rect 131518 5282 131570 5294
rect 132862 5346 132914 5358
rect 132862 5282 132914 5294
rect 138350 5346 138402 5358
rect 138350 5282 138402 5294
rect 12686 5234 12738 5246
rect 12686 5170 12738 5182
rect 21758 5234 21810 5246
rect 21758 5170 21810 5182
rect 22206 5234 22258 5246
rect 41694 5234 41746 5246
rect 53566 5234 53618 5246
rect 35410 5182 35422 5234
rect 35474 5182 35486 5234
rect 46946 5182 46958 5234
rect 47010 5182 47022 5234
rect 22206 5170 22258 5182
rect 41694 5170 41746 5182
rect 53566 5170 53618 5182
rect 54126 5234 54178 5246
rect 54126 5170 54178 5182
rect 54462 5234 54514 5246
rect 89406 5234 89458 5246
rect 59602 5182 59614 5234
rect 59666 5182 59678 5234
rect 62178 5182 62190 5234
rect 62242 5182 62254 5234
rect 54462 5170 54514 5182
rect 89406 5170 89458 5182
rect 90078 5234 90130 5246
rect 90078 5170 90130 5182
rect 91646 5234 91698 5246
rect 91646 5170 91698 5182
rect 92206 5234 92258 5246
rect 92206 5170 92258 5182
rect 93102 5234 93154 5246
rect 93102 5170 93154 5182
rect 101950 5234 102002 5246
rect 101950 5170 102002 5182
rect 102510 5234 102562 5246
rect 102510 5170 102562 5182
rect 105758 5234 105810 5246
rect 105758 5170 105810 5182
rect 116174 5234 116226 5246
rect 116174 5170 116226 5182
rect 120990 5234 121042 5246
rect 126926 5234 126978 5246
rect 125682 5182 125694 5234
rect 125746 5182 125758 5234
rect 120990 5170 121042 5182
rect 126926 5170 126978 5182
rect 132078 5234 132130 5246
rect 132078 5170 132130 5182
rect 138014 5234 138066 5246
rect 138014 5170 138066 5182
rect 139694 5234 139746 5246
rect 139694 5170 139746 5182
rect 140142 5234 140194 5246
rect 140142 5170 140194 5182
rect 140814 5234 140866 5246
rect 140814 5170 140866 5182
rect 141374 5234 141426 5246
rect 144510 5234 144562 5246
rect 142706 5182 142718 5234
rect 142770 5182 142782 5234
rect 141374 5170 141426 5182
rect 144510 5170 144562 5182
rect 145854 5234 145906 5246
rect 145854 5170 145906 5182
rect 146526 5234 146578 5246
rect 146526 5170 146578 5182
rect 11678 5122 11730 5134
rect 15822 5122 15874 5134
rect 7410 5070 7422 5122
rect 7474 5070 7486 5122
rect 7858 5070 7870 5122
rect 7922 5070 7934 5122
rect 10210 5070 10222 5122
rect 10274 5070 10286 5122
rect 15138 5070 15150 5122
rect 15202 5070 15214 5122
rect 11678 5058 11730 5070
rect 15822 5058 15874 5070
rect 16494 5122 16546 5134
rect 16494 5058 16546 5070
rect 17166 5122 17218 5134
rect 29486 5122 29538 5134
rect 17714 5070 17726 5122
rect 17778 5070 17790 5122
rect 25106 5070 25118 5122
rect 25170 5070 25182 5122
rect 25666 5070 25678 5122
rect 25730 5070 25742 5122
rect 17166 5058 17218 5070
rect 29486 5058 29538 5070
rect 30270 5122 30322 5134
rect 32062 5122 32114 5134
rect 31378 5070 31390 5122
rect 31442 5070 31454 5122
rect 30270 5058 30322 5070
rect 32062 5058 32114 5070
rect 32510 5122 32562 5134
rect 41582 5122 41634 5134
rect 40450 5070 40462 5122
rect 40514 5070 40526 5122
rect 41010 5070 41022 5122
rect 41074 5070 41086 5122
rect 32510 5058 32562 5070
rect 41582 5058 41634 5070
rect 42254 5122 42306 5134
rect 48078 5122 48130 5134
rect 44594 5070 44606 5122
rect 44658 5070 44670 5122
rect 42254 5058 42306 5070
rect 48078 5058 48130 5070
rect 48638 5122 48690 5134
rect 52558 5122 52610 5134
rect 52210 5070 52222 5122
rect 52274 5070 52286 5122
rect 48638 5058 48690 5070
rect 52558 5058 52610 5070
rect 53454 5122 53506 5134
rect 69470 5122 69522 5134
rect 76638 5122 76690 5134
rect 84478 5122 84530 5134
rect 60386 5070 60398 5122
rect 60450 5070 60462 5122
rect 66658 5070 66670 5122
rect 66722 5070 66734 5122
rect 70466 5070 70478 5122
rect 70530 5070 70542 5122
rect 76066 5070 76078 5122
rect 76130 5070 76142 5122
rect 77298 5070 77310 5122
rect 77362 5070 77374 5122
rect 53454 5058 53506 5070
rect 69470 5058 69522 5070
rect 76638 5058 76690 5070
rect 84478 5058 84530 5070
rect 85486 5122 85538 5134
rect 89518 5122 89570 5134
rect 85922 5070 85934 5122
rect 85986 5070 85998 5122
rect 85486 5058 85538 5070
rect 89518 5058 89570 5070
rect 93662 5122 93714 5134
rect 93662 5058 93714 5070
rect 95230 5122 95282 5134
rect 104190 5122 104242 5134
rect 109230 5122 109282 5134
rect 112030 5122 112082 5134
rect 117182 5122 117234 5134
rect 120654 5122 120706 5134
rect 127374 5122 127426 5134
rect 95554 5070 95566 5122
rect 95618 5070 95630 5122
rect 105298 5070 105310 5122
rect 105362 5070 105374 5122
rect 108098 5070 108110 5122
rect 108162 5070 108174 5122
rect 110338 5070 110350 5122
rect 110402 5070 110414 5122
rect 112354 5070 112366 5122
rect 112418 5070 112430 5122
rect 117618 5070 117630 5122
rect 117682 5070 117694 5122
rect 125010 5070 125022 5122
rect 125074 5070 125086 5122
rect 95230 5058 95282 5070
rect 104190 5058 104242 5070
rect 109230 5058 109282 5070
rect 112030 5058 112082 5070
rect 117182 5058 117234 5070
rect 120654 5058 120706 5070
rect 127374 5058 127426 5070
rect 127822 5122 127874 5134
rect 131966 5122 132018 5134
rect 136334 5122 136386 5134
rect 141710 5122 141762 5134
rect 128370 5070 128382 5122
rect 128434 5070 128446 5122
rect 135874 5070 135886 5122
rect 135938 5070 135950 5122
rect 139122 5070 139134 5122
rect 139186 5070 139198 5122
rect 127822 5058 127874 5070
rect 131966 5058 132018 5070
rect 136334 5058 136386 5070
rect 141710 5058 141762 5070
rect 142270 5122 142322 5134
rect 142270 5058 142322 5070
rect 143502 5122 143554 5134
rect 145170 5070 145182 5122
rect 145234 5070 145246 5122
rect 143502 5058 143554 5070
rect 11790 5010 11842 5022
rect 11790 4946 11842 4958
rect 12238 5010 12290 5022
rect 36766 5010 36818 5022
rect 14130 4958 14142 5010
rect 14194 4958 14206 5010
rect 34290 4958 34302 5010
rect 34354 4958 34366 5010
rect 12238 4946 12290 4958
rect 36766 4946 36818 4958
rect 38222 5010 38274 5022
rect 49870 5010 49922 5022
rect 43586 4958 43598 5010
rect 43650 4958 43662 5010
rect 45602 4958 45614 5010
rect 45666 4958 45678 5010
rect 38222 4946 38274 4958
rect 49870 4946 49922 4958
rect 56478 5010 56530 5022
rect 56478 4946 56530 4958
rect 57822 5010 57874 5022
rect 57822 4946 57874 4958
rect 58158 5010 58210 5022
rect 71486 5010 71538 5022
rect 67890 4958 67902 5010
rect 67954 4958 67966 5010
rect 68226 4958 68238 5010
rect 68290 4958 68302 5010
rect 58158 4946 58210 4958
rect 71486 4946 71538 4958
rect 71934 5010 71986 5022
rect 90750 5010 90802 5022
rect 82226 4958 82238 5010
rect 82290 4958 82302 5010
rect 71934 4946 71986 4958
rect 90750 4946 90802 4958
rect 91086 5010 91138 5022
rect 91086 4946 91138 4958
rect 94222 5010 94274 5022
rect 94222 4946 94274 4958
rect 94558 5010 94610 5022
rect 94558 4946 94610 4958
rect 111022 5010 111074 5022
rect 111022 4946 111074 4958
rect 137342 5010 137394 5022
rect 138898 4958 138910 5010
rect 138962 4958 138974 5010
rect 145058 4958 145070 5010
rect 145122 4958 145134 5010
rect 137342 4946 137394 4958
rect 11118 4898 11170 4910
rect 11118 4834 11170 4846
rect 16382 4898 16434 4910
rect 21646 4898 21698 4910
rect 33742 4898 33794 4910
rect 20290 4846 20302 4898
rect 20354 4846 20366 4898
rect 28130 4846 28142 4898
rect 28194 4846 28206 4898
rect 16382 4834 16434 4846
rect 21646 4834 21698 4846
rect 33742 4834 33794 4846
rect 36430 4898 36482 4910
rect 36430 4834 36482 4846
rect 48526 4898 48578 4910
rect 48526 4834 48578 4846
rect 55918 4898 55970 4910
rect 55918 4834 55970 4846
rect 56814 4898 56866 4910
rect 56814 4834 56866 4846
rect 57262 4898 57314 4910
rect 57262 4834 57314 4846
rect 58830 4898 58882 4910
rect 58830 4834 58882 4846
rect 71150 4898 71202 4910
rect 71150 4834 71202 4846
rect 72606 4898 72658 4910
rect 91758 4898 91810 4910
rect 102062 4898 102114 4910
rect 73714 4846 73726 4898
rect 73778 4846 73790 4898
rect 88386 4846 88398 4898
rect 88450 4846 88462 4898
rect 97906 4846 97918 4898
rect 97970 4846 97982 4898
rect 72606 4834 72658 4846
rect 91758 4834 91810 4846
rect 102062 4834 102114 4846
rect 108334 4898 108386 4910
rect 108334 4834 108386 4846
rect 111358 4898 111410 4910
rect 137006 4898 137058 4910
rect 114930 4846 114942 4898
rect 114994 4846 115006 4898
rect 120082 4846 120094 4898
rect 120146 4846 120158 4898
rect 130946 4846 130958 4898
rect 131010 4846 131022 4898
rect 133410 4846 133422 4898
rect 133474 4846 133486 4898
rect 111358 4834 111410 4846
rect 137006 4834 137058 4846
rect 144174 4898 144226 4910
rect 144174 4834 144226 4846
rect 1344 4730 148784 4764
rect 1344 4678 38034 4730
rect 38086 4678 38138 4730
rect 38190 4678 38242 4730
rect 38294 4678 74854 4730
rect 74906 4678 74958 4730
rect 75010 4678 75062 4730
rect 75114 4678 111674 4730
rect 111726 4678 111778 4730
rect 111830 4678 111882 4730
rect 111934 4678 148494 4730
rect 148546 4678 148598 4730
rect 148650 4678 148702 4730
rect 148754 4678 148784 4730
rect 1344 4644 148784 4678
rect 12014 4562 12066 4574
rect 16942 4562 16994 4574
rect 16034 4510 16046 4562
rect 16098 4510 16110 4562
rect 12014 4498 12066 4510
rect 16942 4498 16994 4510
rect 28142 4562 28194 4574
rect 39118 4562 39170 4574
rect 48862 4562 48914 4574
rect 38546 4510 38558 4562
rect 38610 4510 38622 4562
rect 48290 4510 48302 4562
rect 48354 4510 48366 4562
rect 28142 4498 28194 4510
rect 39118 4498 39170 4510
rect 48862 4498 48914 4510
rect 51550 4562 51602 4574
rect 51550 4498 51602 4510
rect 55022 4562 55074 4574
rect 55022 4498 55074 4510
rect 60622 4562 60674 4574
rect 64766 4562 64818 4574
rect 64194 4510 64206 4562
rect 64258 4510 64270 4562
rect 60622 4498 60674 4510
rect 64766 4498 64818 4510
rect 81230 4562 81282 4574
rect 81230 4498 81282 4510
rect 81678 4562 81730 4574
rect 81678 4498 81730 4510
rect 85598 4562 85650 4574
rect 85598 4498 85650 4510
rect 86270 4562 86322 4574
rect 92878 4562 92930 4574
rect 92082 4510 92094 4562
rect 92146 4510 92158 4562
rect 86270 4498 86322 4510
rect 92878 4498 92930 4510
rect 97134 4562 97186 4574
rect 97134 4498 97186 4510
rect 97918 4562 97970 4574
rect 97918 4498 97970 4510
rect 98366 4562 98418 4574
rect 107550 4562 107602 4574
rect 116734 4562 116786 4574
rect 102498 4510 102510 4562
rect 102562 4510 102574 4562
rect 111122 4510 111134 4562
rect 111186 4510 111198 4562
rect 116162 4510 116174 4562
rect 116226 4510 116238 4562
rect 98366 4498 98418 4510
rect 107550 4498 107602 4510
rect 116734 4498 116786 4510
rect 118974 4562 119026 4574
rect 118974 4498 119026 4510
rect 124238 4562 124290 4574
rect 128382 4562 128434 4574
rect 134878 4562 134930 4574
rect 127810 4510 127822 4562
rect 127874 4510 127886 4562
rect 131842 4510 131854 4562
rect 131906 4510 131918 4562
rect 124238 4498 124290 4510
rect 128382 4498 128434 4510
rect 134878 4498 134930 4510
rect 135886 4562 135938 4574
rect 135886 4498 135938 4510
rect 143726 4562 143778 4574
rect 143726 4498 143778 4510
rect 146750 4562 146802 4574
rect 146750 4498 146802 4510
rect 12126 4450 12178 4462
rect 33518 4450 33570 4462
rect 59502 4450 59554 4462
rect 86830 4450 86882 4462
rect 7410 4398 7422 4450
rect 7474 4398 7486 4450
rect 10994 4398 11006 4450
rect 11058 4398 11070 4450
rect 21074 4398 21086 4450
rect 21138 4398 21150 4450
rect 22194 4398 22206 4450
rect 22258 4398 22270 4450
rect 26226 4398 26238 4450
rect 26290 4398 26302 4450
rect 28914 4398 28926 4450
rect 28978 4398 28990 4450
rect 32722 4398 32734 4450
rect 32786 4398 32798 4450
rect 41682 4398 41694 4450
rect 41746 4398 41758 4450
rect 49634 4398 49646 4450
rect 49698 4398 49710 4450
rect 53106 4398 53118 4450
rect 53170 4398 53182 4450
rect 57586 4398 57598 4450
rect 57650 4398 57662 4450
rect 68674 4398 68686 4450
rect 68738 4398 68750 4450
rect 80322 4398 80334 4450
rect 80386 4398 80398 4450
rect 12126 4386 12178 4398
rect 33518 4386 33570 4398
rect 59502 4386 59554 4398
rect 86830 4386 86882 4398
rect 97806 4450 97858 4462
rect 97806 4386 97858 4398
rect 103182 4450 103234 4462
rect 103182 4386 103234 4398
rect 119310 4450 119362 4462
rect 119310 4386 119362 4398
rect 119870 4450 119922 4462
rect 119870 4386 119922 4398
rect 135214 4450 135266 4462
rect 135214 4386 135266 4398
rect 136222 4450 136274 4462
rect 144062 4450 144114 4462
rect 137778 4398 137790 4450
rect 137842 4398 137854 4450
rect 141810 4398 141822 4450
rect 141874 4398 141886 4450
rect 145618 4398 145630 4450
rect 145682 4398 145694 4450
rect 145954 4398 145966 4450
rect 146018 4398 146030 4450
rect 136222 4386 136274 4398
rect 144062 4386 144114 4398
rect 12910 4338 12962 4350
rect 59838 4338 59890 4350
rect 5842 4286 5854 4338
rect 5906 4286 5918 4338
rect 13570 4286 13582 4338
rect 13634 4286 13646 4338
rect 19394 4286 19406 4338
rect 19458 4286 19470 4338
rect 35522 4286 35534 4338
rect 35586 4286 35598 4338
rect 36082 4286 36094 4338
rect 36146 4286 36158 4338
rect 39554 4286 39566 4338
rect 39618 4286 39630 4338
rect 45266 4286 45278 4338
rect 45330 4286 45342 4338
rect 45826 4286 45838 4338
rect 45890 4286 45902 4338
rect 56466 4286 56478 4338
rect 56530 4286 56542 4338
rect 12910 4274 12962 4286
rect 59838 4274 59890 4286
rect 61070 4338 61122 4350
rect 89182 4338 89234 4350
rect 99038 4338 99090 4350
rect 61730 4286 61742 4338
rect 61794 4286 61806 4338
rect 69234 4286 69246 4338
rect 69298 4286 69310 4338
rect 72370 4286 72382 4338
rect 72434 4286 72446 4338
rect 74610 4286 74622 4338
rect 74674 4286 74686 4338
rect 75618 4286 75630 4338
rect 75682 4286 75694 4338
rect 85138 4286 85150 4338
rect 85202 4286 85214 4338
rect 88498 4286 88510 4338
rect 88562 4286 88574 4338
rect 89730 4286 89742 4338
rect 89794 4286 89806 4338
rect 94546 4286 94558 4338
rect 94610 4286 94622 4338
rect 96450 4286 96462 4338
rect 96514 4286 96526 4338
rect 61070 4274 61122 4286
rect 89182 4274 89234 4286
rect 99038 4274 99090 4286
rect 99486 4338 99538 4350
rect 108222 4338 108274 4350
rect 112030 4338 112082 4350
rect 100034 4286 100046 4338
rect 100098 4286 100110 4338
rect 108546 4286 108558 4338
rect 108610 4286 108622 4338
rect 99486 4274 99538 4286
rect 108222 4274 108274 4286
rect 112030 4274 112082 4286
rect 113038 4338 113090 4350
rect 119982 4338 120034 4350
rect 124686 4338 124738 4350
rect 129166 4338 129218 4350
rect 136894 4338 136946 4350
rect 113586 4286 113598 4338
rect 113650 4286 113662 4338
rect 118178 4286 118190 4338
rect 118242 4286 118254 4338
rect 121090 4286 121102 4338
rect 121154 4286 121166 4338
rect 125346 4286 125358 4338
rect 125410 4286 125422 4338
rect 129602 4286 129614 4338
rect 129666 4286 129678 4338
rect 134306 4286 134318 4338
rect 134370 4286 134382 4338
rect 113038 4274 113090 4286
rect 119982 4274 120034 4286
rect 124686 4274 124738 4286
rect 129166 4274 129218 4286
rect 136894 4274 136946 4286
rect 145406 4338 145458 4350
rect 145406 4274 145458 4286
rect 6414 4226 6466 4238
rect 4722 4174 4734 4226
rect 4786 4174 4798 4226
rect 6414 4162 6466 4174
rect 6862 4226 6914 4238
rect 17726 4226 17778 4238
rect 25678 4226 25730 4238
rect 28254 4226 28306 4238
rect 30718 4226 30770 4238
rect 52558 4226 52610 4238
rect 111694 4226 111746 4238
rect 141262 4226 141314 4238
rect 147198 4226 147250 4238
rect 8754 4174 8766 4226
rect 8818 4174 8830 4226
rect 9986 4174 9998 4226
rect 10050 4174 10062 4226
rect 18834 4174 18846 4226
rect 18898 4174 18910 4226
rect 20066 4174 20078 4226
rect 20130 4174 20142 4226
rect 23538 4174 23550 4226
rect 23602 4174 23614 4226
rect 27570 4174 27582 4226
rect 27634 4174 27646 4226
rect 30258 4174 30270 4226
rect 30322 4174 30334 4226
rect 31378 4174 31390 4226
rect 31442 4174 31454 4226
rect 40338 4174 40350 4226
rect 40402 4174 40414 4226
rect 42802 4174 42814 4226
rect 42866 4174 42878 4226
rect 50754 4174 50766 4226
rect 50818 4174 50830 4226
rect 54226 4174 54238 4226
rect 54290 4174 54302 4226
rect 55570 4174 55582 4226
rect 55634 4174 55646 4226
rect 58930 4174 58942 4226
rect 58994 4174 59006 4226
rect 71586 4174 71598 4226
rect 71650 4174 71662 4226
rect 73826 4174 73838 4226
rect 73890 4174 73902 4226
rect 84018 4174 84030 4226
rect 84082 4174 84094 4226
rect 87714 4174 87726 4226
rect 87778 4174 87790 4226
rect 93426 4174 93438 4226
rect 93490 4174 93502 4226
rect 95778 4174 95790 4226
rect 95842 4174 95854 4226
rect 117282 4174 117294 4226
rect 117346 4174 117358 4226
rect 121762 4174 121774 4226
rect 121826 4174 121838 4226
rect 133186 4174 133198 4226
rect 133250 4174 133262 4226
rect 138898 4174 138910 4226
rect 138962 4174 138974 4226
rect 143154 4174 143166 4226
rect 143218 4174 143230 4226
rect 6862 4162 6914 4174
rect 17726 4162 17778 4174
rect 25678 4162 25730 4174
rect 28254 4162 28306 4174
rect 30718 4162 30770 4174
rect 52558 4162 52610 4174
rect 111694 4162 111746 4174
rect 141262 4162 141314 4174
rect 147198 4162 147250 4174
rect 16606 4114 16658 4126
rect 16606 4050 16658 4062
rect 132638 4114 132690 4126
rect 132638 4050 132690 4062
rect 145070 4114 145122 4126
rect 145070 4050 145122 4062
rect 1344 3946 148624 3980
rect 1344 3894 19624 3946
rect 19676 3894 19728 3946
rect 19780 3894 19832 3946
rect 19884 3894 56444 3946
rect 56496 3894 56548 3946
rect 56600 3894 56652 3946
rect 56704 3894 93264 3946
rect 93316 3894 93368 3946
rect 93420 3894 93472 3946
rect 93524 3894 130084 3946
rect 130136 3894 130188 3946
rect 130240 3894 130292 3946
rect 130344 3894 148624 3946
rect 1344 3860 148624 3894
rect 14366 3778 14418 3790
rect 9650 3726 9662 3778
rect 9714 3726 9726 3778
rect 14366 3714 14418 3726
rect 63870 3778 63922 3790
rect 63870 3714 63922 3726
rect 67678 3778 67730 3790
rect 67678 3714 67730 3726
rect 68462 3778 68514 3790
rect 68462 3714 68514 3726
rect 71710 3778 71762 3790
rect 71710 3714 71762 3726
rect 75630 3778 75682 3790
rect 75630 3714 75682 3726
rect 79214 3778 79266 3790
rect 79214 3714 79266 3726
rect 80222 3778 80274 3790
rect 80222 3714 80274 3726
rect 80782 3778 80834 3790
rect 80782 3714 80834 3726
rect 84702 3778 84754 3790
rect 84702 3714 84754 3726
rect 88622 3778 88674 3790
rect 88622 3714 88674 3726
rect 92542 3778 92594 3790
rect 92542 3714 92594 3726
rect 111694 3778 111746 3790
rect 111694 3714 111746 3726
rect 115502 3778 115554 3790
rect 115502 3714 115554 3726
rect 116174 3778 116226 3790
rect 116174 3714 116226 3726
rect 119534 3778 119586 3790
rect 131518 3778 131570 3790
rect 119746 3726 119758 3778
rect 119810 3775 119822 3778
rect 120530 3775 120542 3778
rect 119810 3729 120542 3775
rect 119810 3726 119822 3729
rect 120530 3726 120542 3729
rect 120594 3726 120606 3778
rect 119534 3714 119586 3726
rect 131518 3714 131570 3726
rect 132302 3778 132354 3790
rect 132302 3714 132354 3726
rect 6974 3666 7026 3678
rect 13918 3666 13970 3678
rect 30046 3666 30098 3678
rect 40238 3666 40290 3678
rect 64654 3666 64706 3678
rect 8866 3614 8878 3666
rect 8930 3614 8942 3666
rect 11330 3614 11342 3666
rect 11394 3614 11406 3666
rect 15250 3614 15262 3666
rect 15314 3614 15326 3666
rect 18722 3614 18734 3666
rect 18786 3614 18798 3666
rect 23314 3614 23326 3666
rect 23378 3614 23390 3666
rect 28466 3614 28478 3666
rect 28530 3614 28542 3666
rect 31154 3614 31166 3666
rect 31218 3614 31230 3666
rect 34850 3614 34862 3666
rect 34914 3614 34926 3666
rect 39666 3614 39678 3666
rect 39730 3614 39742 3666
rect 43698 3614 43710 3666
rect 43762 3614 43774 3666
rect 47506 3614 47518 3666
rect 47570 3614 47582 3666
rect 51538 3614 51550 3666
rect 51602 3614 51614 3666
rect 55682 3614 55694 3666
rect 55746 3614 55758 3666
rect 59602 3614 59614 3666
rect 59666 3614 59678 3666
rect 6974 3602 7026 3614
rect 13918 3602 13970 3614
rect 30046 3602 30098 3614
rect 40238 3602 40290 3614
rect 64654 3602 64706 3614
rect 68574 3666 68626 3678
rect 68574 3602 68626 3614
rect 76302 3666 76354 3678
rect 76302 3602 76354 3614
rect 76750 3666 76802 3678
rect 79326 3666 79378 3678
rect 78418 3614 78430 3666
rect 78482 3614 78494 3666
rect 76750 3602 76802 3614
rect 79326 3602 79378 3614
rect 80334 3666 80386 3678
rect 80334 3602 80386 3614
rect 95902 3666 95954 3678
rect 108334 3666 108386 3678
rect 119982 3666 120034 3678
rect 98802 3614 98814 3666
rect 98866 3614 98878 3666
rect 102834 3614 102846 3666
rect 102898 3614 102910 3666
rect 106642 3614 106654 3666
rect 106706 3614 106718 3666
rect 110562 3614 110574 3666
rect 110626 3614 110638 3666
rect 113250 3614 113262 3666
rect 113314 3614 113326 3666
rect 117170 3614 117182 3666
rect 117234 3614 117246 3666
rect 95902 3602 95954 3614
rect 108334 3602 108386 3614
rect 119982 3602 120034 3614
rect 120430 3666 120482 3678
rect 128046 3666 128098 3678
rect 121202 3614 121214 3666
rect 121266 3614 121278 3666
rect 125122 3614 125134 3666
rect 125186 3614 125198 3666
rect 120430 3602 120482 3614
rect 128046 3602 128098 3614
rect 128494 3666 128546 3678
rect 131630 3666 131682 3678
rect 129042 3614 129054 3666
rect 129106 3614 129118 3666
rect 128494 3602 128546 3614
rect 131630 3602 131682 3614
rect 132190 3666 132242 3678
rect 135214 3666 135266 3678
rect 134306 3614 134318 3666
rect 134370 3614 134382 3666
rect 132190 3602 132242 3614
rect 135214 3602 135266 3614
rect 139022 3666 139074 3678
rect 139022 3602 139074 3614
rect 139918 3666 139970 3678
rect 141026 3614 141038 3666
rect 141090 3614 141102 3666
rect 144610 3614 144622 3666
rect 144674 3614 144686 3666
rect 147522 3614 147534 3666
rect 147586 3614 147598 3666
rect 139918 3602 139970 3614
rect 6302 3554 6354 3566
rect 6302 3490 6354 3502
rect 6414 3554 6466 3566
rect 6414 3490 6466 3502
rect 6638 3554 6690 3566
rect 6638 3490 6690 3502
rect 10222 3554 10274 3566
rect 19406 3554 19458 3566
rect 60846 3554 60898 3566
rect 14690 3502 14702 3554
rect 14754 3502 14766 3554
rect 29474 3502 29486 3554
rect 29538 3502 29550 3554
rect 10222 3490 10274 3502
rect 19406 3490 19458 3502
rect 60846 3490 60898 3502
rect 72606 3554 72658 3566
rect 72606 3490 72658 3502
rect 111806 3554 111858 3566
rect 123230 3554 123282 3566
rect 112578 3502 112590 3554
rect 112642 3502 112654 3554
rect 111806 3490 111858 3502
rect 123230 3490 123282 3502
rect 135662 3554 135714 3566
rect 144062 3554 144114 3566
rect 137330 3502 137342 3554
rect 137394 3502 137406 3554
rect 140354 3502 140366 3554
rect 140418 3502 140430 3554
rect 146850 3502 146862 3554
rect 146914 3502 146926 3554
rect 135662 3490 135714 3502
rect 144062 3490 144114 3502
rect 6862 3442 6914 3454
rect 10110 3442 10162 3454
rect 7858 3390 7870 3442
rect 7922 3390 7934 3442
rect 6862 3378 6914 3390
rect 10110 3378 10162 3390
rect 10334 3442 10386 3454
rect 14478 3442 14530 3454
rect 21870 3442 21922 3454
rect 12338 3390 12350 3442
rect 12402 3390 12414 3442
rect 16258 3390 16270 3442
rect 16322 3390 16334 3442
rect 17602 3390 17614 3442
rect 17666 3390 17678 3442
rect 10334 3378 10386 3390
rect 14478 3378 14530 3390
rect 21870 3378 21922 3390
rect 22206 3442 22258 3454
rect 25230 3442 25282 3454
rect 24098 3390 24110 3442
rect 24162 3390 24174 3442
rect 22206 3378 22258 3390
rect 25230 3378 25282 3390
rect 26574 3442 26626 3454
rect 33070 3442 33122 3454
rect 36990 3442 37042 3454
rect 27234 3390 27246 3442
rect 27298 3390 27310 3442
rect 32274 3390 32286 3442
rect 32338 3390 32350 3442
rect 36194 3390 36206 3442
rect 36258 3390 36270 3442
rect 26574 3378 26626 3390
rect 33070 3378 33122 3390
rect 36990 3378 37042 3390
rect 37774 3442 37826 3454
rect 41246 3442 41298 3454
rect 38322 3390 38334 3442
rect 38386 3390 38398 3442
rect 37774 3378 37826 3390
rect 41246 3378 41298 3390
rect 41806 3442 41858 3454
rect 45838 3442 45890 3454
rect 48862 3442 48914 3454
rect 42354 3390 42366 3442
rect 42418 3390 42430 3442
rect 46386 3390 46398 3442
rect 46450 3390 46462 3442
rect 41806 3378 41858 3390
rect 45838 3378 45890 3390
rect 48862 3378 48914 3390
rect 49198 3442 49250 3454
rect 49198 3378 49250 3390
rect 49870 3442 49922 3454
rect 53902 3442 53954 3454
rect 56702 3442 56754 3454
rect 50418 3390 50430 3442
rect 50482 3390 50494 3442
rect 54450 3390 54462 3442
rect 54514 3390 54526 3442
rect 49870 3378 49922 3390
rect 53902 3378 53954 3390
rect 56702 3378 56754 3390
rect 57934 3442 57986 3454
rect 84030 3442 84082 3454
rect 87950 3442 88002 3454
rect 91870 3442 91922 3454
rect 96238 3442 96290 3454
rect 58482 3390 58494 3442
rect 58546 3390 58558 3442
rect 61730 3390 61742 3442
rect 61794 3390 61806 3442
rect 65202 3390 65214 3442
rect 65266 3390 65278 3442
rect 69570 3390 69582 3442
rect 69634 3390 69646 3442
rect 73154 3390 73166 3442
rect 73218 3390 73230 3442
rect 77298 3390 77310 3442
rect 77362 3390 77374 3442
rect 82898 3390 82910 3442
rect 82962 3390 82974 3442
rect 86818 3390 86830 3442
rect 86882 3390 86894 3442
rect 91074 3390 91086 3442
rect 91138 3390 91150 3442
rect 94658 3390 94670 3442
rect 94722 3390 94734 3442
rect 57934 3378 57986 3390
rect 84030 3378 84082 3390
rect 87950 3378 88002 3390
rect 91870 3378 91922 3390
rect 96238 3378 96290 3390
rect 96910 3442 96962 3454
rect 100942 3442 100994 3454
rect 104974 3442 105026 3454
rect 108894 3442 108946 3454
rect 112366 3442 112418 3454
rect 115614 3442 115666 3454
rect 97458 3390 97470 3442
rect 97522 3390 97534 3442
rect 101490 3390 101502 3442
rect 101554 3390 101566 3442
rect 105522 3390 105534 3442
rect 105586 3390 105598 3442
rect 109442 3390 109454 3442
rect 109506 3390 109518 3442
rect 114594 3390 114606 3442
rect 114658 3390 114670 3442
rect 96910 3378 96962 3390
rect 100942 3378 100994 3390
rect 104974 3378 105026 3390
rect 108894 3378 108946 3390
rect 112366 3378 112418 3390
rect 115614 3378 115666 3390
rect 116286 3442 116338 3454
rect 119422 3442 119474 3454
rect 123678 3442 123730 3454
rect 127150 3442 127202 3454
rect 135102 3442 135154 3454
rect 138014 3442 138066 3454
rect 118514 3390 118526 3442
rect 118578 3390 118590 3442
rect 122098 3390 122110 3442
rect 122162 3390 122174 3442
rect 126354 3390 126366 3442
rect 126418 3390 126430 3442
rect 130274 3390 130286 3442
rect 130338 3390 130350 3442
rect 133298 3390 133310 3442
rect 133362 3390 133374 3442
rect 136434 3390 136446 3442
rect 136498 3390 136510 3442
rect 145618 3390 145630 3442
rect 145682 3390 145694 3442
rect 116286 3378 116338 3390
rect 119422 3378 119474 3390
rect 123678 3378 123730 3390
rect 127150 3378 127202 3390
rect 135102 3378 135154 3390
rect 138014 3378 138066 3390
rect 29262 3330 29314 3342
rect 29262 3266 29314 3278
rect 57038 3330 57090 3342
rect 57038 3266 57090 3278
rect 143726 3330 143778 3342
rect 143726 3266 143778 3278
rect 1344 3162 148784 3196
rect 1344 3110 38034 3162
rect 38086 3110 38138 3162
rect 38190 3110 38242 3162
rect 38294 3110 74854 3162
rect 74906 3110 74958 3162
rect 75010 3110 75062 3162
rect 75114 3110 111674 3162
rect 111726 3110 111778 3162
rect 111830 3110 111882 3162
rect 111934 3110 148494 3162
rect 148546 3110 148598 3162
rect 148650 3110 148702 3162
rect 148754 3110 148784 3162
rect 1344 3076 148784 3110
<< via1 >>
rect 82574 37326 82626 37378
rect 83806 37326 83858 37378
rect 19624 36822 19676 36874
rect 19728 36822 19780 36874
rect 19832 36822 19884 36874
rect 56444 36822 56496 36874
rect 56548 36822 56600 36874
rect 56652 36822 56704 36874
rect 93264 36822 93316 36874
rect 93368 36822 93420 36874
rect 93472 36822 93524 36874
rect 130084 36822 130136 36874
rect 130188 36822 130240 36874
rect 130292 36822 130344 36874
rect 40798 36654 40850 36706
rect 41358 36654 41410 36706
rect 77534 36654 77586 36706
rect 8878 36542 8930 36594
rect 12798 36542 12850 36594
rect 13918 36542 13970 36594
rect 16718 36542 16770 36594
rect 20638 36542 20690 36594
rect 24222 36542 24274 36594
rect 26910 36542 26962 36594
rect 27694 36542 27746 36594
rect 32286 36542 32338 36594
rect 36318 36542 36370 36594
rect 40238 36542 40290 36594
rect 43934 36542 43986 36594
rect 48078 36542 48130 36594
rect 51998 36542 52050 36594
rect 55694 36542 55746 36594
rect 59726 36542 59778 36594
rect 63646 36542 63698 36594
rect 64766 36542 64818 36594
rect 67230 36542 67282 36594
rect 67678 36542 67730 36594
rect 68462 36542 68514 36594
rect 70814 36542 70866 36594
rect 71710 36542 71762 36594
rect 75518 36542 75570 36594
rect 77198 36542 77250 36594
rect 78990 36542 79042 36594
rect 80222 36542 80274 36594
rect 85822 36542 85874 36594
rect 89742 36542 89794 36594
rect 92766 36542 92818 36594
rect 93550 36542 93602 36594
rect 96238 36542 96290 36594
rect 99822 36542 99874 36594
rect 104414 36542 104466 36594
rect 107886 36542 107938 36594
rect 111582 36542 111634 36594
rect 115502 36542 115554 36594
rect 119422 36542 119474 36594
rect 122222 36542 122274 36594
rect 123342 36542 123394 36594
rect 129054 36542 129106 36594
rect 132638 36542 132690 36594
rect 135102 36542 135154 36594
rect 139022 36542 139074 36594
rect 144174 36542 144226 36594
rect 147534 36542 147586 36594
rect 6638 36430 6690 36482
rect 33518 36430 33570 36482
rect 37438 36430 37490 36482
rect 45950 36430 46002 36482
rect 49198 36430 49250 36482
rect 53118 36430 53170 36482
rect 53790 36430 53842 36482
rect 65102 36430 65154 36482
rect 73502 36430 73554 36482
rect 78206 36430 78258 36482
rect 88398 36430 88450 36482
rect 89070 36430 89122 36482
rect 98366 36430 98418 36482
rect 102734 36430 102786 36482
rect 103630 36430 103682 36482
rect 106878 36430 106930 36482
rect 129838 36430 129890 36482
rect 141822 36430 141874 36482
rect 145742 36430 145794 36482
rect 146862 36430 146914 36482
rect 4846 36318 4898 36370
rect 7870 36318 7922 36370
rect 10782 36318 10834 36370
rect 11678 36318 11730 36370
rect 14702 36318 14754 36370
rect 15374 36318 15426 36370
rect 18286 36318 18338 36370
rect 19294 36318 19346 36370
rect 21422 36318 21474 36370
rect 22206 36318 22258 36370
rect 22878 36318 22930 36370
rect 25566 36318 25618 36370
rect 28142 36318 28194 36370
rect 29262 36318 29314 36370
rect 29822 36318 29874 36370
rect 30942 36318 30994 36370
rect 34302 36318 34354 36370
rect 35086 36318 35138 36370
rect 38222 36318 38274 36370
rect 38894 36318 38946 36370
rect 41918 36318 41970 36370
rect 42590 36318 42642 36370
rect 45278 36318 45330 36370
rect 46846 36318 46898 36370
rect 49646 36318 49698 36370
rect 50990 36318 51042 36370
rect 54798 36318 54850 36370
rect 57486 36318 57538 36370
rect 58494 36318 58546 36370
rect 60846 36318 60898 36370
rect 61630 36318 61682 36370
rect 62302 36318 62354 36370
rect 65886 36318 65938 36370
rect 68910 36318 68962 36370
rect 69470 36318 69522 36370
rect 72382 36318 72434 36370
rect 73166 36318 73218 36370
rect 74510 36318 74562 36370
rect 76414 36318 76466 36370
rect 76862 36318 76914 36370
rect 81230 36318 81282 36370
rect 82238 36318 82290 36370
rect 82574 36318 82626 36370
rect 83022 36318 83074 36370
rect 84142 36318 84194 36370
rect 86830 36318 86882 36370
rect 90750 36318 90802 36370
rect 91982 36318 92034 36370
rect 94558 36318 94610 36370
rect 97470 36318 97522 36370
rect 99038 36318 99090 36370
rect 100830 36318 100882 36370
rect 105310 36318 105362 36370
rect 108894 36318 108946 36370
rect 109902 36318 109954 36370
rect 110238 36318 110290 36370
rect 112590 36318 112642 36370
rect 113598 36318 113650 36370
rect 114382 36318 114434 36370
rect 116510 36318 116562 36370
rect 117518 36318 117570 36370
rect 118302 36318 118354 36370
rect 120430 36318 120482 36370
rect 121774 36318 121826 36370
rect 124350 36318 124402 36370
rect 125358 36318 125410 36370
rect 125694 36318 125746 36370
rect 126142 36318 126194 36370
rect 127710 36318 127762 36370
rect 130398 36318 130450 36370
rect 131294 36318 131346 36370
rect 133534 36318 133586 36370
rect 136110 36318 136162 36370
rect 137118 36318 137170 36370
rect 140030 36318 140082 36370
rect 142158 36318 142210 36370
rect 143054 36318 143106 36370
rect 145294 36318 145346 36370
rect 6078 36206 6130 36258
rect 6862 36206 6914 36258
rect 9998 36206 10050 36258
rect 10446 36206 10498 36258
rect 14366 36206 14418 36258
rect 17838 36206 17890 36258
rect 18622 36206 18674 36258
rect 21870 36206 21922 36258
rect 28478 36206 28530 36258
rect 30158 36206 30210 36258
rect 33966 36206 34018 36258
rect 37886 36206 37938 36258
rect 41134 36206 41186 36258
rect 41582 36206 41634 36258
rect 45726 36206 45778 36258
rect 49982 36206 50034 36258
rect 53566 36206 53618 36258
rect 57038 36206 57090 36258
rect 57822 36206 57874 36258
rect 61294 36206 61346 36258
rect 72494 36206 72546 36258
rect 72718 36206 72770 36258
rect 84478 36206 84530 36258
rect 84926 36206 84978 36258
rect 88622 36206 88674 36258
rect 92318 36206 92370 36258
rect 98590 36206 98642 36258
rect 102174 36206 102226 36258
rect 106318 36206 106370 36258
rect 110686 36206 110738 36258
rect 113934 36206 113986 36258
rect 117854 36206 117906 36258
rect 121438 36206 121490 36258
rect 129614 36206 129666 36258
rect 133198 36206 133250 36258
rect 133982 36206 134034 36258
rect 137454 36206 137506 36258
rect 138014 36206 138066 36258
rect 140926 36206 140978 36258
rect 144958 36206 145010 36258
rect 38034 36038 38086 36090
rect 38138 36038 38190 36090
rect 38242 36038 38294 36090
rect 74854 36038 74906 36090
rect 74958 36038 75010 36090
rect 75062 36038 75114 36090
rect 111674 36038 111726 36090
rect 111778 36038 111830 36090
rect 111882 36038 111934 36090
rect 148494 36038 148546 36090
rect 148598 36038 148650 36090
rect 148702 36038 148754 36090
rect 9662 35870 9714 35922
rect 21422 35870 21474 35922
rect 35758 35870 35810 35922
rect 43598 35870 43650 35922
rect 48414 35870 48466 35922
rect 59502 35870 59554 35922
rect 69694 35870 69746 35922
rect 100382 35870 100434 35922
rect 105086 35870 105138 35922
rect 132190 35870 132242 35922
rect 146862 35870 146914 35922
rect 17838 35758 17890 35810
rect 19742 35758 19794 35810
rect 21982 35758 22034 35810
rect 28254 35758 28306 35810
rect 30606 35758 30658 35810
rect 32510 35758 32562 35810
rect 33742 35758 33794 35810
rect 36542 35758 36594 35810
rect 37214 35758 37266 35810
rect 39342 35758 39394 35810
rect 41694 35758 41746 35810
rect 44158 35758 44210 35810
rect 46174 35758 46226 35810
rect 49758 35758 49810 35810
rect 52222 35758 52274 35810
rect 53342 35758 53394 35810
rect 55582 35758 55634 35810
rect 57598 35758 57650 35810
rect 60510 35758 60562 35810
rect 63646 35758 63698 35810
rect 65662 35758 65714 35810
rect 67678 35758 67730 35810
rect 70254 35758 70306 35810
rect 71262 35758 71314 35810
rect 73502 35758 73554 35810
rect 75630 35758 75682 35810
rect 76078 35758 76130 35810
rect 81678 35758 81730 35810
rect 83806 35758 83858 35810
rect 84926 35758 84978 35810
rect 86718 35758 86770 35810
rect 89518 35758 89570 35810
rect 89966 35758 90018 35810
rect 91422 35758 91474 35810
rect 93326 35758 93378 35810
rect 93774 35758 93826 35810
rect 97918 35758 97970 35810
rect 98702 35758 98754 35810
rect 102622 35758 102674 35810
rect 104078 35758 104130 35810
rect 107102 35758 107154 35810
rect 108446 35758 108498 35810
rect 108894 35758 108946 35810
rect 110910 35758 110962 35810
rect 111694 35758 111746 35810
rect 112030 35758 112082 35810
rect 114270 35758 114322 35810
rect 115614 35758 115666 35810
rect 116062 35758 116114 35810
rect 117854 35758 117906 35810
rect 119198 35758 119250 35810
rect 122110 35758 122162 35810
rect 123118 35758 123170 35810
rect 125022 35758 125074 35810
rect 126142 35758 126194 35810
rect 129502 35758 129554 35810
rect 131406 35758 131458 35810
rect 133982 35758 134034 35810
rect 138014 35758 138066 35810
rect 139358 35758 139410 35810
rect 140254 35758 140306 35810
rect 142942 35758 142994 35810
rect 143166 35758 143218 35810
rect 146190 35758 146242 35810
rect 7198 35646 7250 35698
rect 8990 35646 9042 35698
rect 10446 35646 10498 35698
rect 13358 35646 13410 35698
rect 14142 35646 14194 35698
rect 16942 35646 16994 35698
rect 18958 35646 19010 35698
rect 19630 35646 19682 35698
rect 20414 35646 20466 35698
rect 23102 35646 23154 35698
rect 24782 35646 24834 35698
rect 27582 35646 27634 35698
rect 30830 35646 30882 35698
rect 32846 35646 32898 35698
rect 36206 35646 36258 35698
rect 39230 35646 39282 35698
rect 48750 35646 48802 35698
rect 56478 35646 56530 35698
rect 59838 35646 59890 35698
rect 65550 35646 65602 35698
rect 70590 35646 70642 35698
rect 77310 35646 77362 35698
rect 79102 35646 79154 35698
rect 81342 35646 81394 35698
rect 85822 35646 85874 35698
rect 87614 35646 87666 35698
rect 88286 35646 88338 35698
rect 90190 35646 90242 35698
rect 91310 35646 91362 35698
rect 95006 35646 95058 35698
rect 97582 35646 97634 35698
rect 98590 35646 98642 35698
rect 100942 35646 100994 35698
rect 103742 35646 103794 35698
rect 105534 35646 105586 35698
rect 108110 35646 108162 35698
rect 115278 35646 115330 35698
rect 119086 35646 119138 35698
rect 123454 35646 123506 35698
rect 131630 35646 131682 35698
rect 134990 35646 135042 35698
rect 139022 35646 139074 35698
rect 142606 35646 142658 35698
rect 6414 35534 6466 35586
rect 8318 35534 8370 35586
rect 11006 35534 11058 35586
rect 12686 35534 12738 35586
rect 14590 35534 14642 35586
rect 16270 35534 16322 35586
rect 24222 35534 24274 35586
rect 25566 35534 25618 35586
rect 26798 35534 26850 35586
rect 29598 35534 29650 35586
rect 34862 35534 34914 35586
rect 38558 35534 38610 35586
rect 43038 35534 43090 35586
rect 45502 35534 45554 35586
rect 47294 35534 47346 35586
rect 51102 35534 51154 35586
rect 52670 35534 52722 35586
rect 54462 35534 54514 35586
rect 58942 35534 58994 35586
rect 61630 35534 61682 35586
rect 62638 35534 62690 35586
rect 64654 35534 64706 35586
rect 69022 35534 69074 35586
rect 72382 35534 72434 35586
rect 74846 35534 74898 35586
rect 78094 35534 78146 35586
rect 79774 35534 79826 35586
rect 82126 35534 82178 35586
rect 82798 35534 82850 35586
rect 87838 35534 87890 35586
rect 88174 35534 88226 35586
rect 92094 35534 92146 35586
rect 95902 35534 95954 35586
rect 101614 35534 101666 35586
rect 106094 35534 106146 35586
rect 109678 35534 109730 35586
rect 113262 35534 113314 35586
rect 116846 35534 116898 35586
rect 121102 35534 121154 35586
rect 124014 35534 124066 35586
rect 127486 35534 127538 35586
rect 127934 35534 127986 35586
rect 130622 35534 130674 35586
rect 132974 35534 133026 35586
rect 135662 35534 135714 35586
rect 137006 35534 137058 35586
rect 141598 35534 141650 35586
rect 143950 35534 144002 35586
rect 144958 35534 145010 35586
rect 20750 35422 20802 35474
rect 31278 35422 31330 35474
rect 31614 35422 31666 35474
rect 40014 35422 40066 35474
rect 40350 35422 40402 35474
rect 51662 35422 51714 35474
rect 51998 35422 52050 35474
rect 66334 35422 66386 35474
rect 66670 35422 66722 35474
rect 76302 35422 76354 35474
rect 76638 35422 76690 35474
rect 90526 35422 90578 35474
rect 92430 35422 92482 35474
rect 93998 35422 94050 35474
rect 94334 35422 94386 35474
rect 99374 35422 99426 35474
rect 99710 35422 99762 35474
rect 119870 35422 119922 35474
rect 120206 35422 120258 35474
rect 142270 35422 142322 35474
rect 19624 35254 19676 35306
rect 19728 35254 19780 35306
rect 19832 35254 19884 35306
rect 56444 35254 56496 35306
rect 56548 35254 56600 35306
rect 56652 35254 56704 35306
rect 93264 35254 93316 35306
rect 93368 35254 93420 35306
rect 93472 35254 93524 35306
rect 130084 35254 130136 35306
rect 130188 35254 130240 35306
rect 130292 35254 130344 35306
rect 30046 35086 30098 35138
rect 49758 35086 49810 35138
rect 52670 35086 52722 35138
rect 68126 35086 68178 35138
rect 120654 35086 120706 35138
rect 123118 35086 123170 35138
rect 130734 35086 130786 35138
rect 138798 35086 138850 35138
rect 5854 34974 5906 35026
rect 6974 34974 7026 35026
rect 7534 34974 7586 35026
rect 8430 34974 8482 35026
rect 10334 34974 10386 35026
rect 12910 34974 12962 35026
rect 13918 34974 13970 35026
rect 17166 34974 17218 35026
rect 21870 34974 21922 35026
rect 23774 34974 23826 35026
rect 26126 34974 26178 35026
rect 28142 34974 28194 35026
rect 32398 34974 32450 35026
rect 34190 34974 34242 35026
rect 35982 34974 36034 35026
rect 38446 34974 38498 35026
rect 39902 34974 39954 35026
rect 41806 34974 41858 35026
rect 43486 34974 43538 35026
rect 50878 34974 50930 35026
rect 54238 34974 54290 35026
rect 57710 34974 57762 35026
rect 59502 34974 59554 35026
rect 62974 34974 63026 35026
rect 70366 34974 70418 35026
rect 72270 34974 72322 35026
rect 74510 34974 74562 35026
rect 80782 34974 80834 35026
rect 82574 34974 82626 35026
rect 85934 34974 85986 35026
rect 87950 34974 88002 35026
rect 88958 34974 89010 35026
rect 93326 34974 93378 35026
rect 95790 34974 95842 35026
rect 97582 34974 97634 35026
rect 99262 34974 99314 35026
rect 100270 34974 100322 35026
rect 101838 34974 101890 35026
rect 103630 34974 103682 35026
rect 109790 34974 109842 35026
rect 111582 34974 111634 35026
rect 115502 34974 115554 35026
rect 118414 34974 118466 35026
rect 121550 34974 121602 35026
rect 124014 34974 124066 35026
rect 125134 34974 125186 35026
rect 127710 34974 127762 35026
rect 133646 34974 133698 35026
rect 136334 34974 136386 35026
rect 140142 34974 140194 35026
rect 141710 34974 141762 35026
rect 142830 34974 142882 35026
rect 143278 34974 143330 35026
rect 143726 34974 143778 35026
rect 6750 34862 6802 34914
rect 7534 34862 7586 34914
rect 11230 34862 11282 34914
rect 15038 34862 15090 34914
rect 18286 34862 18338 34914
rect 19070 34862 19122 34914
rect 19742 34862 19794 34914
rect 22878 34862 22930 34914
rect 24894 34862 24946 34914
rect 27022 34862 27074 34914
rect 28814 34862 28866 34914
rect 30830 34862 30882 34914
rect 33182 34862 33234 34914
rect 34974 34862 35026 34914
rect 36766 34862 36818 34914
rect 41022 34862 41074 34914
rect 42814 34862 42866 34914
rect 44606 34862 44658 34914
rect 45614 34862 45666 34914
rect 46398 34862 46450 34914
rect 47854 34862 47906 34914
rect 51998 34862 52050 34914
rect 55358 34862 55410 34914
rect 58718 34862 58770 34914
rect 60622 34862 60674 34914
rect 61742 34862 61794 34914
rect 62190 34862 62242 34914
rect 64094 34862 64146 34914
rect 64878 34862 64930 34914
rect 65550 34862 65602 34914
rect 71486 34862 71538 34914
rect 73278 34862 73330 34914
rect 73838 34862 73890 34914
rect 75742 34862 75794 34914
rect 76190 34862 76242 34914
rect 77422 34862 77474 34914
rect 80110 34862 80162 34914
rect 82014 34862 82066 34914
rect 85262 34862 85314 34914
rect 87278 34862 87330 34914
rect 89966 34862 90018 34914
rect 90414 34862 90466 34914
rect 94222 34862 94274 34914
rect 95118 34862 95170 34914
rect 96798 34862 96850 34914
rect 98590 34862 98642 34914
rect 101166 34862 101218 34914
rect 102958 34862 103010 34914
rect 104862 34862 104914 34914
rect 105422 34862 105474 34914
rect 106878 34862 106930 34914
rect 109230 34862 109282 34914
rect 110910 34862 110962 34914
rect 113822 34862 113874 34914
rect 114830 34862 114882 34914
rect 117742 34862 117794 34914
rect 119982 34862 120034 34914
rect 122670 34862 122722 34914
rect 126030 34862 126082 34914
rect 126814 34862 126866 34914
rect 128830 34862 128882 34914
rect 130062 34862 130114 34914
rect 132974 34862 133026 34914
rect 135662 34862 135714 34914
rect 141150 34862 141202 34914
rect 9326 34750 9378 34802
rect 9662 34750 9714 34802
rect 16158 34750 16210 34802
rect 18958 34750 19010 34802
rect 30606 34750 30658 34802
rect 37662 34750 37714 34802
rect 38222 34750 38274 34802
rect 47070 34750 47122 34802
rect 47518 34750 47570 34802
rect 48974 34750 49026 34802
rect 49534 34750 49586 34802
rect 52558 34750 52610 34802
rect 56702 34750 56754 34802
rect 57038 34750 57090 34802
rect 64766 34750 64818 34802
rect 67342 34750 67394 34802
rect 67902 34750 67954 34802
rect 78206 34750 78258 34802
rect 78542 34750 78594 34802
rect 79438 34750 79490 34802
rect 84030 34750 84082 34802
rect 84366 34750 84418 34802
rect 90526 34750 90578 34802
rect 92094 34750 92146 34802
rect 106094 34750 106146 34802
rect 106654 34750 106706 34802
rect 107886 34750 107938 34802
rect 113150 34750 113202 34802
rect 113486 34750 113538 34802
rect 119870 34750 119922 34802
rect 122334 34750 122386 34802
rect 129950 34750 130002 34802
rect 131742 34750 131794 34802
rect 132078 34750 132130 34802
rect 134766 34750 134818 34802
rect 138014 34750 138066 34802
rect 138574 34750 138626 34802
rect 139694 34750 139746 34802
rect 144734 34750 144786 34802
rect 15598 34638 15650 34690
rect 16494 34638 16546 34690
rect 20078 34638 20130 34690
rect 20750 34638 20802 34690
rect 29710 34638 29762 34690
rect 31502 34638 31554 34690
rect 38782 34638 38834 34690
rect 46062 34638 46114 34690
rect 48190 34638 48242 34690
rect 50094 34638 50146 34690
rect 53678 34638 53730 34690
rect 56254 34638 56306 34690
rect 65886 34638 65938 34690
rect 66782 34638 66834 34690
rect 68462 34638 68514 34690
rect 69470 34638 69522 34690
rect 77646 34638 77698 34690
rect 78990 34638 79042 34690
rect 89630 34638 89682 34690
rect 91310 34638 91362 34690
rect 92430 34638 92482 34690
rect 107214 34638 107266 34690
rect 108222 34638 108274 34690
rect 114158 34638 114210 34690
rect 116958 34638 117010 34690
rect 120990 34638 121042 34690
rect 123454 34638 123506 34690
rect 129278 34638 129330 34690
rect 131070 34638 131122 34690
rect 135102 34638 135154 34690
rect 137342 34638 137394 34690
rect 139134 34638 139186 34690
rect 145630 34638 145682 34690
rect 38034 34470 38086 34522
rect 38138 34470 38190 34522
rect 38242 34470 38294 34522
rect 74854 34470 74906 34522
rect 74958 34470 75010 34522
rect 75062 34470 75114 34522
rect 111674 34470 111726 34522
rect 111778 34470 111830 34522
rect 111882 34470 111934 34522
rect 148494 34470 148546 34522
rect 148598 34470 148650 34522
rect 148702 34470 148754 34522
rect 7758 34302 7810 34354
rect 10894 34302 10946 34354
rect 11678 34302 11730 34354
rect 14254 34302 14306 34354
rect 15934 34302 15986 34354
rect 16718 34302 16770 34354
rect 17838 34302 17890 34354
rect 18286 34302 18338 34354
rect 19182 34302 19234 34354
rect 22766 34302 22818 34354
rect 23662 34302 23714 34354
rect 24446 34302 24498 34354
rect 27358 34302 27410 34354
rect 27918 34302 27970 34354
rect 28366 34302 28418 34354
rect 29374 34302 29426 34354
rect 33518 34302 33570 34354
rect 33966 34302 34018 34354
rect 35646 34302 35698 34354
rect 36654 34302 36706 34354
rect 37102 34302 37154 34354
rect 39902 34302 39954 34354
rect 43150 34302 43202 34354
rect 44270 34302 44322 34354
rect 44718 34302 44770 34354
rect 48750 34302 48802 34354
rect 56366 34302 56418 34354
rect 56814 34302 56866 34354
rect 57486 34302 57538 34354
rect 72718 34302 72770 34354
rect 73726 34302 73778 34354
rect 74174 34302 74226 34354
rect 74734 34302 74786 34354
rect 75630 34302 75682 34354
rect 76302 34302 76354 34354
rect 78654 34302 78706 34354
rect 85486 34302 85538 34354
rect 87614 34302 87666 34354
rect 93774 34302 93826 34354
rect 95566 34302 95618 34354
rect 96462 34302 96514 34354
rect 98926 34302 98978 34354
rect 101502 34302 101554 34354
rect 102062 34302 102114 34354
rect 109230 34302 109282 34354
rect 109566 34302 109618 34354
rect 110126 34302 110178 34354
rect 110910 34302 110962 34354
rect 111358 34302 111410 34354
rect 115054 34302 115106 34354
rect 117742 34302 117794 34354
rect 125246 34302 125298 34354
rect 125694 34302 125746 34354
rect 126254 34302 126306 34354
rect 129390 34302 129442 34354
rect 132638 34302 132690 34354
rect 133870 34302 133922 34354
rect 134318 34302 134370 34354
rect 134766 34302 134818 34354
rect 135326 34302 135378 34354
rect 136334 34302 136386 34354
rect 11230 34190 11282 34242
rect 16270 34190 16322 34242
rect 18622 34190 18674 34242
rect 21870 34190 21922 34242
rect 22206 34190 22258 34242
rect 23214 34190 23266 34242
rect 26126 34190 26178 34242
rect 29934 34190 29986 34242
rect 31726 34190 31778 34242
rect 38110 34190 38162 34242
rect 40462 34190 40514 34242
rect 40798 34190 40850 34242
rect 42478 34190 42530 34242
rect 45278 34190 45330 34242
rect 47070 34190 47122 34242
rect 49646 34190 49698 34242
rect 51438 34190 51490 34242
rect 52446 34190 52498 34242
rect 54126 34190 54178 34242
rect 58942 34190 58994 34242
rect 60734 34190 60786 34242
rect 61406 34190 61458 34242
rect 63646 34190 63698 34242
rect 64542 34190 64594 34242
rect 68126 34190 68178 34242
rect 68574 34190 68626 34242
rect 69918 34190 69970 34242
rect 76862 34190 76914 34242
rect 77198 34190 77250 34242
rect 88622 34190 88674 34242
rect 89294 34190 89346 34242
rect 90414 34190 90466 34242
rect 102622 34190 102674 34242
rect 113374 34190 113426 34242
rect 113822 34190 113874 34242
rect 121438 34190 121490 34242
rect 130622 34190 130674 34242
rect 137006 34190 137058 34242
rect 138350 34190 138402 34242
rect 143054 34190 143106 34242
rect 8094 34078 8146 34130
rect 14590 34078 14642 34130
rect 19406 34078 19458 34130
rect 20190 34078 20242 34130
rect 25790 34078 25842 34130
rect 31054 34078 31106 34130
rect 32846 34078 32898 34130
rect 37438 34078 37490 34130
rect 39118 34078 39170 34130
rect 42142 34078 42194 34130
rect 46286 34078 46338 34130
rect 48190 34078 48242 34130
rect 50766 34078 50818 34130
rect 51774 34078 51826 34130
rect 53566 34078 53618 34130
rect 54462 34078 54514 34130
rect 57822 34078 57874 34130
rect 58606 34078 58658 34130
rect 60398 34078 60450 34130
rect 62526 34078 62578 34130
rect 63310 34078 63362 34130
rect 64318 34078 64370 34130
rect 67342 34078 67394 34130
rect 68798 34078 68850 34130
rect 71038 34078 71090 34130
rect 73502 34078 73554 34130
rect 81902 34078 81954 34130
rect 83806 34078 83858 34130
rect 89630 34078 89682 34130
rect 90302 34078 90354 34130
rect 92206 34078 92258 34130
rect 97246 34078 97298 34130
rect 100046 34078 100098 34130
rect 103182 34078 103234 34130
rect 105198 34078 105250 34130
rect 106990 34078 107042 34130
rect 110462 34078 110514 34130
rect 111918 34078 111970 34130
rect 114158 34078 114210 34130
rect 115950 34078 116002 34130
rect 118078 34078 118130 34130
rect 120094 34078 120146 34130
rect 122558 34078 122610 34130
rect 123118 34078 123170 34130
rect 130510 34078 130562 34130
rect 131294 34078 131346 34130
rect 132302 34078 132354 34130
rect 133534 34078 133586 34130
rect 138574 34078 138626 34130
rect 139022 34078 139074 34130
rect 140030 34078 140082 34130
rect 142942 34078 142994 34130
rect 143726 34078 143778 34130
rect 145070 34078 145122 34130
rect 7198 33966 7250 34018
rect 8542 33966 8594 34018
rect 9886 33966 9938 34018
rect 15038 33966 15090 34018
rect 20750 33966 20802 34018
rect 24894 33966 24946 34018
rect 28814 33966 28866 34018
rect 31054 33966 31106 34018
rect 31390 33966 31442 34018
rect 34526 33966 34578 34018
rect 35198 33966 35250 34018
rect 36094 33966 36146 34018
rect 41582 33966 41634 34018
rect 54910 33966 54962 34018
rect 59502 33966 59554 34018
rect 59838 33966 59890 34018
rect 65662 33966 65714 34018
rect 66446 33966 66498 34018
rect 71038 33966 71090 34018
rect 69134 33854 69186 33906
rect 71486 33966 71538 34018
rect 71934 33966 71986 34018
rect 75070 33966 75122 34018
rect 77646 33966 77698 34018
rect 78206 33966 78258 34018
rect 79102 33966 79154 34018
rect 79774 33966 79826 34018
rect 80558 33966 80610 34018
rect 81454 33966 81506 34018
rect 82686 33966 82738 34018
rect 84590 33966 84642 34018
rect 85150 33966 85202 34018
rect 87054 33966 87106 34018
rect 88174 33966 88226 34018
rect 91086 33966 91138 34018
rect 92766 33966 92818 34018
rect 94222 33966 94274 34018
rect 94782 33966 94834 34018
rect 95118 33966 95170 34018
rect 96014 33966 96066 34018
rect 97918 33966 97970 34018
rect 100494 33966 100546 34018
rect 103854 33966 103906 34018
rect 105870 33966 105922 34018
rect 107662 33966 107714 34018
rect 108670 33966 108722 34018
rect 112478 33966 112530 34018
rect 116622 33966 116674 34018
rect 118526 33966 118578 34018
rect 119310 33966 119362 34018
rect 123790 33966 123842 34018
rect 124798 33966 124850 34018
rect 126590 33966 126642 34018
rect 128942 33966 128994 34018
rect 129950 33966 130002 34018
rect 137342 33966 137394 34018
rect 140702 33966 140754 34018
rect 141822 33966 141874 34018
rect 142382 33966 142434 34018
rect 145630 33966 145682 34018
rect 71486 33854 71538 33906
rect 78206 33854 78258 33906
rect 78766 33854 78818 33906
rect 91422 33854 91474 33906
rect 96014 33854 96066 33906
rect 96686 33854 96738 33906
rect 114494 33854 114546 33906
rect 131630 33854 131682 33906
rect 139358 33854 139410 33906
rect 144062 33854 144114 33906
rect 19624 33686 19676 33738
rect 19728 33686 19780 33738
rect 19832 33686 19884 33738
rect 56444 33686 56496 33738
rect 56548 33686 56600 33738
rect 56652 33686 56704 33738
rect 93264 33686 93316 33738
rect 93368 33686 93420 33738
rect 93472 33686 93524 33738
rect 130084 33686 130136 33738
rect 130188 33686 130240 33738
rect 130292 33686 130344 33738
rect 45502 33518 45554 33570
rect 46174 33518 46226 33570
rect 69246 33518 69298 33570
rect 69806 33518 69858 33570
rect 104862 33518 104914 33570
rect 105422 33518 105474 33570
rect 121774 33518 121826 33570
rect 122222 33518 122274 33570
rect 14926 33406 14978 33458
rect 18846 33406 18898 33458
rect 19742 33406 19794 33458
rect 21534 33406 21586 33458
rect 25230 33406 25282 33458
rect 29486 33406 29538 33458
rect 31838 33406 31890 33458
rect 32622 33406 32674 33458
rect 33406 33406 33458 33458
rect 36878 33406 36930 33458
rect 41806 33406 41858 33458
rect 42142 33406 42194 33458
rect 42702 33406 42754 33458
rect 45502 33406 45554 33458
rect 47518 33406 47570 33458
rect 50766 33406 50818 33458
rect 52446 33406 52498 33458
rect 53454 33406 53506 33458
rect 53902 33406 53954 33458
rect 57150 33406 57202 33458
rect 58270 33406 58322 33458
rect 59166 33406 59218 33458
rect 59614 33406 59666 33458
rect 60174 33406 60226 33458
rect 60734 33406 60786 33458
rect 64990 33406 65042 33458
rect 67118 33406 67170 33458
rect 67678 33406 67730 33458
rect 68126 33406 68178 33458
rect 69358 33406 69410 33458
rect 69806 33406 69858 33458
rect 71374 33406 71426 33458
rect 73726 33406 73778 33458
rect 76078 33406 76130 33458
rect 76526 33406 76578 33458
rect 77982 33406 78034 33458
rect 82574 33406 82626 33458
rect 89070 33406 89122 33458
rect 90750 33406 90802 33458
rect 91870 33406 91922 33458
rect 93214 33406 93266 33458
rect 94110 33406 94162 33458
rect 95230 33406 95282 33458
rect 98254 33406 98306 33458
rect 98590 33406 98642 33458
rect 101054 33406 101106 33458
rect 101614 33406 101666 33458
rect 102734 33406 102786 33458
rect 104078 33406 104130 33458
rect 104974 33406 105026 33458
rect 105422 33406 105474 33458
rect 105870 33406 105922 33458
rect 106318 33406 106370 33458
rect 107662 33406 107714 33458
rect 107998 33406 108050 33458
rect 111918 33406 111970 33458
rect 113038 33406 113090 33458
rect 114606 33406 114658 33458
rect 117070 33406 117122 33458
rect 120654 33406 120706 33458
rect 121102 33406 121154 33458
rect 122894 33406 122946 33458
rect 128606 33406 128658 33458
rect 130510 33406 130562 33458
rect 133198 33406 133250 33458
rect 136782 33406 136834 33458
rect 138126 33406 138178 33458
rect 139582 33406 139634 33458
rect 140142 33406 140194 33458
rect 142718 33406 142770 33458
rect 45950 33294 46002 33346
rect 50206 33294 50258 33346
rect 61518 33294 61570 33346
rect 62078 33294 62130 33346
rect 62638 33294 62690 33346
rect 65886 33294 65938 33346
rect 88174 33294 88226 33346
rect 89966 33294 90018 33346
rect 106766 33294 106818 33346
rect 112366 33294 112418 33346
rect 129614 33294 129666 33346
rect 131406 33294 131458 33346
rect 131966 33294 132018 33346
rect 137454 33294 137506 33346
rect 19406 33182 19458 33234
rect 38670 33182 38722 33234
rect 39902 33182 39954 33234
rect 40462 33182 40514 33234
rect 46398 33182 46450 33234
rect 46734 33182 46786 33234
rect 47966 33182 48018 33234
rect 48302 33182 48354 33234
rect 48862 33182 48914 33234
rect 49198 33182 49250 33234
rect 51214 33182 51266 33234
rect 51550 33182 51602 33234
rect 62974 33182 63026 33234
rect 99822 33182 99874 33234
rect 100270 33182 100322 33234
rect 118414 33182 118466 33234
rect 118750 33182 118802 33234
rect 119646 33182 119698 33234
rect 123902 33182 123954 33234
rect 20526 33070 20578 33122
rect 22094 33070 22146 33122
rect 30830 33070 30882 33122
rect 31390 33070 31442 33122
rect 32286 33070 32338 33122
rect 37662 33070 37714 33122
rect 38110 33070 38162 33122
rect 39006 33070 39058 33122
rect 39566 33070 39618 33122
rect 40798 33070 40850 33122
rect 41246 33070 41298 33122
rect 49870 33070 49922 33122
rect 51998 33070 52050 33122
rect 57822 33070 57874 33122
rect 63422 33070 63474 33122
rect 63870 33070 63922 33122
rect 64318 33070 64370 33122
rect 66670 33070 66722 33122
rect 70814 33070 70866 33122
rect 87726 33070 87778 33122
rect 92206 33070 92258 33122
rect 93550 33070 93602 33122
rect 94782 33070 94834 33122
rect 97246 33070 97298 33122
rect 99486 33070 99538 33122
rect 114046 33070 114098 33122
rect 117406 33070 117458 33122
rect 117854 33070 117906 33122
rect 119310 33070 119362 33122
rect 120094 33070 120146 33122
rect 121774 33070 121826 33122
rect 122110 33070 122162 33122
rect 123566 33070 123618 33122
rect 124910 33070 124962 33122
rect 38034 32902 38086 32954
rect 38138 32902 38190 32954
rect 38242 32902 38294 32954
rect 74854 32902 74906 32954
rect 74958 32902 75010 32954
rect 75062 32902 75114 32954
rect 111674 32902 111726 32954
rect 111778 32902 111830 32954
rect 111882 32902 111934 32954
rect 148494 32902 148546 32954
rect 148598 32902 148650 32954
rect 148702 32902 148754 32954
rect 39454 32734 39506 32786
rect 40126 32734 40178 32786
rect 41582 32734 41634 32786
rect 42030 32734 42082 32786
rect 46510 32734 46562 32786
rect 46958 32734 47010 32786
rect 47630 32734 47682 32786
rect 48190 32734 48242 32786
rect 49422 32734 49474 32786
rect 49870 32734 49922 32786
rect 50542 32734 50594 32786
rect 62302 32734 62354 32786
rect 62862 32734 62914 32786
rect 63198 32734 63250 32786
rect 63982 32734 64034 32786
rect 65438 32734 65490 32786
rect 65774 32734 65826 32786
rect 66222 32734 66274 32786
rect 67118 32734 67170 32786
rect 89294 32734 89346 32786
rect 90750 32734 90802 32786
rect 91198 32734 91250 32786
rect 92430 32734 92482 32786
rect 119758 32734 119810 32786
rect 130958 32734 131010 32786
rect 131406 32734 131458 32786
rect 38446 32622 38498 32674
rect 91646 32622 91698 32674
rect 39006 32510 39058 32562
rect 40798 32510 40850 32562
rect 48526 32510 48578 32562
rect 91982 32510 92034 32562
rect 51326 32398 51378 32450
rect 52558 32398 52610 32450
rect 61854 32398 61906 32450
rect 64430 32398 64482 32450
rect 89742 32398 89794 32450
rect 92990 32398 93042 32450
rect 118750 32398 118802 32450
rect 119310 32398 119362 32450
rect 19624 32118 19676 32170
rect 19728 32118 19780 32170
rect 19832 32118 19884 32170
rect 56444 32118 56496 32170
rect 56548 32118 56600 32170
rect 56652 32118 56704 32170
rect 93264 32118 93316 32170
rect 93368 32118 93420 32170
rect 93472 32118 93524 32170
rect 130084 32118 130136 32170
rect 130188 32118 130240 32170
rect 130292 32118 130344 32170
rect 64878 31838 64930 31890
rect 48974 31502 49026 31554
rect 38034 31334 38086 31386
rect 38138 31334 38190 31386
rect 38242 31334 38294 31386
rect 74854 31334 74906 31386
rect 74958 31334 75010 31386
rect 75062 31334 75114 31386
rect 111674 31334 111726 31386
rect 111778 31334 111830 31386
rect 111882 31334 111934 31386
rect 148494 31334 148546 31386
rect 148598 31334 148650 31386
rect 148702 31334 148754 31386
rect 19624 30550 19676 30602
rect 19728 30550 19780 30602
rect 19832 30550 19884 30602
rect 56444 30550 56496 30602
rect 56548 30550 56600 30602
rect 56652 30550 56704 30602
rect 93264 30550 93316 30602
rect 93368 30550 93420 30602
rect 93472 30550 93524 30602
rect 130084 30550 130136 30602
rect 130188 30550 130240 30602
rect 130292 30550 130344 30602
rect 38034 29766 38086 29818
rect 38138 29766 38190 29818
rect 38242 29766 38294 29818
rect 74854 29766 74906 29818
rect 74958 29766 75010 29818
rect 75062 29766 75114 29818
rect 111674 29766 111726 29818
rect 111778 29766 111830 29818
rect 111882 29766 111934 29818
rect 148494 29766 148546 29818
rect 148598 29766 148650 29818
rect 148702 29766 148754 29818
rect 19624 28982 19676 29034
rect 19728 28982 19780 29034
rect 19832 28982 19884 29034
rect 56444 28982 56496 29034
rect 56548 28982 56600 29034
rect 56652 28982 56704 29034
rect 93264 28982 93316 29034
rect 93368 28982 93420 29034
rect 93472 28982 93524 29034
rect 130084 28982 130136 29034
rect 130188 28982 130240 29034
rect 130292 28982 130344 29034
rect 38034 28198 38086 28250
rect 38138 28198 38190 28250
rect 38242 28198 38294 28250
rect 74854 28198 74906 28250
rect 74958 28198 75010 28250
rect 75062 28198 75114 28250
rect 111674 28198 111726 28250
rect 111778 28198 111830 28250
rect 111882 28198 111934 28250
rect 148494 28198 148546 28250
rect 148598 28198 148650 28250
rect 148702 28198 148754 28250
rect 19624 27414 19676 27466
rect 19728 27414 19780 27466
rect 19832 27414 19884 27466
rect 56444 27414 56496 27466
rect 56548 27414 56600 27466
rect 56652 27414 56704 27466
rect 93264 27414 93316 27466
rect 93368 27414 93420 27466
rect 93472 27414 93524 27466
rect 130084 27414 130136 27466
rect 130188 27414 130240 27466
rect 130292 27414 130344 27466
rect 38034 26630 38086 26682
rect 38138 26630 38190 26682
rect 38242 26630 38294 26682
rect 74854 26630 74906 26682
rect 74958 26630 75010 26682
rect 75062 26630 75114 26682
rect 111674 26630 111726 26682
rect 111778 26630 111830 26682
rect 111882 26630 111934 26682
rect 148494 26630 148546 26682
rect 148598 26630 148650 26682
rect 148702 26630 148754 26682
rect 19624 25846 19676 25898
rect 19728 25846 19780 25898
rect 19832 25846 19884 25898
rect 56444 25846 56496 25898
rect 56548 25846 56600 25898
rect 56652 25846 56704 25898
rect 93264 25846 93316 25898
rect 93368 25846 93420 25898
rect 93472 25846 93524 25898
rect 130084 25846 130136 25898
rect 130188 25846 130240 25898
rect 130292 25846 130344 25898
rect 38034 25062 38086 25114
rect 38138 25062 38190 25114
rect 38242 25062 38294 25114
rect 74854 25062 74906 25114
rect 74958 25062 75010 25114
rect 75062 25062 75114 25114
rect 111674 25062 111726 25114
rect 111778 25062 111830 25114
rect 111882 25062 111934 25114
rect 148494 25062 148546 25114
rect 148598 25062 148650 25114
rect 148702 25062 148754 25114
rect 19624 24278 19676 24330
rect 19728 24278 19780 24330
rect 19832 24278 19884 24330
rect 56444 24278 56496 24330
rect 56548 24278 56600 24330
rect 56652 24278 56704 24330
rect 93264 24278 93316 24330
rect 93368 24278 93420 24330
rect 93472 24278 93524 24330
rect 130084 24278 130136 24330
rect 130188 24278 130240 24330
rect 130292 24278 130344 24330
rect 38034 23494 38086 23546
rect 38138 23494 38190 23546
rect 38242 23494 38294 23546
rect 74854 23494 74906 23546
rect 74958 23494 75010 23546
rect 75062 23494 75114 23546
rect 111674 23494 111726 23546
rect 111778 23494 111830 23546
rect 111882 23494 111934 23546
rect 148494 23494 148546 23546
rect 148598 23494 148650 23546
rect 148702 23494 148754 23546
rect 19624 22710 19676 22762
rect 19728 22710 19780 22762
rect 19832 22710 19884 22762
rect 56444 22710 56496 22762
rect 56548 22710 56600 22762
rect 56652 22710 56704 22762
rect 93264 22710 93316 22762
rect 93368 22710 93420 22762
rect 93472 22710 93524 22762
rect 130084 22710 130136 22762
rect 130188 22710 130240 22762
rect 130292 22710 130344 22762
rect 38034 21926 38086 21978
rect 38138 21926 38190 21978
rect 38242 21926 38294 21978
rect 74854 21926 74906 21978
rect 74958 21926 75010 21978
rect 75062 21926 75114 21978
rect 111674 21926 111726 21978
rect 111778 21926 111830 21978
rect 111882 21926 111934 21978
rect 148494 21926 148546 21978
rect 148598 21926 148650 21978
rect 148702 21926 148754 21978
rect 19624 21142 19676 21194
rect 19728 21142 19780 21194
rect 19832 21142 19884 21194
rect 56444 21142 56496 21194
rect 56548 21142 56600 21194
rect 56652 21142 56704 21194
rect 93264 21142 93316 21194
rect 93368 21142 93420 21194
rect 93472 21142 93524 21194
rect 130084 21142 130136 21194
rect 130188 21142 130240 21194
rect 130292 21142 130344 21194
rect 38034 20358 38086 20410
rect 38138 20358 38190 20410
rect 38242 20358 38294 20410
rect 74854 20358 74906 20410
rect 74958 20358 75010 20410
rect 75062 20358 75114 20410
rect 111674 20358 111726 20410
rect 111778 20358 111830 20410
rect 111882 20358 111934 20410
rect 148494 20358 148546 20410
rect 148598 20358 148650 20410
rect 148702 20358 148754 20410
rect 19624 19574 19676 19626
rect 19728 19574 19780 19626
rect 19832 19574 19884 19626
rect 56444 19574 56496 19626
rect 56548 19574 56600 19626
rect 56652 19574 56704 19626
rect 93264 19574 93316 19626
rect 93368 19574 93420 19626
rect 93472 19574 93524 19626
rect 130084 19574 130136 19626
rect 130188 19574 130240 19626
rect 130292 19574 130344 19626
rect 38034 18790 38086 18842
rect 38138 18790 38190 18842
rect 38242 18790 38294 18842
rect 74854 18790 74906 18842
rect 74958 18790 75010 18842
rect 75062 18790 75114 18842
rect 111674 18790 111726 18842
rect 111778 18790 111830 18842
rect 111882 18790 111934 18842
rect 148494 18790 148546 18842
rect 148598 18790 148650 18842
rect 148702 18790 148754 18842
rect 19624 18006 19676 18058
rect 19728 18006 19780 18058
rect 19832 18006 19884 18058
rect 56444 18006 56496 18058
rect 56548 18006 56600 18058
rect 56652 18006 56704 18058
rect 93264 18006 93316 18058
rect 93368 18006 93420 18058
rect 93472 18006 93524 18058
rect 130084 18006 130136 18058
rect 130188 18006 130240 18058
rect 130292 18006 130344 18058
rect 38034 17222 38086 17274
rect 38138 17222 38190 17274
rect 38242 17222 38294 17274
rect 74854 17222 74906 17274
rect 74958 17222 75010 17274
rect 75062 17222 75114 17274
rect 111674 17222 111726 17274
rect 111778 17222 111830 17274
rect 111882 17222 111934 17274
rect 148494 17222 148546 17274
rect 148598 17222 148650 17274
rect 148702 17222 148754 17274
rect 19624 16438 19676 16490
rect 19728 16438 19780 16490
rect 19832 16438 19884 16490
rect 56444 16438 56496 16490
rect 56548 16438 56600 16490
rect 56652 16438 56704 16490
rect 93264 16438 93316 16490
rect 93368 16438 93420 16490
rect 93472 16438 93524 16490
rect 130084 16438 130136 16490
rect 130188 16438 130240 16490
rect 130292 16438 130344 16490
rect 38034 15654 38086 15706
rect 38138 15654 38190 15706
rect 38242 15654 38294 15706
rect 74854 15654 74906 15706
rect 74958 15654 75010 15706
rect 75062 15654 75114 15706
rect 111674 15654 111726 15706
rect 111778 15654 111830 15706
rect 111882 15654 111934 15706
rect 148494 15654 148546 15706
rect 148598 15654 148650 15706
rect 148702 15654 148754 15706
rect 19624 14870 19676 14922
rect 19728 14870 19780 14922
rect 19832 14870 19884 14922
rect 56444 14870 56496 14922
rect 56548 14870 56600 14922
rect 56652 14870 56704 14922
rect 93264 14870 93316 14922
rect 93368 14870 93420 14922
rect 93472 14870 93524 14922
rect 130084 14870 130136 14922
rect 130188 14870 130240 14922
rect 130292 14870 130344 14922
rect 38034 14086 38086 14138
rect 38138 14086 38190 14138
rect 38242 14086 38294 14138
rect 74854 14086 74906 14138
rect 74958 14086 75010 14138
rect 75062 14086 75114 14138
rect 111674 14086 111726 14138
rect 111778 14086 111830 14138
rect 111882 14086 111934 14138
rect 148494 14086 148546 14138
rect 148598 14086 148650 14138
rect 148702 14086 148754 14138
rect 19624 13302 19676 13354
rect 19728 13302 19780 13354
rect 19832 13302 19884 13354
rect 56444 13302 56496 13354
rect 56548 13302 56600 13354
rect 56652 13302 56704 13354
rect 93264 13302 93316 13354
rect 93368 13302 93420 13354
rect 93472 13302 93524 13354
rect 130084 13302 130136 13354
rect 130188 13302 130240 13354
rect 130292 13302 130344 13354
rect 38034 12518 38086 12570
rect 38138 12518 38190 12570
rect 38242 12518 38294 12570
rect 74854 12518 74906 12570
rect 74958 12518 75010 12570
rect 75062 12518 75114 12570
rect 111674 12518 111726 12570
rect 111778 12518 111830 12570
rect 111882 12518 111934 12570
rect 148494 12518 148546 12570
rect 148598 12518 148650 12570
rect 148702 12518 148754 12570
rect 19624 11734 19676 11786
rect 19728 11734 19780 11786
rect 19832 11734 19884 11786
rect 56444 11734 56496 11786
rect 56548 11734 56600 11786
rect 56652 11734 56704 11786
rect 93264 11734 93316 11786
rect 93368 11734 93420 11786
rect 93472 11734 93524 11786
rect 130084 11734 130136 11786
rect 130188 11734 130240 11786
rect 130292 11734 130344 11786
rect 38034 10950 38086 11002
rect 38138 10950 38190 11002
rect 38242 10950 38294 11002
rect 74854 10950 74906 11002
rect 74958 10950 75010 11002
rect 75062 10950 75114 11002
rect 111674 10950 111726 11002
rect 111778 10950 111830 11002
rect 111882 10950 111934 11002
rect 148494 10950 148546 11002
rect 148598 10950 148650 11002
rect 148702 10950 148754 11002
rect 19624 10166 19676 10218
rect 19728 10166 19780 10218
rect 19832 10166 19884 10218
rect 56444 10166 56496 10218
rect 56548 10166 56600 10218
rect 56652 10166 56704 10218
rect 93264 10166 93316 10218
rect 93368 10166 93420 10218
rect 93472 10166 93524 10218
rect 130084 10166 130136 10218
rect 130188 10166 130240 10218
rect 130292 10166 130344 10218
rect 128718 9886 128770 9938
rect 129278 9550 129330 9602
rect 38034 9382 38086 9434
rect 38138 9382 38190 9434
rect 38242 9382 38294 9434
rect 74854 9382 74906 9434
rect 74958 9382 75010 9434
rect 75062 9382 75114 9434
rect 111674 9382 111726 9434
rect 111778 9382 111830 9434
rect 111882 9382 111934 9434
rect 148494 9382 148546 9434
rect 148598 9382 148650 9434
rect 148702 9382 148754 9434
rect 67230 9214 67282 9266
rect 64654 9102 64706 9154
rect 66110 9102 66162 9154
rect 66446 9102 66498 9154
rect 128270 9102 128322 9154
rect 130174 9102 130226 9154
rect 131294 9102 131346 9154
rect 65886 8990 65938 9042
rect 128046 8990 128098 9042
rect 129166 8990 129218 9042
rect 129502 8990 129554 9042
rect 130286 8990 130338 9042
rect 130846 8990 130898 9042
rect 64318 8878 64370 8930
rect 65550 8766 65602 8818
rect 19624 8598 19676 8650
rect 19728 8598 19780 8650
rect 19832 8598 19884 8650
rect 56444 8598 56496 8650
rect 56548 8598 56600 8650
rect 56652 8598 56704 8650
rect 93264 8598 93316 8650
rect 93368 8598 93420 8650
rect 93472 8598 93524 8650
rect 130084 8598 130136 8650
rect 130188 8598 130240 8650
rect 130292 8598 130344 8650
rect 67678 8318 67730 8370
rect 63646 8206 63698 8258
rect 64206 8206 64258 8258
rect 119198 8206 119250 8258
rect 120542 8206 120594 8258
rect 131294 8206 131346 8258
rect 131854 8206 131906 8258
rect 118302 8094 118354 8146
rect 119422 8094 119474 8146
rect 119870 8094 119922 8146
rect 127374 8094 127426 8146
rect 63198 7982 63250 8034
rect 66782 7982 66834 8034
rect 67342 7982 67394 8034
rect 68238 7982 68290 8034
rect 88958 7982 89010 8034
rect 118862 7982 118914 8034
rect 121102 7982 121154 8034
rect 121438 7982 121490 8034
rect 126814 7982 126866 8034
rect 127710 7982 127762 8034
rect 128158 7982 128210 8034
rect 128942 7982 128994 8034
rect 132302 7982 132354 8034
rect 132862 7982 132914 8034
rect 38034 7814 38086 7866
rect 38138 7814 38190 7866
rect 38242 7814 38294 7866
rect 74854 7814 74906 7866
rect 74958 7814 75010 7866
rect 75062 7814 75114 7866
rect 111674 7814 111726 7866
rect 111778 7814 111830 7866
rect 111882 7814 111934 7866
rect 148494 7814 148546 7866
rect 148598 7814 148650 7866
rect 148702 7814 148754 7866
rect 19966 7646 20018 7698
rect 78318 7646 78370 7698
rect 90862 7646 90914 7698
rect 113598 7646 113650 7698
rect 123342 7646 123394 7698
rect 126366 7646 126418 7698
rect 127038 7646 127090 7698
rect 19070 7534 19122 7586
rect 28366 7534 28418 7586
rect 50318 7534 50370 7586
rect 62526 7534 62578 7586
rect 62862 7534 62914 7586
rect 63086 7534 63138 7586
rect 63310 7534 63362 7586
rect 63534 7534 63586 7586
rect 66110 7534 66162 7586
rect 66446 7534 66498 7586
rect 67790 7534 67842 7586
rect 76302 7534 76354 7586
rect 76750 7534 76802 7586
rect 99598 7534 99650 7586
rect 118078 7534 118130 7586
rect 119646 7534 119698 7586
rect 120206 7534 120258 7586
rect 121326 7534 121378 7586
rect 126030 7534 126082 7586
rect 128046 7534 128098 7586
rect 129726 7534 129778 7586
rect 141486 7534 141538 7586
rect 142382 7534 142434 7586
rect 18510 7422 18562 7474
rect 18958 7422 19010 7474
rect 28702 7422 28754 7474
rect 48750 7422 48802 7474
rect 50542 7422 50594 7474
rect 51550 7422 51602 7474
rect 63870 7422 63922 7474
rect 65550 7422 65602 7474
rect 65886 7422 65938 7474
rect 68126 7422 68178 7474
rect 76974 7422 77026 7474
rect 88510 7422 88562 7474
rect 99262 7422 99314 7474
rect 118414 7422 118466 7474
rect 119086 7422 119138 7474
rect 119422 7422 119474 7474
rect 121214 7422 121266 7474
rect 121998 7422 122050 7474
rect 128158 7422 128210 7474
rect 132078 7422 132130 7474
rect 132638 7422 132690 7474
rect 141822 7422 141874 7474
rect 142606 7422 142658 7474
rect 20302 7310 20354 7362
rect 20750 7310 20802 7362
rect 26350 7310 26402 7362
rect 29150 7310 29202 7362
rect 39230 7310 39282 7362
rect 39790 7310 39842 7362
rect 48414 7310 48466 7362
rect 49758 7310 49810 7362
rect 51102 7310 51154 7362
rect 64654 7310 64706 7362
rect 67230 7310 67282 7362
rect 68686 7310 68738 7362
rect 69134 7310 69186 7362
rect 69470 7310 69522 7362
rect 69918 7310 69970 7362
rect 75070 7310 75122 7362
rect 75518 7310 75570 7362
rect 77870 7310 77922 7362
rect 89182 7310 89234 7362
rect 89630 7310 89682 7362
rect 90414 7310 90466 7362
rect 91422 7310 91474 7362
rect 113038 7310 113090 7362
rect 114158 7310 114210 7362
rect 115950 7310 116002 7362
rect 116734 7310 116786 7362
rect 117518 7310 117570 7362
rect 122894 7310 122946 7362
rect 133086 7310 133138 7362
rect 133534 7310 133586 7362
rect 18174 7198 18226 7250
rect 64542 7198 64594 7250
rect 77310 7198 77362 7250
rect 77646 7198 77698 7250
rect 78206 7198 78258 7250
rect 113374 7198 113426 7250
rect 114158 7198 114210 7250
rect 122334 7198 122386 7250
rect 127374 7198 127426 7250
rect 128942 7198 128994 7250
rect 19624 7030 19676 7082
rect 19728 7030 19780 7082
rect 19832 7030 19884 7082
rect 56444 7030 56496 7082
rect 56548 7030 56600 7082
rect 56652 7030 56704 7082
rect 93264 7030 93316 7082
rect 93368 7030 93420 7082
rect 93472 7030 93524 7082
rect 130084 7030 130136 7082
rect 130188 7030 130240 7082
rect 130292 7030 130344 7082
rect 27134 6862 27186 6914
rect 29710 6862 29762 6914
rect 30046 6862 30098 6914
rect 47854 6862 47906 6914
rect 50206 6862 50258 6914
rect 68126 6862 68178 6914
rect 68462 6862 68514 6914
rect 87390 6862 87442 6914
rect 89742 6862 89794 6914
rect 91198 6862 91250 6914
rect 99150 6862 99202 6914
rect 99486 6862 99538 6914
rect 126590 6862 126642 6914
rect 127374 6862 127426 6914
rect 141822 6862 141874 6914
rect 142158 6862 142210 6914
rect 39118 6750 39170 6802
rect 40126 6750 40178 6802
rect 114382 6750 114434 6802
rect 115726 6750 115778 6802
rect 7422 6638 7474 6690
rect 7870 6638 7922 6690
rect 16158 6638 16210 6690
rect 16718 6638 16770 6690
rect 20414 6638 20466 6690
rect 20862 6638 20914 6690
rect 27806 6638 27858 6690
rect 31502 6638 31554 6690
rect 49534 6638 49586 6690
rect 51214 6638 51266 6690
rect 62302 6638 62354 6690
rect 62862 6638 62914 6690
rect 71262 6638 71314 6690
rect 78206 6638 78258 6690
rect 81118 6638 81170 6690
rect 89182 6638 89234 6690
rect 91982 6638 92034 6690
rect 93102 6638 93154 6690
rect 98478 6638 98530 6690
rect 100270 6638 100322 6690
rect 101054 6638 101106 6690
rect 111582 6638 111634 6690
rect 113374 6638 113426 6690
rect 115166 6638 115218 6690
rect 117630 6638 117682 6690
rect 118302 6638 118354 6690
rect 122110 6638 122162 6690
rect 127038 6638 127090 6690
rect 128046 6638 128098 6690
rect 128382 6638 128434 6690
rect 133646 6638 133698 6690
rect 143950 6638 144002 6690
rect 10894 6526 10946 6578
rect 26126 6526 26178 6578
rect 26798 6526 26850 6578
rect 27918 6526 27970 6578
rect 28814 6526 28866 6578
rect 30270 6526 30322 6578
rect 30830 6526 30882 6578
rect 38334 6526 38386 6578
rect 38894 6526 38946 6578
rect 48078 6526 48130 6578
rect 48414 6526 48466 6578
rect 49422 6526 49474 6578
rect 50542 6526 50594 6578
rect 52110 6526 52162 6578
rect 66334 6526 66386 6578
rect 66670 6526 66722 6578
rect 67566 6526 67618 6578
rect 67902 6526 67954 6578
rect 69470 6526 69522 6578
rect 73278 6526 73330 6578
rect 77646 6526 77698 6578
rect 79998 6526 80050 6578
rect 81566 6526 81618 6578
rect 87614 6526 87666 6578
rect 88174 6526 88226 6578
rect 89070 6526 89122 6578
rect 91870 6526 91922 6578
rect 100046 6526 100098 6578
rect 112254 6526 112306 6578
rect 115054 6526 115106 6578
rect 131966 6526 132018 6578
rect 132078 6526 132130 6578
rect 133086 6526 133138 6578
rect 133758 6526 133810 6578
rect 142494 6526 142546 6578
rect 142718 6526 142770 6578
rect 10334 6414 10386 6466
rect 11230 6414 11282 6466
rect 19182 6414 19234 6466
rect 19854 6414 19906 6466
rect 21534 6414 21586 6466
rect 25790 6414 25842 6466
rect 39454 6414 39506 6466
rect 40462 6414 40514 6466
rect 47518 6414 47570 6466
rect 51550 6414 51602 6466
rect 52446 6414 52498 6466
rect 61854 6414 61906 6466
rect 65326 6414 65378 6466
rect 65886 6414 65938 6466
rect 69358 6414 69410 6466
rect 69918 6414 69970 6466
rect 70702 6414 70754 6466
rect 77310 6414 77362 6466
rect 78542 6414 78594 6466
rect 87054 6414 87106 6466
rect 90078 6414 90130 6466
rect 90862 6414 90914 6466
rect 93662 6414 93714 6466
rect 101614 6414 101666 6466
rect 110462 6414 110514 6466
rect 111022 6414 111074 6466
rect 114046 6414 114098 6466
rect 116286 6414 116338 6466
rect 117182 6414 117234 6466
rect 120542 6414 120594 6466
rect 121326 6414 121378 6466
rect 121774 6414 121826 6466
rect 127374 6414 127426 6466
rect 130958 6414 131010 6466
rect 131518 6414 131570 6466
rect 132974 6414 133026 6466
rect 134206 6414 134258 6466
rect 141262 6414 141314 6466
rect 143502 6414 143554 6466
rect 38034 6246 38086 6298
rect 38138 6246 38190 6298
rect 38242 6246 38294 6298
rect 74854 6246 74906 6298
rect 74958 6246 75010 6298
rect 75062 6246 75114 6298
rect 111674 6246 111726 6298
rect 111778 6246 111830 6298
rect 111882 6246 111934 6298
rect 148494 6246 148546 6298
rect 148598 6246 148650 6298
rect 148702 6246 148754 6298
rect 8094 6078 8146 6130
rect 11342 6078 11394 6130
rect 14926 6078 14978 6130
rect 16046 6078 16098 6130
rect 17838 6078 17890 6130
rect 20526 6078 20578 6130
rect 30942 6078 30994 6130
rect 31502 6078 31554 6130
rect 50318 6078 50370 6130
rect 51102 6078 51154 6130
rect 59950 6078 60002 6130
rect 60846 6078 60898 6130
rect 65550 6078 65602 6130
rect 70142 6078 70194 6130
rect 72158 6078 72210 6130
rect 73502 6078 73554 6130
rect 74062 6078 74114 6130
rect 75742 6078 75794 6130
rect 87390 6078 87442 6130
rect 88510 6078 88562 6130
rect 90414 6078 90466 6130
rect 101726 6078 101778 6130
rect 107886 6078 107938 6130
rect 110350 6078 110402 6130
rect 113374 6078 113426 6130
rect 117070 6078 117122 6130
rect 126478 6078 126530 6130
rect 132078 6078 132130 6130
rect 140254 6078 140306 6130
rect 143726 6078 143778 6130
rect 145294 6078 145346 6130
rect 16606 5966 16658 6018
rect 16942 5966 16994 6018
rect 18958 5966 19010 6018
rect 19518 5966 19570 6018
rect 21982 5966 22034 6018
rect 38446 5966 38498 6018
rect 39678 5966 39730 6018
rect 46622 5966 46674 6018
rect 46958 5966 47010 6018
rect 61518 5966 61570 6018
rect 71150 5966 71202 6018
rect 74734 5966 74786 6018
rect 75182 5966 75234 6018
rect 77086 5966 77138 6018
rect 86158 5966 86210 6018
rect 86494 5966 86546 6018
rect 89630 5966 89682 6018
rect 91534 5966 91586 6018
rect 91870 5966 91922 6018
rect 108558 5966 108610 6018
rect 109678 5966 109730 6018
rect 112030 5966 112082 6018
rect 112366 5966 112418 6018
rect 115054 5966 115106 6018
rect 115614 5966 115666 6018
rect 133086 5966 133138 6018
rect 134094 5966 134146 6018
rect 137902 5966 137954 6018
rect 138686 5966 138738 6018
rect 139134 5966 139186 6018
rect 142718 5966 142770 6018
rect 144846 5966 144898 6018
rect 8430 5854 8482 5906
rect 15822 5854 15874 5906
rect 18398 5854 18450 5906
rect 18734 5854 18786 5906
rect 26910 5854 26962 5906
rect 28030 5854 28082 5906
rect 28366 5854 28418 5906
rect 31838 5854 31890 5906
rect 36766 5854 36818 5906
rect 37886 5854 37938 5906
rect 38670 5854 38722 5906
rect 39454 5854 39506 5906
rect 41470 5854 41522 5906
rect 48750 5854 48802 5906
rect 49758 5854 49810 5906
rect 52894 5854 52946 5906
rect 53342 5854 53394 5906
rect 64654 5854 64706 5906
rect 66110 5854 66162 5906
rect 67006 5854 67058 5906
rect 67678 5854 67730 5906
rect 70702 5854 70754 5906
rect 75406 5854 75458 5906
rect 79326 5854 79378 5906
rect 79998 5854 80050 5906
rect 87950 5854 88002 5906
rect 89406 5854 89458 5906
rect 90974 5854 91026 5906
rect 101278 5854 101330 5906
rect 108894 5854 108946 5906
rect 109566 5854 109618 5906
rect 114270 5854 114322 5906
rect 114942 5854 114994 5906
rect 116510 5854 116562 5906
rect 119646 5854 119698 5906
rect 119982 5854 120034 5906
rect 127150 5854 127202 5906
rect 129166 5854 129218 5906
rect 129614 5854 129666 5906
rect 133310 5854 133362 5906
rect 139358 5854 139410 5906
rect 140814 5854 140866 5906
rect 141374 5854 141426 5906
rect 142606 5854 142658 5906
rect 143390 5854 143442 5906
rect 9774 5742 9826 5794
rect 10110 5742 10162 5794
rect 11902 5742 11954 5794
rect 12462 5742 12514 5794
rect 20638 5742 20690 5794
rect 21198 5742 21250 5794
rect 21534 5742 21586 5794
rect 25790 5742 25842 5794
rect 27470 5742 27522 5794
rect 35646 5742 35698 5794
rect 40238 5742 40290 5794
rect 40910 5742 40962 5794
rect 45278 5742 45330 5794
rect 47630 5742 47682 5794
rect 51774 5742 51826 5794
rect 56478 5742 56530 5794
rect 57486 5742 57538 5794
rect 60510 5742 60562 5794
rect 62638 5742 62690 5794
rect 63534 5742 63586 5794
rect 66670 5742 66722 5794
rect 71262 5742 71314 5794
rect 71710 5742 71762 5794
rect 72606 5742 72658 5794
rect 80446 5742 80498 5794
rect 92430 5742 92482 5794
rect 94894 5742 94946 5794
rect 100158 5742 100210 5794
rect 110686 5742 110738 5794
rect 111134 5742 111186 5794
rect 116174 5742 116226 5794
rect 120990 5742 121042 5794
rect 128158 5742 128210 5794
rect 134542 5742 134594 5794
rect 134990 5742 135042 5794
rect 135438 5742 135490 5794
rect 137454 5742 137506 5794
rect 141934 5742 141986 5794
rect 37550 5630 37602 5682
rect 40350 5630 40402 5682
rect 60510 5630 60562 5682
rect 61182 5630 61234 5682
rect 76302 5630 76354 5682
rect 113934 5630 113986 5682
rect 132638 5630 132690 5682
rect 133982 5630 134034 5682
rect 139694 5630 139746 5682
rect 19624 5462 19676 5514
rect 19728 5462 19780 5514
rect 19832 5462 19884 5514
rect 56444 5462 56496 5514
rect 56548 5462 56600 5514
rect 56652 5462 56704 5514
rect 93264 5462 93316 5514
rect 93368 5462 93420 5514
rect 93472 5462 93524 5514
rect 130084 5462 130136 5514
rect 130188 5462 130240 5514
rect 130292 5462 130344 5514
rect 20862 5294 20914 5346
rect 28702 5294 28754 5346
rect 31950 5294 32002 5346
rect 37438 5294 37490 5346
rect 49086 5294 49138 5346
rect 67342 5294 67394 5346
rect 67678 5294 67730 5346
rect 72942 5294 72994 5346
rect 88958 5294 89010 5346
rect 98702 5294 98754 5346
rect 115502 5294 115554 5346
rect 116286 5294 116338 5346
rect 131518 5294 131570 5346
rect 132862 5294 132914 5346
rect 138350 5294 138402 5346
rect 12686 5182 12738 5234
rect 21758 5182 21810 5234
rect 22206 5182 22258 5234
rect 35422 5182 35474 5234
rect 41694 5182 41746 5234
rect 46958 5182 47010 5234
rect 53566 5182 53618 5234
rect 54126 5182 54178 5234
rect 54462 5182 54514 5234
rect 59614 5182 59666 5234
rect 62190 5182 62242 5234
rect 89406 5182 89458 5234
rect 90078 5182 90130 5234
rect 91646 5182 91698 5234
rect 92206 5182 92258 5234
rect 93102 5182 93154 5234
rect 101950 5182 102002 5234
rect 102510 5182 102562 5234
rect 105758 5182 105810 5234
rect 116174 5182 116226 5234
rect 120990 5182 121042 5234
rect 125694 5182 125746 5234
rect 126926 5182 126978 5234
rect 132078 5182 132130 5234
rect 138014 5182 138066 5234
rect 139694 5182 139746 5234
rect 140142 5182 140194 5234
rect 140814 5182 140866 5234
rect 141374 5182 141426 5234
rect 142718 5182 142770 5234
rect 144510 5182 144562 5234
rect 145854 5182 145906 5234
rect 146526 5182 146578 5234
rect 7422 5070 7474 5122
rect 7870 5070 7922 5122
rect 10222 5070 10274 5122
rect 11678 5070 11730 5122
rect 15150 5070 15202 5122
rect 15822 5070 15874 5122
rect 16494 5070 16546 5122
rect 17166 5070 17218 5122
rect 17726 5070 17778 5122
rect 25118 5070 25170 5122
rect 25678 5070 25730 5122
rect 29486 5070 29538 5122
rect 30270 5070 30322 5122
rect 31390 5070 31442 5122
rect 32062 5070 32114 5122
rect 32510 5070 32562 5122
rect 40462 5070 40514 5122
rect 41022 5070 41074 5122
rect 41582 5070 41634 5122
rect 42254 5070 42306 5122
rect 44606 5070 44658 5122
rect 48078 5070 48130 5122
rect 48638 5070 48690 5122
rect 52222 5070 52274 5122
rect 52558 5070 52610 5122
rect 53454 5070 53506 5122
rect 60398 5070 60450 5122
rect 66670 5070 66722 5122
rect 69470 5070 69522 5122
rect 70478 5070 70530 5122
rect 76078 5070 76130 5122
rect 76638 5070 76690 5122
rect 77310 5070 77362 5122
rect 84478 5070 84530 5122
rect 85486 5070 85538 5122
rect 85934 5070 85986 5122
rect 89518 5070 89570 5122
rect 93662 5070 93714 5122
rect 95230 5070 95282 5122
rect 95566 5070 95618 5122
rect 104190 5070 104242 5122
rect 105310 5070 105362 5122
rect 108110 5070 108162 5122
rect 109230 5070 109282 5122
rect 110350 5070 110402 5122
rect 112030 5070 112082 5122
rect 112366 5070 112418 5122
rect 117182 5070 117234 5122
rect 117630 5070 117682 5122
rect 120654 5070 120706 5122
rect 125022 5070 125074 5122
rect 127374 5070 127426 5122
rect 127822 5070 127874 5122
rect 128382 5070 128434 5122
rect 131966 5070 132018 5122
rect 135886 5070 135938 5122
rect 136334 5070 136386 5122
rect 139134 5070 139186 5122
rect 141710 5070 141762 5122
rect 142270 5070 142322 5122
rect 143502 5070 143554 5122
rect 145182 5070 145234 5122
rect 11790 4958 11842 5010
rect 12238 4958 12290 5010
rect 14142 4958 14194 5010
rect 34302 4958 34354 5010
rect 36766 4958 36818 5010
rect 38222 4958 38274 5010
rect 43598 4958 43650 5010
rect 45614 4958 45666 5010
rect 49870 4958 49922 5010
rect 56478 4958 56530 5010
rect 57822 4958 57874 5010
rect 58158 4958 58210 5010
rect 67902 4958 67954 5010
rect 68238 4958 68290 5010
rect 71486 4958 71538 5010
rect 71934 4958 71986 5010
rect 82238 4958 82290 5010
rect 90750 4958 90802 5010
rect 91086 4958 91138 5010
rect 94222 4958 94274 5010
rect 94558 4958 94610 5010
rect 111022 4958 111074 5010
rect 137342 4958 137394 5010
rect 138910 4958 138962 5010
rect 145070 4958 145122 5010
rect 11118 4846 11170 4898
rect 16382 4846 16434 4898
rect 20302 4846 20354 4898
rect 21646 4846 21698 4898
rect 28142 4846 28194 4898
rect 33742 4846 33794 4898
rect 36430 4846 36482 4898
rect 48526 4846 48578 4898
rect 55918 4846 55970 4898
rect 56814 4846 56866 4898
rect 57262 4846 57314 4898
rect 58830 4846 58882 4898
rect 71150 4846 71202 4898
rect 72606 4846 72658 4898
rect 73726 4846 73778 4898
rect 88398 4846 88450 4898
rect 91758 4846 91810 4898
rect 97918 4846 97970 4898
rect 102062 4846 102114 4898
rect 108334 4846 108386 4898
rect 111358 4846 111410 4898
rect 114942 4846 114994 4898
rect 120094 4846 120146 4898
rect 130958 4846 131010 4898
rect 133422 4846 133474 4898
rect 137006 4846 137058 4898
rect 144174 4846 144226 4898
rect 38034 4678 38086 4730
rect 38138 4678 38190 4730
rect 38242 4678 38294 4730
rect 74854 4678 74906 4730
rect 74958 4678 75010 4730
rect 75062 4678 75114 4730
rect 111674 4678 111726 4730
rect 111778 4678 111830 4730
rect 111882 4678 111934 4730
rect 148494 4678 148546 4730
rect 148598 4678 148650 4730
rect 148702 4678 148754 4730
rect 12014 4510 12066 4562
rect 16046 4510 16098 4562
rect 16942 4510 16994 4562
rect 28142 4510 28194 4562
rect 38558 4510 38610 4562
rect 39118 4510 39170 4562
rect 48302 4510 48354 4562
rect 48862 4510 48914 4562
rect 51550 4510 51602 4562
rect 55022 4510 55074 4562
rect 60622 4510 60674 4562
rect 64206 4510 64258 4562
rect 64766 4510 64818 4562
rect 81230 4510 81282 4562
rect 81678 4510 81730 4562
rect 85598 4510 85650 4562
rect 86270 4510 86322 4562
rect 92094 4510 92146 4562
rect 92878 4510 92930 4562
rect 97134 4510 97186 4562
rect 97918 4510 97970 4562
rect 98366 4510 98418 4562
rect 102510 4510 102562 4562
rect 107550 4510 107602 4562
rect 111134 4510 111186 4562
rect 116174 4510 116226 4562
rect 116734 4510 116786 4562
rect 118974 4510 119026 4562
rect 124238 4510 124290 4562
rect 127822 4510 127874 4562
rect 128382 4510 128434 4562
rect 131854 4510 131906 4562
rect 134878 4510 134930 4562
rect 135886 4510 135938 4562
rect 143726 4510 143778 4562
rect 146750 4510 146802 4562
rect 7422 4398 7474 4450
rect 11006 4398 11058 4450
rect 12126 4398 12178 4450
rect 21086 4398 21138 4450
rect 22206 4398 22258 4450
rect 26238 4398 26290 4450
rect 28926 4398 28978 4450
rect 32734 4398 32786 4450
rect 33518 4398 33570 4450
rect 41694 4398 41746 4450
rect 49646 4398 49698 4450
rect 53118 4398 53170 4450
rect 57598 4398 57650 4450
rect 59502 4398 59554 4450
rect 68686 4398 68738 4450
rect 80334 4398 80386 4450
rect 86830 4398 86882 4450
rect 97806 4398 97858 4450
rect 103182 4398 103234 4450
rect 119310 4398 119362 4450
rect 119870 4398 119922 4450
rect 135214 4398 135266 4450
rect 136222 4398 136274 4450
rect 137790 4398 137842 4450
rect 141822 4398 141874 4450
rect 144062 4398 144114 4450
rect 145630 4398 145682 4450
rect 145966 4398 146018 4450
rect 5854 4286 5906 4338
rect 12910 4286 12962 4338
rect 13582 4286 13634 4338
rect 19406 4286 19458 4338
rect 35534 4286 35586 4338
rect 36094 4286 36146 4338
rect 39566 4286 39618 4338
rect 45278 4286 45330 4338
rect 45838 4286 45890 4338
rect 56478 4286 56530 4338
rect 59838 4286 59890 4338
rect 61070 4286 61122 4338
rect 61742 4286 61794 4338
rect 69246 4286 69298 4338
rect 72382 4286 72434 4338
rect 74622 4286 74674 4338
rect 75630 4286 75682 4338
rect 85150 4286 85202 4338
rect 88510 4286 88562 4338
rect 89182 4286 89234 4338
rect 89742 4286 89794 4338
rect 94558 4286 94610 4338
rect 96462 4286 96514 4338
rect 99038 4286 99090 4338
rect 99486 4286 99538 4338
rect 100046 4286 100098 4338
rect 108222 4286 108274 4338
rect 108558 4286 108610 4338
rect 112030 4286 112082 4338
rect 113038 4286 113090 4338
rect 113598 4286 113650 4338
rect 118190 4286 118242 4338
rect 119982 4286 120034 4338
rect 121102 4286 121154 4338
rect 124686 4286 124738 4338
rect 125358 4286 125410 4338
rect 129166 4286 129218 4338
rect 129614 4286 129666 4338
rect 134318 4286 134370 4338
rect 136894 4286 136946 4338
rect 145406 4286 145458 4338
rect 4734 4174 4786 4226
rect 6414 4174 6466 4226
rect 6862 4174 6914 4226
rect 8766 4174 8818 4226
rect 9998 4174 10050 4226
rect 17726 4174 17778 4226
rect 18846 4174 18898 4226
rect 20078 4174 20130 4226
rect 23550 4174 23602 4226
rect 25678 4174 25730 4226
rect 27582 4174 27634 4226
rect 28254 4174 28306 4226
rect 30270 4174 30322 4226
rect 30718 4174 30770 4226
rect 31390 4174 31442 4226
rect 40350 4174 40402 4226
rect 42814 4174 42866 4226
rect 50766 4174 50818 4226
rect 52558 4174 52610 4226
rect 54238 4174 54290 4226
rect 55582 4174 55634 4226
rect 58942 4174 58994 4226
rect 71598 4174 71650 4226
rect 73838 4174 73890 4226
rect 84030 4174 84082 4226
rect 87726 4174 87778 4226
rect 93438 4174 93490 4226
rect 95790 4174 95842 4226
rect 111694 4174 111746 4226
rect 117294 4174 117346 4226
rect 121774 4174 121826 4226
rect 133198 4174 133250 4226
rect 138910 4174 138962 4226
rect 141262 4174 141314 4226
rect 143166 4174 143218 4226
rect 147198 4174 147250 4226
rect 16606 4062 16658 4114
rect 132638 4062 132690 4114
rect 145070 4062 145122 4114
rect 19624 3894 19676 3946
rect 19728 3894 19780 3946
rect 19832 3894 19884 3946
rect 56444 3894 56496 3946
rect 56548 3894 56600 3946
rect 56652 3894 56704 3946
rect 93264 3894 93316 3946
rect 93368 3894 93420 3946
rect 93472 3894 93524 3946
rect 130084 3894 130136 3946
rect 130188 3894 130240 3946
rect 130292 3894 130344 3946
rect 9662 3726 9714 3778
rect 14366 3726 14418 3778
rect 63870 3726 63922 3778
rect 67678 3726 67730 3778
rect 68462 3726 68514 3778
rect 71710 3726 71762 3778
rect 75630 3726 75682 3778
rect 79214 3726 79266 3778
rect 80222 3726 80274 3778
rect 80782 3726 80834 3778
rect 84702 3726 84754 3778
rect 88622 3726 88674 3778
rect 92542 3726 92594 3778
rect 111694 3726 111746 3778
rect 115502 3726 115554 3778
rect 116174 3726 116226 3778
rect 119534 3726 119586 3778
rect 119758 3726 119810 3778
rect 120542 3726 120594 3778
rect 131518 3726 131570 3778
rect 132302 3726 132354 3778
rect 6974 3614 7026 3666
rect 8878 3614 8930 3666
rect 11342 3614 11394 3666
rect 13918 3614 13970 3666
rect 15262 3614 15314 3666
rect 18734 3614 18786 3666
rect 23326 3614 23378 3666
rect 28478 3614 28530 3666
rect 30046 3614 30098 3666
rect 31166 3614 31218 3666
rect 34862 3614 34914 3666
rect 39678 3614 39730 3666
rect 40238 3614 40290 3666
rect 43710 3614 43762 3666
rect 47518 3614 47570 3666
rect 51550 3614 51602 3666
rect 55694 3614 55746 3666
rect 59614 3614 59666 3666
rect 64654 3614 64706 3666
rect 68574 3614 68626 3666
rect 76302 3614 76354 3666
rect 76750 3614 76802 3666
rect 78430 3614 78482 3666
rect 79326 3614 79378 3666
rect 80334 3614 80386 3666
rect 95902 3614 95954 3666
rect 98814 3614 98866 3666
rect 102846 3614 102898 3666
rect 106654 3614 106706 3666
rect 108334 3614 108386 3666
rect 110574 3614 110626 3666
rect 113262 3614 113314 3666
rect 117182 3614 117234 3666
rect 119982 3614 120034 3666
rect 120430 3614 120482 3666
rect 121214 3614 121266 3666
rect 125134 3614 125186 3666
rect 128046 3614 128098 3666
rect 128494 3614 128546 3666
rect 129054 3614 129106 3666
rect 131630 3614 131682 3666
rect 132190 3614 132242 3666
rect 134318 3614 134370 3666
rect 135214 3614 135266 3666
rect 139022 3614 139074 3666
rect 139918 3614 139970 3666
rect 141038 3614 141090 3666
rect 144622 3614 144674 3666
rect 147534 3614 147586 3666
rect 6302 3502 6354 3554
rect 6414 3502 6466 3554
rect 6638 3502 6690 3554
rect 10222 3502 10274 3554
rect 14702 3502 14754 3554
rect 19406 3502 19458 3554
rect 29486 3502 29538 3554
rect 60846 3502 60898 3554
rect 72606 3502 72658 3554
rect 111806 3502 111858 3554
rect 112590 3502 112642 3554
rect 123230 3502 123282 3554
rect 135662 3502 135714 3554
rect 137342 3502 137394 3554
rect 140366 3502 140418 3554
rect 144062 3502 144114 3554
rect 146862 3502 146914 3554
rect 6862 3390 6914 3442
rect 7870 3390 7922 3442
rect 10110 3390 10162 3442
rect 10334 3390 10386 3442
rect 12350 3390 12402 3442
rect 14478 3390 14530 3442
rect 16270 3390 16322 3442
rect 17614 3390 17666 3442
rect 21870 3390 21922 3442
rect 22206 3390 22258 3442
rect 24110 3390 24162 3442
rect 25230 3390 25282 3442
rect 26574 3390 26626 3442
rect 27246 3390 27298 3442
rect 32286 3390 32338 3442
rect 33070 3390 33122 3442
rect 36206 3390 36258 3442
rect 36990 3390 37042 3442
rect 37774 3390 37826 3442
rect 38334 3390 38386 3442
rect 41246 3390 41298 3442
rect 41806 3390 41858 3442
rect 42366 3390 42418 3442
rect 45838 3390 45890 3442
rect 46398 3390 46450 3442
rect 48862 3390 48914 3442
rect 49198 3390 49250 3442
rect 49870 3390 49922 3442
rect 50430 3390 50482 3442
rect 53902 3390 53954 3442
rect 54462 3390 54514 3442
rect 56702 3390 56754 3442
rect 57934 3390 57986 3442
rect 58494 3390 58546 3442
rect 61742 3390 61794 3442
rect 65214 3390 65266 3442
rect 69582 3390 69634 3442
rect 73166 3390 73218 3442
rect 77310 3390 77362 3442
rect 82910 3390 82962 3442
rect 84030 3390 84082 3442
rect 86830 3390 86882 3442
rect 87950 3390 88002 3442
rect 91086 3390 91138 3442
rect 91870 3390 91922 3442
rect 94670 3390 94722 3442
rect 96238 3390 96290 3442
rect 96910 3390 96962 3442
rect 97470 3390 97522 3442
rect 100942 3390 100994 3442
rect 101502 3390 101554 3442
rect 104974 3390 105026 3442
rect 105534 3390 105586 3442
rect 108894 3390 108946 3442
rect 109454 3390 109506 3442
rect 112366 3390 112418 3442
rect 114606 3390 114658 3442
rect 115614 3390 115666 3442
rect 116286 3390 116338 3442
rect 118526 3390 118578 3442
rect 119422 3390 119474 3442
rect 122110 3390 122162 3442
rect 123678 3390 123730 3442
rect 126366 3390 126418 3442
rect 127150 3390 127202 3442
rect 130286 3390 130338 3442
rect 133310 3390 133362 3442
rect 135102 3390 135154 3442
rect 136446 3390 136498 3442
rect 138014 3390 138066 3442
rect 145630 3390 145682 3442
rect 29262 3278 29314 3330
rect 57038 3278 57090 3330
rect 143726 3278 143778 3330
rect 38034 3110 38086 3162
rect 38138 3110 38190 3162
rect 38242 3110 38294 3162
rect 74854 3110 74906 3162
rect 74958 3110 75010 3162
rect 75062 3110 75114 3162
rect 111674 3110 111726 3162
rect 111778 3110 111830 3162
rect 111882 3110 111934 3162
rect 148494 3110 148546 3162
rect 148598 3110 148650 3162
rect 148702 3110 148754 3162
<< metal2 >>
rect 4592 39200 4704 40000
rect 5488 39200 5600 40000
rect 6384 39200 6496 40000
rect 7280 39200 7392 40000
rect 8176 39200 8288 40000
rect 9072 39200 9184 40000
rect 9968 39200 10080 40000
rect 10864 39200 10976 40000
rect 11760 39200 11872 40000
rect 12656 39200 12768 40000
rect 13552 39200 13664 40000
rect 14448 39200 14560 40000
rect 15344 39200 15456 40000
rect 16240 39200 16352 40000
rect 17136 39200 17248 40000
rect 18032 39200 18144 40000
rect 18928 39200 19040 40000
rect 19824 39200 19936 40000
rect 20720 39200 20832 40000
rect 21616 39200 21728 40000
rect 22512 39200 22624 40000
rect 23408 39200 23520 40000
rect 24304 39200 24416 40000
rect 25200 39200 25312 40000
rect 26096 39200 26208 40000
rect 26992 39200 27104 40000
rect 27888 39200 28000 40000
rect 28784 39200 28896 40000
rect 29680 39200 29792 40000
rect 30576 39200 30688 40000
rect 31472 39200 31584 40000
rect 32368 39200 32480 40000
rect 33264 39200 33376 40000
rect 34160 39200 34272 40000
rect 35056 39200 35168 40000
rect 35952 39200 36064 40000
rect 36848 39200 36960 40000
rect 37744 39200 37856 40000
rect 38640 39200 38752 40000
rect 39536 39200 39648 40000
rect 40432 39200 40544 40000
rect 41328 39200 41440 40000
rect 42224 39200 42336 40000
rect 43120 39200 43232 40000
rect 44016 39200 44128 40000
rect 44912 39200 45024 40000
rect 45808 39200 45920 40000
rect 46704 39200 46816 40000
rect 47600 39200 47712 40000
rect 48496 39200 48608 40000
rect 49392 39200 49504 40000
rect 50288 39200 50400 40000
rect 51184 39200 51296 40000
rect 52080 39200 52192 40000
rect 52976 39200 53088 40000
rect 53872 39200 53984 40000
rect 54768 39200 54880 40000
rect 55664 39200 55776 40000
rect 56560 39200 56672 40000
rect 57456 39200 57568 40000
rect 58352 39200 58464 40000
rect 59248 39200 59360 40000
rect 60144 39200 60256 40000
rect 61040 39200 61152 40000
rect 61936 39200 62048 40000
rect 62832 39200 62944 40000
rect 63728 39200 63840 40000
rect 64624 39200 64736 40000
rect 65520 39200 65632 40000
rect 66416 39200 66528 40000
rect 67312 39200 67424 40000
rect 68208 39200 68320 40000
rect 69104 39200 69216 40000
rect 70000 39200 70112 40000
rect 70896 39200 71008 40000
rect 71792 39200 71904 40000
rect 72688 39200 72800 40000
rect 73052 39228 73444 39284
rect 4620 36372 4676 39200
rect 4844 36372 4900 36382
rect 4620 36370 4900 36372
rect 4620 36318 4846 36370
rect 4898 36318 4900 36370
rect 4620 36316 4900 36318
rect 4844 36306 4900 36316
rect 5516 35028 5572 39200
rect 6076 36260 6132 36270
rect 6076 36166 6132 36204
rect 6412 35586 6468 39200
rect 6412 35534 6414 35586
rect 6466 35534 6468 35586
rect 6412 35522 6468 35534
rect 6636 36482 6692 36494
rect 6636 36430 6638 36482
rect 6690 36430 6692 36482
rect 6636 36260 6692 36430
rect 5852 35028 5908 35038
rect 5516 35026 5908 35028
rect 5516 34974 5854 35026
rect 5906 34974 5908 35026
rect 5516 34972 5908 34974
rect 5852 34962 5908 34972
rect 6636 34692 6692 36204
rect 6860 36258 6916 36270
rect 6860 36206 6862 36258
rect 6914 36206 6916 36258
rect 6860 35028 6916 36206
rect 7196 35698 7252 35710
rect 7196 35646 7198 35698
rect 7250 35646 7252 35698
rect 6972 35028 7028 35038
rect 6860 35026 7028 35028
rect 6860 34974 6974 35026
rect 7026 34974 7028 35026
rect 6860 34972 7028 34974
rect 6972 34962 7028 34972
rect 6636 34626 6692 34636
rect 6748 34914 6804 34926
rect 6748 34862 6750 34914
rect 6802 34862 6804 34914
rect 6748 34020 6804 34862
rect 7196 34692 7252 35646
rect 7308 35140 7364 39200
rect 8204 37268 8260 39200
rect 7868 37212 8260 37268
rect 7868 36370 7924 37212
rect 7868 36318 7870 36370
rect 7922 36318 7924 36370
rect 7868 35924 7924 36318
rect 7868 35858 7924 35868
rect 8428 36932 8484 36942
rect 8316 35588 8372 35598
rect 8428 35588 8484 36876
rect 9100 36932 9156 39200
rect 9100 36866 9156 36876
rect 9996 36820 10052 39200
rect 9884 36764 10052 36820
rect 8316 35586 8484 35588
rect 8316 35534 8318 35586
rect 8370 35534 8484 35586
rect 8316 35532 8484 35534
rect 8876 36594 8932 36606
rect 8876 36542 8878 36594
rect 8930 36542 8932 36594
rect 8316 35522 8372 35532
rect 7308 35074 7364 35084
rect 8428 35140 8484 35150
rect 7532 35026 7588 35038
rect 7532 34974 7534 35026
rect 7586 34974 7588 35026
rect 7532 34914 7588 34974
rect 8428 35026 8484 35084
rect 8428 34974 8430 35026
rect 8482 34974 8484 35026
rect 8428 34962 8484 34974
rect 7532 34862 7534 34914
rect 7586 34862 7588 34914
rect 7532 34850 7588 34862
rect 8876 34804 8932 36542
rect 9660 35924 9716 35934
rect 9660 35830 9716 35868
rect 8988 35700 9044 35710
rect 8988 35698 9380 35700
rect 8988 35646 8990 35698
rect 9042 35646 9380 35698
rect 8988 35644 9380 35646
rect 8988 35634 9044 35644
rect 8876 34738 8932 34748
rect 9324 34802 9380 35644
rect 9884 35028 9940 36764
rect 10780 36370 10836 36382
rect 10780 36318 10782 36370
rect 10834 36318 10836 36370
rect 9996 36260 10052 36270
rect 9996 36166 10052 36204
rect 10444 36258 10500 36270
rect 10444 36206 10446 36258
rect 10498 36206 10500 36258
rect 10444 35698 10500 36206
rect 10444 35646 10446 35698
rect 10498 35646 10500 35698
rect 10444 35634 10500 35646
rect 10780 36260 10836 36318
rect 9884 34962 9940 34972
rect 10332 35028 10388 35038
rect 10332 34934 10388 34972
rect 10780 34916 10836 36204
rect 10892 35588 10948 39200
rect 11676 36372 11732 36382
rect 11788 36372 11844 39200
rect 11676 36370 11788 36372
rect 11676 36318 11678 36370
rect 11730 36318 11788 36370
rect 11676 36316 11788 36318
rect 11676 36306 11732 36316
rect 11788 36240 11844 36316
rect 11004 35588 11060 35598
rect 10892 35586 11060 35588
rect 10892 35534 11006 35586
rect 11058 35534 11060 35586
rect 10892 35532 11060 35534
rect 11004 35522 11060 35532
rect 12684 35586 12740 39200
rect 12796 36594 12852 36606
rect 12796 36542 12798 36594
rect 12850 36542 12852 36594
rect 12796 35812 12852 36542
rect 13580 36484 13636 39200
rect 13916 36596 13972 36606
rect 13916 36502 13972 36540
rect 13580 36428 13860 36484
rect 12796 35746 12852 35756
rect 12908 36372 12964 36382
rect 12684 35534 12686 35586
rect 12738 35534 12740 35586
rect 12684 35522 12740 35534
rect 11676 35028 11732 35038
rect 11228 34916 11284 34926
rect 10780 34850 10836 34860
rect 10892 34914 11284 34916
rect 10892 34862 11230 34914
rect 11282 34862 11284 34914
rect 10892 34860 11284 34862
rect 9324 34750 9326 34802
rect 9378 34750 9380 34802
rect 9324 34738 9380 34750
rect 9660 34802 9716 34814
rect 9660 34750 9662 34802
rect 9714 34750 9716 34802
rect 7196 34636 7812 34692
rect 7756 34354 7812 34636
rect 7756 34302 7758 34354
rect 7810 34302 7812 34354
rect 7756 34290 7812 34302
rect 8092 34130 8148 34142
rect 8092 34078 8094 34130
rect 8146 34078 8148 34130
rect 7196 34020 7252 34030
rect 6748 34018 7252 34020
rect 6748 33966 7198 34018
rect 7250 33966 7252 34018
rect 6748 33964 7252 33966
rect 7196 31892 7252 33964
rect 8092 33908 8148 34078
rect 8092 33842 8148 33852
rect 8540 34018 8596 34030
rect 8540 33966 8542 34018
rect 8594 33966 8596 34018
rect 8540 33908 8596 33966
rect 9660 34020 9716 34750
rect 10892 34354 10948 34860
rect 11228 34850 11284 34860
rect 11676 34356 11732 34972
rect 12908 35026 12964 36316
rect 13356 35698 13412 35710
rect 13356 35646 13358 35698
rect 13410 35646 13412 35698
rect 13356 35364 13412 35646
rect 13356 35298 13412 35308
rect 12908 34974 12910 35026
rect 12962 34974 12964 35026
rect 12908 34962 12964 34974
rect 13804 35028 13860 36428
rect 14364 36258 14420 36270
rect 14364 36206 14366 36258
rect 14418 36206 14420 36258
rect 14140 35700 14196 35710
rect 14364 35700 14420 36206
rect 14140 35698 14420 35700
rect 14140 35646 14142 35698
rect 14194 35646 14420 35698
rect 14140 35644 14420 35646
rect 14140 35634 14196 35644
rect 14476 35588 14532 39200
rect 15372 36596 15428 39200
rect 14700 36370 14756 36382
rect 14700 36318 14702 36370
rect 14754 36318 14756 36370
rect 14588 35588 14644 35598
rect 14476 35586 14644 35588
rect 14476 35534 14590 35586
rect 14642 35534 14644 35586
rect 14476 35532 14644 35534
rect 14588 35522 14644 35532
rect 14252 35364 14308 35374
rect 13916 35028 13972 35038
rect 13804 35026 13972 35028
rect 13804 34974 13918 35026
rect 13970 34974 13972 35026
rect 13804 34972 13972 34974
rect 13916 34962 13972 34972
rect 10892 34302 10894 34354
rect 10946 34302 10948 34354
rect 10892 34290 10948 34302
rect 11228 34354 11732 34356
rect 11228 34302 11678 34354
rect 11730 34302 11732 34354
rect 11228 34300 11732 34302
rect 11228 34242 11284 34300
rect 11676 34290 11732 34300
rect 14252 34354 14308 35308
rect 14700 34580 14756 36318
rect 15372 36370 15428 36540
rect 15372 36318 15374 36370
rect 15426 36318 15428 36370
rect 15372 36306 15428 36318
rect 16268 35586 16324 39200
rect 16268 35534 16270 35586
rect 16322 35534 16324 35586
rect 16268 35522 16324 35534
rect 16604 37044 16660 37054
rect 15036 34914 15092 34926
rect 15036 34862 15038 34914
rect 15090 34862 15092 34914
rect 14924 34580 14980 34590
rect 14700 34524 14924 34580
rect 14252 34302 14254 34354
rect 14306 34302 14308 34354
rect 14252 34290 14308 34302
rect 11228 34190 11230 34242
rect 11282 34190 11284 34242
rect 11228 34178 11284 34190
rect 14588 34130 14644 34142
rect 14588 34078 14590 34130
rect 14642 34078 14644 34130
rect 9884 34020 9940 34030
rect 9660 34018 9940 34020
rect 9660 33966 9886 34018
rect 9938 33966 9940 34018
rect 9660 33964 9940 33966
rect 8540 33842 8596 33852
rect 9884 32676 9940 33964
rect 14588 34020 14644 34078
rect 14588 33954 14644 33964
rect 14924 33458 14980 34524
rect 15036 34356 15092 34862
rect 16156 34802 16212 34814
rect 16156 34750 16158 34802
rect 16210 34750 16212 34802
rect 15036 34290 15092 34300
rect 15596 34692 15652 34702
rect 15036 34020 15092 34030
rect 15036 33926 15092 33964
rect 14924 33406 14926 33458
rect 14978 33406 14980 33458
rect 14924 33394 14980 33406
rect 9884 32610 9940 32620
rect 11676 32676 11732 32686
rect 7196 31826 7252 31836
rect 11676 6804 11732 32620
rect 15596 8428 15652 34636
rect 16156 34692 16212 34750
rect 16156 34626 16212 34636
rect 16492 34692 16548 34702
rect 16492 34598 16548 34636
rect 15932 34356 15988 34366
rect 16604 34356 16660 36988
rect 16716 36596 16772 36606
rect 16716 36594 16884 36596
rect 16716 36542 16718 36594
rect 16770 36542 16884 36594
rect 16716 36540 16884 36542
rect 16716 36530 16772 36540
rect 16828 34468 16884 36540
rect 16828 34402 16884 34412
rect 16940 35698 16996 35710
rect 16940 35646 16942 35698
rect 16994 35646 16996 35698
rect 16716 34356 16772 34366
rect 15932 34262 15988 34300
rect 16268 34354 16772 34356
rect 16268 34302 16718 34354
rect 16770 34302 16772 34354
rect 16268 34300 16772 34302
rect 16268 34242 16324 34300
rect 16716 34290 16772 34300
rect 16940 34356 16996 35646
rect 17164 35026 17220 39200
rect 18060 36484 18116 39200
rect 17724 36428 18116 36484
rect 18956 36484 19012 39200
rect 19852 37044 19908 39200
rect 19852 36988 20020 37044
rect 19622 36876 19886 36886
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19622 36810 19886 36820
rect 18956 36428 19348 36484
rect 17724 35812 17780 36428
rect 18284 36372 18340 36382
rect 18172 36370 18340 36372
rect 18172 36318 18286 36370
rect 18338 36318 18340 36370
rect 18172 36316 18340 36318
rect 17836 36260 17892 36270
rect 18172 36260 18228 36316
rect 18284 36306 18340 36316
rect 19292 36370 19348 36428
rect 19292 36318 19294 36370
rect 19346 36318 19348 36370
rect 17836 36258 18228 36260
rect 17836 36206 17838 36258
rect 17890 36206 18228 36258
rect 17836 36204 18228 36206
rect 17836 36194 17892 36204
rect 17836 35812 17892 35822
rect 17724 35810 17892 35812
rect 17724 35758 17838 35810
rect 17890 35758 17892 35810
rect 17724 35756 17892 35758
rect 17836 35746 17892 35756
rect 17164 34974 17166 35026
rect 17218 34974 17220 35026
rect 17164 34962 17220 34974
rect 16940 34290 16996 34300
rect 17836 34804 17892 34814
rect 17836 34354 17892 34748
rect 17836 34302 17838 34354
rect 17890 34302 17892 34354
rect 17836 34290 17892 34302
rect 16268 34190 16270 34242
rect 16322 34190 16324 34242
rect 16268 34178 16324 34190
rect 18172 33236 18228 36204
rect 18620 36260 18676 36270
rect 18620 36166 18676 36204
rect 18284 36036 18340 36046
rect 18284 34914 18340 35980
rect 18956 35700 19012 35710
rect 18956 35698 19236 35700
rect 18956 35646 18958 35698
rect 19010 35646 19236 35698
rect 18956 35644 19236 35646
rect 18956 35634 19012 35644
rect 19068 35476 19124 35486
rect 18284 34862 18286 34914
rect 18338 34862 18340 34914
rect 18284 34850 18340 34862
rect 18620 35140 18676 35150
rect 18396 34692 18452 34702
rect 18284 34356 18340 34366
rect 18284 34262 18340 34300
rect 18172 33170 18228 33180
rect 18396 29652 18452 34636
rect 18620 34242 18676 35084
rect 19068 34914 19124 35420
rect 19068 34862 19070 34914
rect 19122 34862 19124 34914
rect 18956 34804 19012 34814
rect 18956 34710 19012 34748
rect 18620 34190 18622 34242
rect 18674 34190 18676 34242
rect 18620 33460 18676 34190
rect 18844 33460 18900 33470
rect 18620 33458 18900 33460
rect 18620 33406 18846 33458
rect 18898 33406 18900 33458
rect 18620 33404 18900 33406
rect 18844 33394 18900 33404
rect 19068 33012 19124 34862
rect 19180 34354 19236 35644
rect 19180 34302 19182 34354
rect 19234 34302 19236 34354
rect 19180 34290 19236 34302
rect 19292 33236 19348 36318
rect 19740 35812 19796 35822
rect 19740 35718 19796 35756
rect 19628 35698 19684 35710
rect 19628 35646 19630 35698
rect 19682 35646 19684 35698
rect 19628 35476 19684 35646
rect 19628 35410 19684 35420
rect 19622 35308 19886 35318
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19622 35242 19886 35252
rect 19740 34914 19796 34926
rect 19740 34862 19742 34914
rect 19794 34862 19796 34914
rect 19740 34692 19796 34862
rect 19740 34626 19796 34636
rect 19852 34916 19908 34926
rect 19852 34468 19908 34860
rect 19404 34130 19460 34142
rect 19404 34078 19406 34130
rect 19458 34078 19460 34130
rect 19404 33460 19460 34078
rect 19852 34020 19908 34412
rect 19964 34244 20020 36988
rect 20636 36594 20692 36606
rect 20636 36542 20638 36594
rect 20690 36542 20692 36594
rect 20636 36484 20692 36542
rect 20636 36418 20692 36428
rect 20188 36260 20244 36270
rect 19964 34178 20020 34188
rect 20076 34690 20132 34702
rect 20076 34638 20078 34690
rect 20130 34638 20132 34690
rect 19852 33964 20020 34020
rect 19622 33740 19886 33750
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19622 33674 19886 33684
rect 19740 33460 19796 33470
rect 19404 33458 19796 33460
rect 19404 33406 19742 33458
rect 19794 33406 19796 33458
rect 19404 33404 19796 33406
rect 19404 33236 19460 33246
rect 19292 33234 19460 33236
rect 19292 33182 19406 33234
rect 19458 33182 19460 33234
rect 19292 33180 19460 33182
rect 19404 33170 19460 33180
rect 19740 33124 19796 33404
rect 19740 33058 19796 33068
rect 19068 32946 19124 32956
rect 19622 32172 19886 32182
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19622 32106 19886 32116
rect 19622 30604 19886 30614
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19622 30538 19886 30548
rect 18396 29586 18452 29596
rect 19622 29036 19886 29046
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19622 28970 19886 28980
rect 19622 27468 19886 27478
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19622 27402 19886 27412
rect 18508 26068 18564 26078
rect 15260 8372 15652 8428
rect 17948 17668 18004 17678
rect 15148 7588 15204 7598
rect 11676 6738 11732 6748
rect 14924 7476 14980 7486
rect 7420 6690 7476 6702
rect 7420 6638 7422 6690
rect 7474 6638 7476 6690
rect 7420 6468 7476 6638
rect 7868 6692 7924 6702
rect 7868 6690 8148 6692
rect 7868 6638 7870 6690
rect 7922 6638 8148 6690
rect 7868 6636 8148 6638
rect 7868 6626 7924 6636
rect 7420 5122 7476 6412
rect 8092 6130 8148 6636
rect 10892 6580 10948 6590
rect 10892 6486 10948 6524
rect 13580 6580 13636 6590
rect 8092 6078 8094 6130
rect 8146 6078 8148 6130
rect 8092 6066 8148 6078
rect 10332 6466 10388 6478
rect 10332 6414 10334 6466
rect 10386 6414 10388 6466
rect 8428 5908 8484 5918
rect 8428 5906 9716 5908
rect 8428 5854 8430 5906
rect 8482 5854 9716 5906
rect 8428 5852 9716 5854
rect 8428 5842 8484 5852
rect 7420 5070 7422 5122
rect 7474 5070 7476 5122
rect 7420 5058 7476 5070
rect 7868 5122 7924 5134
rect 7868 5070 7870 5122
rect 7922 5070 7924 5122
rect 6860 4452 6916 4462
rect 5852 4338 5908 4350
rect 5852 4286 5854 4338
rect 5906 4286 5908 4338
rect 4732 4228 4788 4238
rect 4396 4226 4788 4228
rect 4396 4174 4734 4226
rect 4786 4174 4788 4226
rect 4396 4172 4788 4174
rect 4396 800 4452 4172
rect 4732 4162 4788 4172
rect 5852 4004 5908 4286
rect 5852 3938 5908 3948
rect 6412 4226 6468 4238
rect 6412 4174 6414 4226
rect 6466 4174 6468 4226
rect 6412 4004 6468 4174
rect 6412 3938 6468 3948
rect 6636 4228 6692 4238
rect 6860 4228 6916 4396
rect 7420 4452 7476 4462
rect 7420 4358 7476 4396
rect 6412 3668 6468 3678
rect 6300 3556 6356 3566
rect 6300 3462 6356 3500
rect 6412 3554 6468 3612
rect 6412 3502 6414 3554
rect 6466 3502 6468 3554
rect 6412 3490 6468 3502
rect 6636 3554 6692 4172
rect 6636 3502 6638 3554
rect 6690 3502 6692 3554
rect 6636 3490 6692 3502
rect 6748 4226 6916 4228
rect 6748 4174 6862 4226
rect 6914 4174 6916 4226
rect 6748 4172 6916 4174
rect 6748 2772 6804 4172
rect 6860 4162 6916 4172
rect 6972 3668 7028 3678
rect 7868 3668 7924 5070
rect 6972 3666 7924 3668
rect 6972 3614 6974 3666
rect 7026 3614 7924 3666
rect 6972 3612 7924 3614
rect 8316 4564 8372 4574
rect 6972 3602 7028 3612
rect 6860 3444 6916 3454
rect 6860 3350 6916 3388
rect 7868 3444 7924 3454
rect 8316 3444 8372 4508
rect 8764 4228 8820 4238
rect 8764 4134 8820 4172
rect 9660 3778 9716 5852
rect 9660 3726 9662 3778
rect 9714 3726 9716 3778
rect 9660 3714 9716 3726
rect 9772 5794 9828 5806
rect 9772 5742 9774 5794
rect 9826 5742 9828 5794
rect 9772 4452 9828 5742
rect 10108 5794 10164 5806
rect 10108 5742 10110 5794
rect 10162 5742 10164 5794
rect 10108 4564 10164 5742
rect 10220 5124 10276 5134
rect 10220 5030 10276 5068
rect 10108 4498 10164 4508
rect 10332 4564 10388 6414
rect 11228 6468 11284 6478
rect 11228 6132 11284 6412
rect 12908 6468 12964 6478
rect 11340 6132 11396 6142
rect 11228 6130 11396 6132
rect 11228 6078 11342 6130
rect 11394 6078 11396 6130
rect 11228 6076 11396 6078
rect 11340 6066 11396 6076
rect 11900 5794 11956 5806
rect 11900 5742 11902 5794
rect 11954 5742 11956 5794
rect 11676 5124 11732 5134
rect 11676 5030 11732 5068
rect 11788 5012 11844 5022
rect 11788 4918 11844 4956
rect 11116 4900 11172 4910
rect 11116 4806 11172 4844
rect 10332 4498 10388 4508
rect 8876 3666 8932 3678
rect 8876 3614 8878 3666
rect 8930 3614 8932 3666
rect 7868 3442 8484 3444
rect 7868 3390 7870 3442
rect 7922 3390 8484 3442
rect 7868 3388 8484 3390
rect 7868 3378 7924 3388
rect 6748 2716 7140 2772
rect 5740 2548 5796 2558
rect 5740 800 5796 2492
rect 7084 800 7140 2716
rect 8428 800 8484 3388
rect 8876 3220 8932 3614
rect 8876 3154 8932 3164
rect 9772 800 9828 4396
rect 11004 4452 11060 4462
rect 11004 4358 11060 4396
rect 9996 4228 10052 4238
rect 9884 4226 10052 4228
rect 9884 4174 9998 4226
rect 10050 4174 10052 4226
rect 9884 4172 10052 4174
rect 9884 3444 9940 4172
rect 9996 4162 10052 4172
rect 10220 4228 10276 4238
rect 10220 3554 10276 4172
rect 11340 3668 11396 3678
rect 11340 3574 11396 3612
rect 10220 3502 10222 3554
rect 10274 3502 10276 3554
rect 10220 3490 10276 3502
rect 11116 3556 11172 3566
rect 9884 3378 9940 3388
rect 10108 3444 10164 3454
rect 10108 3350 10164 3388
rect 10332 3442 10388 3454
rect 10332 3390 10334 3442
rect 10386 3390 10388 3442
rect 10332 3332 10388 3390
rect 10332 3266 10388 3276
rect 11116 800 11172 3500
rect 11900 3556 11956 5742
rect 12460 5794 12516 5806
rect 12460 5742 12462 5794
rect 12514 5742 12516 5794
rect 12236 5012 12292 5022
rect 12012 4564 12068 4574
rect 12012 4470 12068 4508
rect 12124 4452 12180 4462
rect 12236 4452 12292 4956
rect 12460 5012 12516 5742
rect 12684 5236 12740 5246
rect 12684 5142 12740 5180
rect 12460 4946 12516 4956
rect 12124 4450 12292 4452
rect 12124 4398 12126 4450
rect 12178 4398 12292 4450
rect 12124 4396 12292 4398
rect 12124 4386 12180 4396
rect 12908 4338 12964 6412
rect 12908 4286 12910 4338
rect 12962 4286 12964 4338
rect 12908 4274 12964 4286
rect 13580 5236 13636 6524
rect 14924 6132 14980 7420
rect 13580 4338 13636 5180
rect 14700 6130 14980 6132
rect 14700 6078 14926 6130
rect 14978 6078 14980 6130
rect 14700 6076 14980 6078
rect 14140 5012 14196 5022
rect 13580 4286 13582 4338
rect 13634 4286 13636 4338
rect 13580 4274 13636 4286
rect 13804 5010 14196 5012
rect 13804 4958 14142 5010
rect 14194 4958 14196 5010
rect 13804 4956 14196 4958
rect 11900 3490 11956 3500
rect 12348 3556 12404 3566
rect 12348 3442 12404 3500
rect 12348 3390 12350 3442
rect 12402 3390 12404 3442
rect 12348 3378 12404 3390
rect 13804 800 13860 4956
rect 14140 4946 14196 4956
rect 13916 4004 13972 4014
rect 13916 3666 13972 3948
rect 14364 4004 14420 4014
rect 14364 3778 14420 3948
rect 14364 3726 14366 3778
rect 14418 3726 14420 3778
rect 14364 3714 14420 3726
rect 13916 3614 13918 3666
rect 13970 3614 13972 3666
rect 13916 3602 13972 3614
rect 14700 3554 14756 6076
rect 14924 6066 14980 6076
rect 15148 5122 15204 7532
rect 15148 5070 15150 5122
rect 15202 5070 15204 5122
rect 15148 5058 15204 5070
rect 15260 3666 15316 8372
rect 16604 7252 16660 7262
rect 16156 6690 16212 6702
rect 16156 6638 16158 6690
rect 16210 6638 16212 6690
rect 16156 6468 16212 6638
rect 16156 6402 16212 6412
rect 16044 6132 16100 6142
rect 16044 6038 16100 6076
rect 16604 6018 16660 7196
rect 16716 6690 16772 6702
rect 16716 6638 16718 6690
rect 16770 6638 16772 6690
rect 16716 6132 16772 6638
rect 16716 6066 16772 6076
rect 16828 6468 16884 6478
rect 16604 5966 16606 6018
rect 16658 5966 16660 6018
rect 16604 5954 16660 5966
rect 15820 5908 15876 5918
rect 15820 5814 15876 5852
rect 15820 5122 15876 5134
rect 15820 5070 15822 5122
rect 15874 5070 15876 5122
rect 15820 5012 15876 5070
rect 15820 4946 15876 4956
rect 16492 5122 16548 5134
rect 16492 5070 16494 5122
rect 16546 5070 16548 5122
rect 16492 5012 16548 5070
rect 16380 4900 16436 4910
rect 16044 4898 16436 4900
rect 16044 4846 16382 4898
rect 16434 4846 16436 4898
rect 16044 4844 16436 4846
rect 16044 4562 16100 4844
rect 16380 4834 16436 4844
rect 16044 4510 16046 4562
rect 16098 4510 16100 4562
rect 16044 4498 16100 4510
rect 16492 3780 16548 4956
rect 16828 5124 16884 6412
rect 17836 6132 17892 6142
rect 17836 6038 17892 6076
rect 16940 6018 16996 6030
rect 16940 5966 16942 6018
rect 16994 5966 16996 6018
rect 16940 5572 16996 5966
rect 16940 5516 17332 5572
rect 17164 5124 17220 5134
rect 16828 5122 17220 5124
rect 16828 5070 17166 5122
rect 17218 5070 17220 5122
rect 16828 5068 17220 5070
rect 17276 5124 17332 5516
rect 17724 5124 17780 5134
rect 17276 5122 17780 5124
rect 17276 5070 17726 5122
rect 17778 5070 17780 5122
rect 17276 5068 17780 5070
rect 16828 4564 16884 5068
rect 17164 5058 17220 5068
rect 17724 5058 17780 5068
rect 17948 4900 18004 17612
rect 18508 7700 18564 26012
rect 19622 25900 19886 25910
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19622 25834 19886 25844
rect 19622 24332 19886 24342
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19622 24266 19886 24276
rect 19622 22764 19886 22774
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19622 22698 19886 22708
rect 19622 21196 19886 21206
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19622 21130 19886 21140
rect 19964 20188 20020 33964
rect 20076 26068 20132 34638
rect 20188 34130 20244 36204
rect 20748 36148 20804 39200
rect 21420 36372 21476 36382
rect 21420 36278 21476 36316
rect 20636 36092 20804 36148
rect 20412 35700 20468 35710
rect 20412 35606 20468 35644
rect 20636 35140 20692 36092
rect 21420 35924 21476 35934
rect 21420 35830 21476 35868
rect 21644 35812 21700 39200
rect 22204 36372 22260 36382
rect 22540 36372 22596 39200
rect 22260 36316 22372 36372
rect 21868 36258 21924 36270
rect 21868 36206 21870 36258
rect 21922 36206 21924 36258
rect 22204 36240 22260 36316
rect 21868 36036 21924 36206
rect 21868 35970 21924 35980
rect 21980 35812 22036 35822
rect 21644 35810 22036 35812
rect 21644 35758 21982 35810
rect 22034 35758 22036 35810
rect 21644 35756 22036 35758
rect 21980 35746 22036 35756
rect 20748 35476 20804 35486
rect 20748 35474 21364 35476
rect 20748 35422 20750 35474
rect 20802 35422 21364 35474
rect 20748 35420 21364 35422
rect 20748 35410 20804 35420
rect 20636 35074 20692 35084
rect 20748 34692 20804 34702
rect 20748 34598 20804 34636
rect 20188 34078 20190 34130
rect 20242 34078 20244 34130
rect 20188 34066 20244 34078
rect 20748 34244 20804 34254
rect 20748 34018 20804 34188
rect 20748 33966 20750 34018
rect 20802 33966 20804 34018
rect 20748 33954 20804 33966
rect 20524 33122 20580 33134
rect 20524 33070 20526 33122
rect 20578 33070 20580 33122
rect 20524 33012 20580 33070
rect 20524 32946 20580 32956
rect 20076 26002 20132 26012
rect 19964 20132 20132 20188
rect 19622 19628 19886 19638
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19622 19562 19886 19572
rect 19622 18060 19886 18070
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19622 17994 19886 18004
rect 19622 16492 19886 16502
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19622 16426 19886 16436
rect 19622 14924 19886 14934
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19622 14858 19886 14868
rect 19622 13356 19886 13366
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19622 13290 19886 13300
rect 19622 11788 19886 11798
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19622 11722 19886 11732
rect 19622 10220 19886 10230
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19622 10154 19886 10164
rect 19622 8652 19886 8662
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19622 8586 19886 8596
rect 18508 7474 18564 7644
rect 19964 7700 20020 7710
rect 19964 7606 20020 7644
rect 19068 7588 19124 7598
rect 18508 7422 18510 7474
rect 18562 7422 18564 7474
rect 18508 7410 18564 7422
rect 18956 7474 19012 7486
rect 18956 7422 18958 7474
rect 19010 7422 19012 7474
rect 18172 7252 18228 7262
rect 18172 7158 18228 7196
rect 18620 6804 18676 6814
rect 18396 5908 18452 5918
rect 18396 5814 18452 5852
rect 17948 4834 18004 4844
rect 16940 4564 16996 4574
rect 16828 4562 16996 4564
rect 16828 4510 16942 4562
rect 16994 4510 16996 4562
rect 16828 4508 16996 4510
rect 16940 4498 16996 4508
rect 17724 4228 17780 4238
rect 17612 4226 17780 4228
rect 17612 4174 17726 4226
rect 17778 4174 17780 4226
rect 17612 4172 17780 4174
rect 16604 4114 16660 4126
rect 16604 4062 16606 4114
rect 16658 4062 16660 4114
rect 16604 4004 16660 4062
rect 16604 3938 16660 3948
rect 16492 3714 16548 3724
rect 15260 3614 15262 3666
rect 15314 3614 15316 3666
rect 15260 3602 15316 3614
rect 14700 3502 14702 3554
rect 14754 3502 14756 3554
rect 14700 3490 14756 3502
rect 14476 3444 14532 3454
rect 14476 3350 14532 3388
rect 15148 3444 15204 3454
rect 15148 800 15204 3388
rect 16268 3444 16324 3454
rect 16268 3350 16324 3388
rect 16492 3444 16548 3454
rect 16492 800 16548 3388
rect 17612 3444 17668 4172
rect 17724 4162 17780 4172
rect 18620 3668 18676 6748
rect 18956 6692 19012 7422
rect 19068 6804 19124 7532
rect 19622 7084 19886 7094
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19622 7018 19886 7028
rect 19068 6738 19124 6748
rect 18956 6132 19012 6636
rect 18732 6020 18788 6030
rect 18732 5906 18788 5964
rect 18956 6018 19012 6076
rect 19180 6466 19236 6478
rect 19180 6414 19182 6466
rect 19234 6414 19236 6466
rect 19180 6132 19236 6414
rect 19180 6066 19236 6076
rect 19852 6466 19908 6478
rect 19852 6414 19854 6466
rect 19906 6414 19908 6466
rect 18956 5966 18958 6018
rect 19010 5966 19012 6018
rect 18956 5954 19012 5966
rect 19516 6020 19572 6030
rect 19852 6020 19908 6414
rect 19516 6018 19908 6020
rect 19516 5966 19518 6018
rect 19570 5966 19908 6018
rect 19516 5964 19908 5966
rect 18732 5854 18734 5906
rect 18786 5854 18788 5906
rect 18732 5842 18788 5854
rect 19516 5684 19572 5964
rect 19404 5628 19572 5684
rect 19404 4338 19460 5628
rect 19622 5516 19886 5526
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19622 5450 19886 5460
rect 19404 4286 19406 4338
rect 19458 4286 19460 4338
rect 19404 4274 19460 4286
rect 18844 4228 18900 4238
rect 18844 4226 19236 4228
rect 18844 4174 18846 4226
rect 18898 4174 19236 4226
rect 18844 4172 19236 4174
rect 18844 4162 18900 4172
rect 18732 3668 18788 3678
rect 18620 3666 18788 3668
rect 18620 3614 18734 3666
rect 18786 3614 18788 3666
rect 18620 3612 18788 3614
rect 18732 3602 18788 3612
rect 17612 3350 17668 3388
rect 19180 800 19236 4172
rect 20076 4226 20132 20132
rect 20300 7362 20356 7374
rect 20300 7310 20302 7362
rect 20354 7310 20356 7362
rect 20300 6692 20356 7310
rect 20748 7362 20804 7374
rect 20748 7310 20750 7362
rect 20802 7310 20804 7362
rect 20300 6626 20356 6636
rect 20412 7252 20468 7262
rect 20412 6690 20468 7196
rect 20748 7252 20804 7310
rect 20748 7186 20804 7196
rect 20412 6638 20414 6690
rect 20466 6638 20468 6690
rect 20412 6580 20468 6638
rect 20412 6514 20468 6524
rect 20748 6804 20804 6814
rect 20524 6132 20580 6142
rect 20524 6038 20580 6076
rect 20636 5796 20692 5806
rect 20636 5702 20692 5740
rect 20748 5348 20804 6748
rect 20860 6692 20916 6702
rect 20860 6598 20916 6636
rect 21308 6020 21364 35420
rect 21868 35140 21924 35150
rect 21868 35026 21924 35084
rect 21868 34974 21870 35026
rect 21922 34974 21924 35026
rect 21868 34962 21924 34974
rect 21532 34468 21588 34478
rect 21532 33458 21588 34412
rect 21868 34468 21924 34478
rect 21868 34242 21924 34412
rect 21868 34190 21870 34242
rect 21922 34190 21924 34242
rect 21868 34178 21924 34190
rect 22204 34242 22260 34254
rect 22204 34190 22206 34242
rect 22258 34190 22260 34242
rect 21532 33406 21534 33458
rect 21586 33406 21588 33458
rect 21532 33394 21588 33406
rect 22092 33122 22148 33134
rect 22092 33070 22094 33122
rect 22146 33070 22148 33122
rect 22092 33012 22148 33070
rect 22092 32946 22148 32956
rect 22204 29988 22260 34190
rect 22204 29922 22260 29932
rect 22316 10948 22372 36316
rect 22540 35924 22596 36316
rect 22540 35858 22596 35868
rect 22764 38948 22820 38958
rect 22764 35700 22820 38892
rect 22876 36372 22932 36382
rect 22876 36278 22932 36316
rect 22764 34354 22820 35644
rect 23100 35698 23156 35710
rect 23100 35646 23102 35698
rect 23154 35646 23156 35698
rect 23100 35588 23156 35646
rect 23100 35522 23156 35532
rect 23436 35028 23492 39200
rect 24220 36708 24276 36718
rect 24220 36594 24276 36652
rect 24220 36542 24222 36594
rect 24274 36542 24276 36594
rect 24220 36530 24276 36542
rect 23884 35588 23940 35598
rect 23772 35028 23828 35038
rect 23436 35026 23828 35028
rect 23436 34974 23774 35026
rect 23826 34974 23828 35026
rect 23436 34972 23828 34974
rect 23772 34962 23828 34972
rect 22764 34302 22766 34354
rect 22818 34302 22820 34354
rect 22764 34290 22820 34302
rect 22876 34914 22932 34926
rect 22876 34862 22878 34914
rect 22930 34862 22932 34914
rect 22876 34244 22932 34862
rect 23660 34356 23716 34366
rect 23884 34356 23940 35532
rect 24220 35588 24276 35598
rect 24332 35588 24388 39200
rect 25228 36484 25284 39200
rect 25228 36428 25620 36484
rect 24220 35586 24388 35588
rect 24220 35534 24222 35586
rect 24274 35534 24388 35586
rect 24220 35532 24388 35534
rect 24780 35698 24836 35710
rect 24780 35646 24782 35698
rect 24834 35646 24836 35698
rect 24220 35522 24276 35532
rect 23660 34354 23940 34356
rect 23660 34302 23662 34354
rect 23714 34302 23940 34354
rect 23660 34300 23940 34302
rect 24220 34692 24276 34702
rect 23660 34290 23716 34300
rect 22876 34178 22932 34188
rect 23212 34244 23268 34254
rect 23212 34150 23268 34188
rect 22316 10882 22372 10892
rect 23884 34020 23940 34030
rect 21308 5954 21364 5964
rect 21532 6468 21588 6478
rect 21196 5796 21252 5806
rect 20860 5348 20916 5358
rect 20748 5346 20916 5348
rect 20748 5294 20862 5346
rect 20914 5294 20916 5346
rect 20748 5292 20916 5294
rect 20860 5282 20916 5292
rect 21196 5236 21252 5740
rect 21196 5170 21252 5180
rect 21532 5794 21588 6412
rect 21980 6020 22036 6030
rect 21980 5926 22036 5964
rect 21532 5742 21534 5794
rect 21586 5742 21588 5794
rect 21532 5124 21588 5742
rect 21756 5236 21812 5246
rect 21756 5142 21812 5180
rect 22204 5236 22260 5246
rect 22204 5142 22260 5180
rect 21532 5058 21588 5068
rect 20300 4900 20356 4910
rect 20300 4806 20356 4844
rect 21644 4900 21700 4910
rect 21644 4806 21700 4844
rect 20076 4174 20078 4226
rect 20130 4174 20132 4226
rect 20076 4162 20132 4174
rect 20524 4452 20580 4462
rect 19622 3948 19886 3958
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19622 3882 19886 3892
rect 19404 3556 19460 3566
rect 19404 3462 19460 3500
rect 20524 3444 20580 4396
rect 21084 4452 21140 4462
rect 22204 4452 22260 4462
rect 21084 4358 21140 4396
rect 21868 4450 22260 4452
rect 21868 4398 22206 4450
rect 22258 4398 22260 4450
rect 21868 4396 22260 4398
rect 20524 800 20580 3388
rect 21868 3442 21924 4396
rect 22204 4386 22260 4396
rect 23548 4228 23604 4238
rect 23884 4228 23940 33964
rect 24220 27636 24276 34636
rect 24444 34468 24500 34478
rect 24444 34354 24500 34412
rect 24780 34468 24836 35646
rect 24892 35364 24948 35374
rect 24892 34914 24948 35308
rect 24892 34862 24894 34914
rect 24946 34862 24948 34914
rect 24892 34850 24948 34862
rect 24780 34402 24836 34412
rect 24444 34302 24446 34354
rect 24498 34302 24500 34354
rect 24444 34290 24500 34302
rect 24892 34020 24948 34030
rect 24892 33926 24948 33964
rect 25228 33458 25284 36428
rect 25564 36370 25620 36428
rect 25564 36318 25566 36370
rect 25618 36318 25620 36370
rect 25564 36306 25620 36318
rect 25564 35586 25620 35598
rect 25564 35534 25566 35586
rect 25618 35534 25620 35586
rect 25564 35364 25620 35534
rect 25564 35298 25620 35308
rect 26124 35026 26180 39200
rect 26908 36594 26964 36606
rect 26908 36542 26910 36594
rect 26962 36542 26964 36594
rect 26908 36484 26964 36542
rect 26908 36418 26964 36428
rect 27020 36260 27076 39200
rect 27692 36596 27748 36606
rect 27916 36596 27972 39200
rect 27916 36540 28308 36596
rect 27692 36502 27748 36540
rect 28140 36370 28196 36382
rect 28140 36318 28142 36370
rect 28194 36318 28196 36370
rect 26796 36204 27076 36260
rect 27580 36260 27636 36270
rect 26796 35586 26852 36204
rect 26796 35534 26798 35586
rect 26850 35534 26852 35586
rect 26796 35522 26852 35534
rect 27020 35924 27076 35934
rect 26124 34974 26126 35026
rect 26178 34974 26180 35026
rect 26124 34962 26180 34974
rect 27020 34916 27076 35868
rect 27580 35698 27636 36204
rect 28140 35924 28196 36318
rect 27580 35646 27582 35698
rect 27634 35646 27636 35698
rect 27580 35634 27636 35646
rect 27804 35868 28196 35924
rect 27804 35252 27860 35868
rect 28252 35812 28308 36540
rect 27804 35186 27860 35196
rect 27916 35810 28308 35812
rect 27916 35758 28254 35810
rect 28306 35758 28308 35810
rect 27916 35756 28308 35758
rect 27020 34914 27412 34916
rect 27020 34862 27022 34914
rect 27074 34862 27412 34914
rect 27020 34860 27412 34862
rect 27020 34850 27076 34860
rect 27356 34354 27412 34860
rect 27356 34302 27358 34354
rect 27410 34302 27412 34354
rect 27356 34290 27412 34302
rect 27916 34354 27972 35756
rect 28252 35746 28308 35756
rect 28476 36258 28532 36270
rect 28476 36206 28478 36258
rect 28530 36206 28532 36258
rect 28364 35252 28420 35262
rect 28140 35140 28196 35150
rect 28140 35026 28196 35084
rect 28140 34974 28142 35026
rect 28194 34974 28196 35026
rect 28140 34962 28196 34974
rect 27916 34302 27918 34354
rect 27970 34302 27972 34354
rect 27916 34290 27972 34302
rect 28364 34354 28420 35196
rect 28364 34302 28366 34354
rect 28418 34302 28420 34354
rect 26124 34242 26180 34254
rect 26124 34190 26126 34242
rect 26178 34190 26180 34242
rect 25788 34130 25844 34142
rect 25788 34078 25790 34130
rect 25842 34078 25844 34130
rect 25788 34020 25844 34078
rect 25788 33954 25844 33964
rect 25228 33406 25230 33458
rect 25282 33406 25284 33458
rect 25228 33394 25284 33406
rect 26012 33796 26068 33806
rect 24220 27570 24276 27580
rect 26012 33124 26068 33740
rect 25004 10052 25060 10062
rect 23548 4226 23940 4228
rect 23548 4174 23550 4226
rect 23602 4174 23940 4226
rect 23548 4172 23940 4174
rect 24556 5796 24612 5806
rect 23548 4162 23604 4172
rect 23324 3668 23380 3678
rect 23324 3574 23380 3612
rect 21868 3390 21870 3442
rect 21922 3390 21924 3442
rect 21868 800 21924 3390
rect 22204 3444 22260 3454
rect 22204 3350 22260 3388
rect 23212 3444 23268 3454
rect 23212 800 23268 3388
rect 24108 3444 24164 3454
rect 24108 3350 24164 3388
rect 24556 800 24612 5740
rect 25004 3668 25060 9996
rect 25788 6468 25844 6478
rect 25676 6466 25844 6468
rect 25676 6414 25790 6466
rect 25842 6414 25844 6466
rect 25676 6412 25844 6414
rect 25116 5124 25172 5134
rect 25116 5030 25172 5068
rect 25676 5122 25732 6412
rect 25788 6402 25844 6412
rect 25788 5796 25844 5806
rect 25788 5702 25844 5740
rect 25676 5070 25678 5122
rect 25730 5070 25732 5122
rect 25676 5058 25732 5070
rect 26012 4900 26068 33068
rect 26124 26180 26180 34190
rect 28364 34020 28420 34302
rect 28364 33954 28420 33964
rect 28476 26516 28532 36206
rect 28812 35140 28868 39200
rect 29708 36596 29764 39200
rect 30044 38836 30100 38846
rect 29708 36540 29988 36596
rect 29260 36372 29316 36382
rect 29260 36278 29316 36316
rect 29820 36370 29876 36382
rect 29820 36318 29822 36370
rect 29874 36318 29876 36370
rect 29596 36148 29652 36158
rect 29596 35586 29652 36092
rect 29596 35534 29598 35586
rect 29650 35534 29652 35586
rect 29596 35522 29652 35534
rect 28812 35074 28868 35084
rect 28812 34914 28868 34926
rect 28812 34862 28814 34914
rect 28866 34862 28868 34914
rect 28476 26450 28532 26460
rect 28588 34020 28644 34030
rect 26124 26114 26180 26124
rect 28364 7586 28420 7598
rect 28364 7534 28366 7586
rect 28418 7534 28420 7586
rect 26348 7362 26404 7374
rect 26348 7310 26350 7362
rect 26402 7310 26404 7362
rect 26348 6804 26404 7310
rect 27132 7364 27188 7374
rect 27132 6914 27188 7308
rect 27132 6862 27134 6914
rect 27186 6862 27188 6914
rect 27132 6850 27188 6862
rect 26348 6738 26404 6748
rect 27804 6690 27860 6702
rect 27804 6638 27806 6690
rect 27858 6638 27860 6690
rect 26124 6580 26180 6590
rect 26796 6580 26852 6590
rect 26124 6578 26852 6580
rect 26124 6526 26126 6578
rect 26178 6526 26798 6578
rect 26850 6526 26852 6578
rect 26124 6524 26852 6526
rect 26124 6514 26180 6524
rect 26796 6514 26852 6524
rect 27804 6580 27860 6638
rect 27804 6514 27860 6524
rect 27916 6578 27972 6590
rect 27916 6526 27918 6578
rect 27970 6526 27972 6578
rect 26908 5906 26964 5918
rect 26908 5854 26910 5906
rect 26962 5854 26964 5906
rect 26908 5796 26964 5854
rect 26908 5730 26964 5740
rect 27468 5794 27524 5806
rect 27468 5742 27470 5794
rect 27522 5742 27524 5794
rect 26012 4834 26068 4844
rect 26236 4452 26292 4462
rect 25900 4450 26292 4452
rect 25900 4398 26238 4450
rect 26290 4398 26292 4450
rect 25900 4396 26292 4398
rect 25676 4228 25732 4238
rect 25900 4228 25956 4396
rect 26236 4386 26292 4396
rect 27468 4452 27524 5742
rect 27916 5796 27972 6526
rect 28028 5908 28084 5918
rect 28028 5814 28084 5852
rect 28364 5906 28420 7534
rect 28364 5854 28366 5906
rect 28418 5854 28420 5906
rect 28364 5842 28420 5854
rect 27916 5348 27972 5740
rect 27916 5282 27972 5292
rect 28252 5236 28308 5246
rect 28140 4898 28196 4910
rect 28140 4846 28142 4898
rect 28194 4846 28196 4898
rect 28140 4562 28196 4846
rect 28140 4510 28142 4562
rect 28194 4510 28196 4562
rect 28140 4498 28196 4510
rect 27468 4386 27524 4396
rect 25676 4226 25956 4228
rect 25676 4174 25678 4226
rect 25730 4174 25956 4226
rect 25676 4172 25956 4174
rect 25676 4162 25732 4172
rect 25004 3602 25060 3612
rect 25228 3444 25284 3454
rect 25228 3350 25284 3388
rect 25900 800 25956 4172
rect 27580 4228 27636 4238
rect 27580 4134 27636 4172
rect 28252 4226 28308 5180
rect 28252 4174 28254 4226
rect 28306 4174 28308 4226
rect 28252 4116 28308 4174
rect 28252 4050 28308 4060
rect 28476 3668 28532 3678
rect 28588 3668 28644 33964
rect 28812 34018 28868 34862
rect 29708 34692 29764 34702
rect 28812 33966 28814 34018
rect 28866 33966 28868 34018
rect 28812 33348 28868 33966
rect 28812 33282 28868 33292
rect 29148 34690 29764 34692
rect 29148 34638 29710 34690
rect 29762 34638 29764 34690
rect 29148 34636 29764 34638
rect 28700 7476 28756 7486
rect 28700 7474 29092 7476
rect 28700 7422 28702 7474
rect 28754 7422 29092 7474
rect 28700 7420 29092 7422
rect 28700 7410 28756 7420
rect 29036 7028 29092 7420
rect 29148 7364 29204 34636
rect 29708 34626 29764 34636
rect 29372 34356 29428 34366
rect 29372 34262 29428 34300
rect 29484 33908 29540 33918
rect 29484 33458 29540 33852
rect 29820 33908 29876 36318
rect 29932 34242 29988 36540
rect 29932 34190 29934 34242
rect 29986 34190 29988 34242
rect 29932 34178 29988 34190
rect 30044 35138 30100 38780
rect 30604 37380 30660 39200
rect 30604 37324 30996 37380
rect 30940 36596 30996 37324
rect 30604 36372 30660 36382
rect 30044 35086 30046 35138
rect 30098 35086 30100 35138
rect 29820 33842 29876 33852
rect 29484 33406 29486 33458
rect 29538 33406 29540 33458
rect 29484 10052 29540 33406
rect 30044 33460 30100 35086
rect 30044 33394 30100 33404
rect 30156 36258 30212 36270
rect 30156 36206 30158 36258
rect 30210 36206 30212 36258
rect 30156 24724 30212 36206
rect 30604 35810 30660 36316
rect 30940 36370 30996 36540
rect 30940 36318 30942 36370
rect 30994 36318 30996 36370
rect 30940 36306 30996 36318
rect 31500 35924 31556 39200
rect 32284 36596 32340 36606
rect 32284 36502 32340 36540
rect 31500 35868 31780 35924
rect 30604 35758 30606 35810
rect 30658 35758 30660 35810
rect 30604 35746 30660 35758
rect 30828 35698 30884 35710
rect 30828 35646 30830 35698
rect 30882 35646 30884 35698
rect 30828 34914 30884 35646
rect 30828 34862 30830 34914
rect 30882 34862 30884 34914
rect 30604 34802 30660 34814
rect 30604 34750 30606 34802
rect 30658 34750 30660 34802
rect 30604 34356 30660 34750
rect 30604 34290 30660 34300
rect 30828 33124 30884 34862
rect 31276 35474 31332 35486
rect 31276 35422 31278 35474
rect 31330 35422 31332 35474
rect 31052 34130 31108 34142
rect 31052 34078 31054 34130
rect 31106 34078 31108 34130
rect 31052 34018 31108 34078
rect 31052 33966 31054 34018
rect 31106 33966 31108 34018
rect 31052 33954 31108 33966
rect 30828 33030 30884 33068
rect 31276 32900 31332 35422
rect 31612 35474 31668 35486
rect 31612 35422 31614 35474
rect 31666 35422 31668 35474
rect 31500 34804 31556 34814
rect 31500 34690 31556 34748
rect 31500 34638 31502 34690
rect 31554 34638 31556 34690
rect 31276 32834 31332 32844
rect 31388 34018 31444 34030
rect 31388 33966 31390 34018
rect 31442 33966 31444 34018
rect 31388 33122 31444 33966
rect 31388 33070 31390 33122
rect 31442 33070 31444 33122
rect 31388 32340 31444 33070
rect 31388 32274 31444 32284
rect 30156 24658 30212 24668
rect 29484 9986 29540 9996
rect 30492 12740 30548 12750
rect 29148 7270 29204 7308
rect 29820 9380 29876 9390
rect 29036 6972 29764 7028
rect 29708 6914 29764 6972
rect 29708 6862 29710 6914
rect 29762 6862 29764 6914
rect 29708 6850 29764 6862
rect 28812 6580 28868 6590
rect 28812 6486 28868 6524
rect 28700 5348 28756 5358
rect 28700 5254 28756 5292
rect 29484 5124 29540 5134
rect 29484 5030 29540 5068
rect 28476 3666 28644 3668
rect 28476 3614 28478 3666
rect 28530 3614 28644 3666
rect 28476 3612 28644 3614
rect 28924 4452 28980 4462
rect 28476 3602 28532 3612
rect 26572 3444 26628 3454
rect 26572 3350 26628 3388
rect 27244 3444 27300 3454
rect 28924 3444 28980 4396
rect 29820 4228 29876 9324
rect 30044 6916 30100 6926
rect 30044 6822 30100 6860
rect 30268 6580 30324 6590
rect 30268 6486 30324 6524
rect 30268 5124 30324 5134
rect 29820 4162 29876 4172
rect 29932 5122 30324 5124
rect 29932 5070 30270 5122
rect 30322 5070 30324 5122
rect 29932 5068 30324 5070
rect 27244 800 27300 3388
rect 28588 3388 28980 3444
rect 29260 4116 29316 4126
rect 28588 800 28644 3388
rect 29260 3330 29316 4060
rect 29484 3780 29540 3790
rect 29484 3554 29540 3724
rect 29484 3502 29486 3554
rect 29538 3502 29540 3554
rect 29484 3490 29540 3502
rect 29260 3278 29262 3330
rect 29314 3278 29316 3330
rect 29260 3266 29316 3278
rect 29932 800 29988 5068
rect 30268 5058 30324 5068
rect 30268 4228 30324 4238
rect 30492 4228 30548 12684
rect 31500 7700 31556 34638
rect 31500 7634 31556 7644
rect 31612 6916 31668 35422
rect 31724 34242 31780 35868
rect 32396 35026 32452 39200
rect 32508 35810 32564 35822
rect 32508 35758 32510 35810
rect 32562 35758 32564 35810
rect 32508 35588 32564 35758
rect 33292 35812 33348 39200
rect 33516 36484 33572 36494
rect 33516 36390 33572 36428
rect 33964 36260 34020 36270
rect 33964 36166 34020 36204
rect 33740 35812 33796 35822
rect 33292 35810 33796 35812
rect 33292 35758 33742 35810
rect 33794 35758 33796 35810
rect 33292 35756 33796 35758
rect 32508 35522 32564 35532
rect 32844 35698 32900 35710
rect 32844 35646 32846 35698
rect 32898 35646 32900 35698
rect 32396 34974 32398 35026
rect 32450 34974 32452 35026
rect 32396 34962 32452 34974
rect 32844 34804 32900 35646
rect 32844 34738 32900 34748
rect 33180 34914 33236 34926
rect 33180 34862 33182 34914
rect 33234 34862 33236 34914
rect 33180 34692 33236 34862
rect 33180 34626 33236 34636
rect 33292 34804 33348 34814
rect 31724 34190 31726 34242
rect 31778 34190 31780 34242
rect 31724 34178 31780 34190
rect 32844 34356 32900 34366
rect 32844 34130 32900 34300
rect 32844 34078 32846 34130
rect 32898 34078 32900 34130
rect 32844 34066 32900 34078
rect 33292 34020 33348 34748
rect 33292 33954 33348 33964
rect 32620 33572 32676 33582
rect 31836 33460 31892 33470
rect 31836 33366 31892 33404
rect 32620 33458 32676 33516
rect 32620 33406 32622 33458
rect 32674 33406 32676 33458
rect 32284 33122 32340 33134
rect 32284 33070 32286 33122
rect 32338 33070 32340 33122
rect 31948 33012 32004 33022
rect 31836 32900 31892 32910
rect 31836 24948 31892 32844
rect 31948 31108 32004 32956
rect 32284 32900 32340 33070
rect 32620 33124 32676 33406
rect 33404 33458 33460 35756
rect 33740 35746 33796 35756
rect 34188 35026 34244 39200
rect 35084 36484 35140 39200
rect 34188 34974 34190 35026
rect 34242 34974 34244 35026
rect 34188 34962 34244 34974
rect 34300 36370 34356 36382
rect 34300 36318 34302 36370
rect 34354 36318 34356 36370
rect 33964 34692 34020 34702
rect 33516 34356 33572 34366
rect 33516 34262 33572 34300
rect 33964 34354 34020 34636
rect 33964 34302 33966 34354
rect 34018 34302 34020 34354
rect 33964 34290 34020 34302
rect 34300 34020 34356 36318
rect 35084 36370 35140 36428
rect 35084 36318 35086 36370
rect 35138 36318 35140 36370
rect 35084 36306 35140 36318
rect 35756 36708 35812 36718
rect 35756 35922 35812 36652
rect 35756 35870 35758 35922
rect 35810 35870 35812 35922
rect 35756 35812 35812 35870
rect 35756 35746 35812 35756
rect 34860 35586 34916 35598
rect 34860 35534 34862 35586
rect 34914 35534 34916 35586
rect 34524 34020 34580 34030
rect 34300 34018 34580 34020
rect 34300 33966 34526 34018
rect 34578 33966 34580 34018
rect 34300 33964 34580 33966
rect 33404 33406 33406 33458
rect 33458 33406 33460 33458
rect 33404 33394 33460 33406
rect 34524 33908 34580 33964
rect 32620 33058 32676 33068
rect 32284 32834 32340 32844
rect 31948 31042 32004 31052
rect 31836 24882 31892 24892
rect 31500 6692 31556 6702
rect 31612 6692 31668 6860
rect 31500 6690 31668 6692
rect 31500 6638 31502 6690
rect 31554 6638 31668 6690
rect 31500 6636 31668 6638
rect 32956 10836 33012 10846
rect 31500 6626 31556 6636
rect 30828 6580 30884 6590
rect 30828 6578 31444 6580
rect 30828 6526 30830 6578
rect 30882 6526 31444 6578
rect 30828 6524 31444 6526
rect 30828 6514 30884 6524
rect 30940 6130 30996 6142
rect 30940 6078 30942 6130
rect 30994 6078 30996 6130
rect 30940 5348 30996 6078
rect 30940 5282 30996 5292
rect 31388 6132 31444 6524
rect 31500 6132 31556 6142
rect 31388 6130 31556 6132
rect 31388 6078 31502 6130
rect 31554 6078 31556 6130
rect 31388 6076 31556 6078
rect 31388 5122 31444 6076
rect 31500 6066 31556 6076
rect 31836 5908 31892 5918
rect 31836 5814 31892 5852
rect 31948 5348 32004 5358
rect 31948 5254 32004 5292
rect 31388 5070 31390 5122
rect 31442 5070 31444 5122
rect 31388 5058 31444 5070
rect 32060 5124 32116 5134
rect 32508 5124 32564 5134
rect 32060 5122 32564 5124
rect 32060 5070 32062 5122
rect 32114 5070 32510 5122
rect 32562 5070 32564 5122
rect 32060 5068 32564 5070
rect 31388 4900 31444 4910
rect 31276 4452 31332 4462
rect 30268 4226 30548 4228
rect 30268 4174 30270 4226
rect 30322 4174 30548 4226
rect 30268 4172 30548 4174
rect 30716 4228 30772 4238
rect 30268 4162 30324 4172
rect 30716 4134 30772 4172
rect 30044 3780 30100 3790
rect 30044 3666 30100 3724
rect 30044 3614 30046 3666
rect 30098 3614 30100 3666
rect 30044 3556 30100 3614
rect 31164 3668 31220 3678
rect 31164 3574 31220 3612
rect 30044 3490 30100 3500
rect 31276 800 31332 4396
rect 31388 4226 31444 4844
rect 31388 4174 31390 4226
rect 31442 4174 31444 4226
rect 31388 4162 31444 4174
rect 32060 4228 32116 5068
rect 32508 5058 32564 5068
rect 32732 4452 32788 4462
rect 32732 4358 32788 4396
rect 32060 4162 32116 4172
rect 32956 3668 33012 10780
rect 34524 9268 34580 33852
rect 34860 32004 34916 35534
rect 35980 35026 36036 39200
rect 36316 37940 36372 37950
rect 36316 36594 36372 37884
rect 36316 36542 36318 36594
rect 36370 36542 36372 36594
rect 36316 36530 36372 36542
rect 36652 36372 36708 36382
rect 36540 35812 36596 35822
rect 36428 35810 36596 35812
rect 36428 35758 36542 35810
rect 36594 35758 36596 35810
rect 36428 35756 36596 35758
rect 35980 34974 35982 35026
rect 36034 34974 36036 35026
rect 35980 34962 36036 34974
rect 36204 35698 36260 35710
rect 36204 35646 36206 35698
rect 36258 35646 36260 35698
rect 34972 34916 35028 34926
rect 34972 34914 35252 34916
rect 34972 34862 34974 34914
rect 35026 34862 35252 34914
rect 34972 34860 35252 34862
rect 34972 34850 35028 34860
rect 35196 34018 35252 34860
rect 35196 33966 35198 34018
rect 35250 33966 35252 34018
rect 35196 33124 35252 33966
rect 35196 33058 35252 33068
rect 35644 34580 35700 34590
rect 35644 34354 35700 34524
rect 36204 34580 36260 35646
rect 36204 34514 36260 34524
rect 35644 34302 35646 34354
rect 35698 34302 35700 34354
rect 34860 31938 34916 31948
rect 35420 16100 35476 16110
rect 34524 9202 34580 9212
rect 34972 10948 35028 10958
rect 34972 8428 35028 10892
rect 34972 8372 35140 8428
rect 35084 8306 35140 8316
rect 32956 3602 33012 3612
rect 33404 7700 33460 7710
rect 33404 3668 33460 7644
rect 35420 5234 35476 16044
rect 35644 9380 35700 34302
rect 36092 34018 36148 34030
rect 36092 33966 36094 34018
rect 36146 33966 36148 34018
rect 36092 33460 36148 33966
rect 36092 33394 36148 33404
rect 36428 31948 36484 35756
rect 36540 35746 36596 35756
rect 36652 34804 36708 36316
rect 36876 35812 36932 39200
rect 37436 36484 37492 36494
rect 37436 36390 37492 36428
rect 37212 35812 37268 35822
rect 36876 35810 37268 35812
rect 36876 35758 37214 35810
rect 37266 35758 37268 35810
rect 36876 35756 37268 35758
rect 36652 34354 36708 34748
rect 36652 34302 36654 34354
rect 36706 34302 36708 34354
rect 36652 34290 36708 34302
rect 36764 34914 36820 34926
rect 36764 34862 36766 34914
rect 36818 34862 36820 34914
rect 36764 33460 36820 34862
rect 36764 33394 36820 33404
rect 36876 33458 36932 35756
rect 37212 35746 37268 35756
rect 36988 35028 37044 35038
rect 36988 34244 37044 34972
rect 37660 34804 37716 34814
rect 37660 34710 37716 34748
rect 37100 34468 37156 34478
rect 37100 34354 37156 34412
rect 37100 34302 37102 34354
rect 37154 34302 37156 34354
rect 37100 34290 37156 34302
rect 37772 34244 37828 39200
rect 38668 37380 38724 39200
rect 39004 37604 39060 37614
rect 38668 37324 38948 37380
rect 38892 36484 38948 37324
rect 38220 36370 38276 36382
rect 38220 36318 38222 36370
rect 38274 36318 38276 36370
rect 37884 36258 37940 36270
rect 37884 36206 37886 36258
rect 37938 36206 37940 36258
rect 37884 35028 37940 36206
rect 38220 36260 38276 36318
rect 38892 36370 38948 36428
rect 38892 36318 38894 36370
rect 38946 36318 38948 36370
rect 38892 36306 38948 36318
rect 38220 36204 38500 36260
rect 38032 36092 38296 36102
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38032 36026 38296 36036
rect 38444 35364 38500 36204
rect 38556 35588 38612 35598
rect 39004 35588 39060 37548
rect 39564 37044 39620 39200
rect 39564 36988 39956 37044
rect 38556 35586 39060 35588
rect 38556 35534 38558 35586
rect 38610 35534 39060 35586
rect 38556 35532 39060 35534
rect 39116 36036 39172 36046
rect 38556 35522 38612 35532
rect 38444 35308 38612 35364
rect 37884 34962 37940 34972
rect 38444 35028 38500 35038
rect 38444 34934 38500 34972
rect 38220 34802 38276 34814
rect 38220 34750 38222 34802
rect 38274 34750 38276 34802
rect 38220 34692 38276 34750
rect 38220 34636 38500 34692
rect 38032 34524 38296 34534
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38032 34458 38296 34468
rect 38108 34244 38164 34254
rect 37772 34242 38164 34244
rect 37772 34190 38110 34242
rect 38162 34190 38164 34242
rect 37772 34188 38164 34190
rect 36988 34178 37044 34188
rect 38108 34178 38164 34188
rect 36876 33406 36878 33458
rect 36930 33406 36932 33458
rect 36876 33394 36932 33406
rect 37436 34130 37492 34142
rect 37436 34078 37438 34130
rect 37490 34078 37492 34130
rect 37436 33124 37492 34078
rect 38444 33572 38500 34636
rect 38108 33236 38164 33246
rect 37660 33124 37716 33134
rect 38108 33124 38164 33180
rect 37436 33122 37716 33124
rect 37436 33070 37662 33122
rect 37714 33070 37716 33122
rect 37436 33068 37716 33070
rect 36428 31892 36596 31948
rect 36540 27300 36596 31892
rect 37660 27748 37716 33068
rect 37884 33122 38164 33124
rect 37884 33070 38110 33122
rect 38162 33070 38164 33122
rect 37884 33068 38164 33070
rect 37884 32676 37940 33068
rect 38108 33058 38164 33068
rect 38032 32956 38296 32966
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38032 32890 38296 32900
rect 38444 32900 38500 33516
rect 38444 32834 38500 32844
rect 37884 32610 37940 32620
rect 38444 32676 38500 32686
rect 38556 32676 38612 35308
rect 38780 34690 38836 34702
rect 38780 34638 38782 34690
rect 38834 34638 38836 34690
rect 38668 33236 38724 33246
rect 38668 33142 38724 33180
rect 38500 32620 38612 32676
rect 38032 31388 38296 31398
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38032 31322 38296 31332
rect 38032 29820 38296 29830
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38032 29754 38296 29764
rect 38032 28252 38296 28262
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38032 28186 38296 28196
rect 37660 27682 37716 27692
rect 36540 27234 36596 27244
rect 38032 26684 38296 26694
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38032 26618 38296 26628
rect 38032 25116 38296 25126
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38032 25050 38296 25060
rect 38032 23548 38296 23558
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38032 23482 38296 23492
rect 38032 21980 38296 21990
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38032 21914 38296 21924
rect 38032 20412 38296 20422
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38032 20346 38296 20356
rect 38032 18844 38296 18854
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38032 18778 38296 18788
rect 38032 17276 38296 17286
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38032 17210 38296 17220
rect 38032 15708 38296 15718
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38032 15642 38296 15652
rect 38444 15092 38500 32620
rect 38780 20188 38836 34638
rect 39116 34130 39172 35980
rect 39340 35812 39396 35822
rect 39340 35718 39396 35756
rect 39116 34078 39118 34130
rect 39170 34078 39172 34130
rect 39116 34066 39172 34078
rect 39228 35698 39284 35710
rect 39228 35646 39230 35698
rect 39282 35646 39284 35698
rect 39004 33124 39060 33134
rect 39004 33122 39172 33124
rect 39004 33070 39006 33122
rect 39058 33070 39172 33122
rect 39004 33068 39172 33070
rect 39004 33058 39060 33068
rect 39004 32900 39060 32910
rect 39004 32564 39060 32844
rect 39004 32470 39060 32508
rect 39116 27860 39172 33068
rect 39228 32900 39284 35646
rect 39228 32834 39284 32844
rect 39452 35028 39508 35038
rect 39452 32786 39508 34972
rect 39900 35026 39956 36988
rect 40460 36708 40516 39200
rect 41356 37044 41412 39200
rect 41356 36988 41860 37044
rect 40796 36708 40852 36718
rect 40460 36706 40852 36708
rect 40460 36654 40798 36706
rect 40850 36654 40852 36706
rect 40460 36652 40852 36654
rect 40796 36642 40852 36652
rect 41356 36708 41412 36718
rect 41356 36706 41748 36708
rect 41356 36654 41358 36706
rect 41410 36654 41748 36706
rect 41356 36652 41748 36654
rect 41356 36642 41412 36652
rect 40236 36596 40292 36606
rect 40236 36594 40404 36596
rect 40236 36542 40238 36594
rect 40290 36542 40404 36594
rect 40236 36540 40404 36542
rect 40236 36530 40292 36540
rect 40348 36484 40404 36540
rect 40348 36418 40404 36428
rect 41132 36260 41188 36270
rect 41132 36166 41188 36204
rect 41580 36258 41636 36270
rect 41580 36206 41582 36258
rect 41634 36206 41636 36258
rect 40012 35476 40068 35486
rect 40348 35476 40404 35486
rect 40012 35382 40068 35420
rect 40236 35474 40404 35476
rect 40236 35422 40350 35474
rect 40402 35422 40404 35474
rect 40236 35420 40404 35422
rect 39900 34974 39902 35026
rect 39954 34974 39956 35026
rect 39900 34962 39956 34974
rect 39788 34916 39844 34926
rect 39788 34356 39844 34860
rect 39900 34356 39956 34366
rect 39788 34354 39956 34356
rect 39788 34302 39902 34354
rect 39954 34302 39956 34354
rect 39788 34300 39956 34302
rect 39452 32734 39454 32786
rect 39506 32734 39508 32786
rect 39452 32722 39508 32734
rect 39564 33122 39620 33134
rect 39564 33070 39566 33122
rect 39618 33070 39620 33122
rect 39564 32340 39620 33070
rect 39564 32274 39620 32284
rect 39788 31948 39844 34300
rect 39900 34244 39956 34300
rect 39900 34178 39956 34188
rect 39900 33234 39956 33246
rect 39900 33182 39902 33234
rect 39954 33182 39956 33234
rect 39900 32788 39956 33182
rect 40124 32788 40180 32798
rect 39900 32786 40180 32788
rect 39900 32734 40126 32786
rect 40178 32734 40180 32786
rect 39900 32732 40180 32734
rect 39788 31892 39956 31948
rect 39116 27794 39172 27804
rect 38780 20132 39284 20188
rect 38444 15026 38500 15036
rect 38032 14140 38296 14150
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38032 14074 38296 14084
rect 38032 12572 38296 12582
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38032 12506 38296 12516
rect 38032 11004 38296 11014
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38032 10938 38296 10948
rect 38032 9436 38296 9446
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38032 9370 38296 9380
rect 35644 9314 35700 9324
rect 38032 7868 38296 7878
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38032 7802 38296 7812
rect 37884 7364 37940 7374
rect 37436 6580 37492 6590
rect 36764 6020 36820 6030
rect 36764 5906 36820 5964
rect 36764 5854 36766 5906
rect 36818 5854 36820 5906
rect 36764 5842 36820 5854
rect 37436 6020 37492 6524
rect 35420 5182 35422 5234
rect 35474 5182 35476 5234
rect 35420 5170 35476 5182
rect 35644 5794 35700 5806
rect 35644 5742 35646 5794
rect 35698 5742 35700 5794
rect 35532 5124 35588 5134
rect 34300 5010 34356 5022
rect 34300 4958 34302 5010
rect 34354 4958 34356 5010
rect 33740 4900 33796 4910
rect 34300 4900 34356 4958
rect 33740 4898 34356 4900
rect 33740 4846 33742 4898
rect 33794 4846 34356 4898
rect 33740 4844 34356 4846
rect 33740 4834 33796 4844
rect 33516 4452 33572 4462
rect 33516 4358 33572 4396
rect 33404 3602 33460 3612
rect 32284 3444 32340 3454
rect 33068 3444 33124 3454
rect 32284 3442 33124 3444
rect 32284 3390 32286 3442
rect 32338 3390 33070 3442
rect 33122 3390 33124 3442
rect 32284 3388 33124 3390
rect 32284 3378 32340 3388
rect 32620 800 32676 3388
rect 33068 3378 33124 3388
rect 33964 800 34020 4844
rect 35532 4338 35588 5068
rect 35532 4286 35534 4338
rect 35586 4286 35588 4338
rect 34860 3668 34916 3678
rect 34860 3574 34916 3612
rect 35532 3668 35588 4286
rect 35532 3602 35588 3612
rect 35644 980 35700 5742
rect 36764 5684 36820 5694
rect 36764 5010 36820 5628
rect 37436 5346 37492 5964
rect 37884 5906 37940 7308
rect 39228 7364 39284 20132
rect 39900 12740 39956 31892
rect 40124 31892 40180 32732
rect 40124 31826 40180 31836
rect 39900 12674 39956 12684
rect 39228 7270 39284 7308
rect 39788 7362 39844 7374
rect 39788 7310 39790 7362
rect 39842 7310 39844 7362
rect 39116 6804 39172 6814
rect 39116 6710 39172 6748
rect 38332 6580 38388 6590
rect 38332 6486 38388 6524
rect 38892 6578 38948 6590
rect 38892 6526 38894 6578
rect 38946 6526 38948 6578
rect 38892 6468 38948 6526
rect 38032 6300 38296 6310
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38032 6234 38296 6244
rect 37884 5854 37886 5906
rect 37938 5854 37940 5906
rect 37884 5842 37940 5854
rect 38444 6018 38500 6030
rect 38444 5966 38446 6018
rect 38498 5966 38500 6018
rect 37548 5684 37604 5694
rect 37548 5590 37604 5628
rect 38220 5684 38276 5694
rect 37436 5294 37438 5346
rect 37490 5294 37492 5346
rect 37436 5282 37492 5294
rect 36764 4958 36766 5010
rect 36818 4958 36820 5010
rect 36764 4946 36820 4958
rect 38220 5010 38276 5628
rect 38220 4958 38222 5010
rect 38274 4958 38276 5010
rect 38220 4946 38276 4958
rect 36428 4900 36484 4910
rect 36092 4898 36484 4900
rect 36092 4846 36430 4898
rect 36482 4846 36484 4898
rect 36092 4844 36484 4846
rect 36092 4338 36148 4844
rect 36428 4834 36484 4844
rect 38032 4732 38296 4742
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38032 4666 38296 4676
rect 38444 4564 38500 5966
rect 38668 5908 38724 5918
rect 38892 5908 38948 6412
rect 38668 5906 38948 5908
rect 38668 5854 38670 5906
rect 38722 5854 38948 5906
rect 38668 5852 38948 5854
rect 39452 6466 39508 6478
rect 39452 6414 39454 6466
rect 39506 6414 39508 6466
rect 39452 5906 39508 6414
rect 39788 6468 39844 7310
rect 40124 6804 40180 6814
rect 40236 6804 40292 35420
rect 40348 35410 40404 35420
rect 41580 35364 41636 36206
rect 41580 35298 41636 35308
rect 41692 35810 41748 36652
rect 41692 35758 41694 35810
rect 41746 35758 41748 35810
rect 41020 34914 41076 34926
rect 41020 34862 41022 34914
rect 41074 34862 41076 34914
rect 40460 34244 40516 34254
rect 40460 34150 40516 34188
rect 40796 34242 40852 34254
rect 40796 34190 40798 34242
rect 40850 34190 40852 34242
rect 40796 34132 40852 34190
rect 40796 34066 40852 34076
rect 41020 33684 41076 34862
rect 41580 34018 41636 34030
rect 41580 33966 41582 34018
rect 41634 33966 41636 34018
rect 41580 33796 41636 33966
rect 41580 33730 41636 33740
rect 41020 33618 41076 33628
rect 40460 33234 40516 33246
rect 40460 33182 40462 33234
rect 40514 33182 40516 33234
rect 40460 32788 40516 33182
rect 40796 33124 40852 33134
rect 40796 33122 40964 33124
rect 40796 33070 40798 33122
rect 40850 33070 40964 33122
rect 40796 33068 40964 33070
rect 40796 33058 40852 33068
rect 40460 32722 40516 32732
rect 40796 32564 40852 32574
rect 40796 32470 40852 32508
rect 40908 29316 40964 33068
rect 40908 29250 40964 29260
rect 41244 33122 41300 33134
rect 41244 33070 41246 33122
rect 41298 33070 41300 33122
rect 41244 32788 41300 33070
rect 40180 6748 40292 6804
rect 40572 10948 40628 10958
rect 40572 8372 40628 10892
rect 41244 10836 41300 32732
rect 41580 32788 41636 32798
rect 41692 32788 41748 35758
rect 41804 35026 41860 36988
rect 41804 34974 41806 35026
rect 41858 34974 41860 35026
rect 41804 34962 41860 34974
rect 41916 36370 41972 36382
rect 41916 36318 41918 36370
rect 41970 36318 41972 36370
rect 41804 33684 41860 33694
rect 41804 33458 41860 33628
rect 41916 33572 41972 36318
rect 42252 36372 42308 39200
rect 43036 38052 43092 38062
rect 42588 36372 42644 36382
rect 42252 36370 42644 36372
rect 42252 36318 42590 36370
rect 42642 36318 42644 36370
rect 42252 36316 42644 36318
rect 41916 33506 41972 33516
rect 42028 35476 42084 35486
rect 41804 33406 41806 33458
rect 41858 33406 41860 33458
rect 41804 33394 41860 33406
rect 41580 32786 41748 32788
rect 41580 32734 41582 32786
rect 41634 32734 41748 32786
rect 41580 32732 41748 32734
rect 42028 32786 42084 35420
rect 42476 34242 42532 34254
rect 42476 34190 42478 34242
rect 42530 34190 42532 34242
rect 42140 34130 42196 34142
rect 42140 34078 42142 34130
rect 42194 34078 42196 34130
rect 42140 33796 42196 34078
rect 42140 33730 42196 33740
rect 42028 32734 42030 32786
rect 42082 32734 42084 32786
rect 41580 32722 41636 32732
rect 42028 24836 42084 32734
rect 42028 24770 42084 24780
rect 42140 33572 42196 33582
rect 42140 33458 42196 33516
rect 42140 33406 42142 33458
rect 42194 33406 42196 33458
rect 42140 33012 42196 33406
rect 42364 33572 42420 33582
rect 42364 33124 42420 33516
rect 42364 33058 42420 33068
rect 42140 13412 42196 32956
rect 42476 27188 42532 34190
rect 42588 33460 42644 36316
rect 43036 35586 43092 37996
rect 43148 37044 43204 39200
rect 43932 38724 43988 38734
rect 43148 36988 43540 37044
rect 43036 35534 43038 35586
rect 43090 35534 43092 35586
rect 43036 35522 43092 35534
rect 42812 35140 42868 35150
rect 42812 34914 42868 35084
rect 42812 34862 42814 34914
rect 42866 34862 42868 34914
rect 42812 34850 42868 34862
rect 43148 35140 43204 35150
rect 43148 34354 43204 35084
rect 43484 35026 43540 36988
rect 43932 36594 43988 38668
rect 43932 36542 43934 36594
rect 43986 36542 43988 36594
rect 43932 36530 43988 36542
rect 44044 36260 44100 39200
rect 43820 36204 44100 36260
rect 43596 35924 43652 35934
rect 43820 35924 43876 36204
rect 43596 35922 43876 35924
rect 43596 35870 43598 35922
rect 43650 35870 43876 35922
rect 43596 35868 43876 35870
rect 43596 35858 43652 35868
rect 44044 35812 44100 36204
rect 44604 37268 44660 37278
rect 44156 35812 44212 35822
rect 44044 35810 44212 35812
rect 44044 35758 44158 35810
rect 44210 35758 44212 35810
rect 44044 35756 44212 35758
rect 44156 35746 44212 35756
rect 43484 34974 43486 35026
rect 43538 34974 43540 35026
rect 43484 34962 43540 34974
rect 44604 34916 44660 37212
rect 44940 36260 44996 39200
rect 45276 37044 45332 37054
rect 45276 36372 45332 36988
rect 45836 36708 45892 39200
rect 45836 36652 46228 36708
rect 45948 36484 46004 36494
rect 44940 36204 45220 36260
rect 43148 34302 43150 34354
rect 43202 34302 43204 34354
rect 43148 34290 43204 34302
rect 44268 34914 44660 34916
rect 44268 34862 44606 34914
rect 44658 34862 44660 34914
rect 44268 34860 44660 34862
rect 44268 34354 44324 34860
rect 44604 34850 44660 34860
rect 44716 36148 44772 36158
rect 44268 34302 44270 34354
rect 44322 34302 44324 34354
rect 44268 34290 44324 34302
rect 44716 34692 44772 36092
rect 44716 34354 44772 34636
rect 44716 34302 44718 34354
rect 44770 34302 44772 34354
rect 44716 34290 44772 34302
rect 45164 34244 45220 36204
rect 45276 34468 45332 36316
rect 45836 36482 46004 36484
rect 45836 36430 45950 36482
rect 46002 36430 46004 36482
rect 45836 36428 46004 36430
rect 45724 36258 45780 36270
rect 45724 36206 45726 36258
rect 45778 36206 45780 36258
rect 45724 36036 45780 36206
rect 45724 35970 45780 35980
rect 45836 36260 45892 36428
rect 45948 36418 46004 36428
rect 45500 35588 45556 35598
rect 45500 35586 45780 35588
rect 45500 35534 45502 35586
rect 45554 35534 45780 35586
rect 45500 35532 45780 35534
rect 45500 35522 45556 35532
rect 45612 34916 45668 34926
rect 45612 34822 45668 34860
rect 45276 34412 45444 34468
rect 45276 34244 45332 34254
rect 45164 34242 45332 34244
rect 45164 34190 45278 34242
rect 45330 34190 45332 34242
rect 45164 34188 45332 34190
rect 45276 34178 45332 34188
rect 44604 34132 44660 34142
rect 43596 33796 43652 33806
rect 43148 33740 43596 33796
rect 43148 33684 43204 33740
rect 43596 33730 43652 33740
rect 43148 33618 43204 33628
rect 42700 33460 42756 33470
rect 42588 33458 42756 33460
rect 42588 33406 42702 33458
rect 42754 33406 42756 33458
rect 42588 33404 42756 33406
rect 42700 33394 42756 33404
rect 44604 31220 44660 34076
rect 45388 34020 45444 34412
rect 45276 33964 45444 34020
rect 44604 31154 44660 31164
rect 45052 31892 45108 31902
rect 42476 27122 42532 27132
rect 42812 27748 42868 27758
rect 42140 13346 42196 13356
rect 41244 10770 41300 10780
rect 40124 6672 40180 6748
rect 39788 6402 39844 6412
rect 40460 6468 40516 6478
rect 40460 6374 40516 6412
rect 39676 6020 39732 6030
rect 39676 5926 39732 5964
rect 40460 6020 40516 6030
rect 39452 5854 39454 5906
rect 39506 5854 39508 5906
rect 38668 5842 38724 5852
rect 39452 5842 39508 5854
rect 40236 5796 40292 5806
rect 40236 5702 40292 5740
rect 40348 5684 40404 5694
rect 40348 5590 40404 5628
rect 38444 4498 38500 4508
rect 38556 5124 38612 5134
rect 38556 4562 38612 5068
rect 40460 5122 40516 5964
rect 40460 5070 40462 5122
rect 40514 5070 40516 5122
rect 40460 5058 40516 5070
rect 38556 4510 38558 4562
rect 38610 4510 38612 4562
rect 38556 4498 38612 4510
rect 39116 4564 39172 4574
rect 39116 4470 39172 4508
rect 39564 4564 39620 4574
rect 36092 4286 36094 4338
rect 36146 4286 36148 4338
rect 36092 4274 36148 4286
rect 39564 4338 39620 4508
rect 39564 4286 39566 4338
rect 39618 4286 39620 4338
rect 39564 4274 39620 4286
rect 40236 4340 40292 4350
rect 39340 4228 39396 4238
rect 36204 3444 36260 3454
rect 36204 3350 36260 3388
rect 36876 3444 36932 3454
rect 36988 3444 37044 3454
rect 36932 3442 37044 3444
rect 36932 3390 36990 3442
rect 37042 3390 37044 3442
rect 36932 3388 37044 3390
rect 36876 2212 36932 3388
rect 36988 3378 37044 3388
rect 37772 3444 37828 3454
rect 37772 2324 37828 3388
rect 38332 3444 38388 3454
rect 38332 3350 38388 3388
rect 38032 3164 38296 3174
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38032 3098 38296 3108
rect 37772 2268 38052 2324
rect 35308 924 35700 980
rect 36652 2156 36932 2212
rect 35308 800 35364 924
rect 36652 800 36708 2156
rect 37996 800 38052 2268
rect 39340 800 39396 4172
rect 39676 3780 39732 3790
rect 39676 3666 39732 3724
rect 39676 3614 39678 3666
rect 39730 3614 39732 3666
rect 39676 3602 39732 3614
rect 40236 3668 40292 4284
rect 40348 4228 40404 4238
rect 40348 4134 40404 4172
rect 40572 3780 40628 8316
rect 41020 5908 41076 5918
rect 40908 5796 40964 5806
rect 40908 5236 40964 5740
rect 40908 5170 40964 5180
rect 41020 5122 41076 5852
rect 41468 5908 41524 5918
rect 41468 5814 41524 5852
rect 41692 5236 41748 5246
rect 41692 5142 41748 5180
rect 41020 5070 41022 5122
rect 41074 5070 41076 5122
rect 41020 5058 41076 5070
rect 41580 5124 41636 5134
rect 41580 5030 41636 5068
rect 42252 5124 42308 5134
rect 42252 5030 42308 5068
rect 40572 3714 40628 3724
rect 41692 4450 41748 4462
rect 41692 4398 41694 4450
rect 41746 4398 41748 4450
rect 40236 3574 40292 3612
rect 40684 3444 40740 3454
rect 40684 800 40740 3388
rect 41244 3444 41300 3454
rect 41244 3350 41300 3388
rect 41692 3444 41748 4398
rect 42812 4226 42868 27692
rect 45052 23380 45108 31836
rect 43932 15092 43988 15102
rect 43596 5012 43652 5022
rect 42812 4174 42814 4226
rect 42866 4174 42868 4226
rect 42812 4162 42868 4174
rect 43372 5010 43652 5012
rect 43372 4958 43598 5010
rect 43650 4958 43652 5010
rect 43372 4956 43652 4958
rect 41692 3378 41748 3388
rect 41804 3444 41860 3454
rect 42364 3444 42420 3454
rect 41804 3442 42420 3444
rect 41804 3390 41806 3442
rect 41858 3390 42366 3442
rect 42418 3390 42420 3442
rect 41804 3388 42420 3390
rect 41804 3378 41860 3388
rect 42028 800 42084 3388
rect 42364 3378 42420 3388
rect 43372 800 43428 4956
rect 43596 4946 43652 4956
rect 43708 3668 43764 3678
rect 43932 3668 43988 15036
rect 44604 5460 44660 5470
rect 44604 5122 44660 5404
rect 44604 5070 44606 5122
rect 44658 5070 44660 5122
rect 44604 5058 44660 5070
rect 43708 3666 43988 3668
rect 43708 3614 43710 3666
rect 43762 3614 43988 3666
rect 43708 3612 43988 3614
rect 44716 5012 44772 5022
rect 43708 3602 43764 3612
rect 44716 800 44772 4956
rect 45052 4228 45108 23324
rect 45276 16100 45332 33964
rect 45500 33570 45556 33582
rect 45500 33518 45502 33570
rect 45554 33518 45556 33570
rect 45500 33458 45556 33518
rect 45500 33406 45502 33458
rect 45554 33406 45556 33458
rect 45500 33394 45556 33406
rect 45388 33124 45444 33134
rect 45388 31780 45444 33068
rect 45388 31714 45444 31724
rect 45724 20132 45780 35532
rect 45836 23044 45892 36204
rect 46172 35810 46228 36652
rect 46732 36596 46788 39200
rect 47404 36596 47460 36606
rect 46732 36540 47012 36596
rect 46844 36372 46900 36382
rect 46844 36278 46900 36316
rect 46172 35758 46174 35810
rect 46226 35758 46228 35810
rect 46060 34690 46116 34702
rect 46060 34638 46062 34690
rect 46114 34638 46116 34690
rect 46060 34356 46116 34638
rect 46060 34290 46116 34300
rect 46172 33570 46228 35758
rect 46172 33518 46174 33570
rect 46226 33518 46228 33570
rect 46172 33506 46228 33518
rect 46284 36148 46340 36158
rect 46284 34130 46340 36092
rect 46396 35364 46452 35374
rect 46396 34916 46452 35308
rect 46396 34914 46564 34916
rect 46396 34862 46398 34914
rect 46450 34862 46564 34914
rect 46396 34860 46564 34862
rect 46396 34850 46452 34860
rect 46284 34078 46286 34130
rect 46338 34078 46340 34130
rect 45948 33348 46004 33358
rect 46284 33348 46340 34078
rect 45948 33346 46340 33348
rect 45948 33294 45950 33346
rect 46002 33294 46340 33346
rect 45948 33292 46340 33294
rect 46396 34468 46452 34478
rect 45948 33282 46004 33292
rect 46396 33234 46452 34412
rect 46396 33182 46398 33234
rect 46450 33182 46452 33234
rect 46396 33170 46452 33182
rect 45836 22978 45892 22988
rect 46508 32786 46564 34860
rect 46956 34244 47012 36540
rect 47292 35588 47348 35598
rect 47180 35586 47348 35588
rect 47180 35534 47294 35586
rect 47346 35534 47348 35586
rect 47180 35532 47348 35534
rect 47068 34802 47124 34814
rect 47068 34750 47070 34802
rect 47122 34750 47124 34802
rect 47068 34692 47124 34750
rect 47068 34626 47124 34636
rect 47068 34244 47124 34254
rect 46956 34242 47124 34244
rect 46956 34190 47070 34242
rect 47122 34190 47124 34242
rect 46956 34188 47124 34190
rect 47068 34178 47124 34188
rect 46508 32734 46510 32786
rect 46562 32734 46564 32786
rect 45724 20066 45780 20076
rect 45276 16034 45332 16044
rect 46508 14420 46564 32734
rect 46732 33234 46788 33246
rect 46732 33182 46734 33234
rect 46786 33182 46788 33234
rect 46732 32788 46788 33182
rect 46956 32788 47012 32798
rect 46732 32786 47012 32788
rect 46732 32734 46958 32786
rect 47010 32734 47012 32786
rect 46732 32732 47012 32734
rect 46956 32116 47012 32732
rect 46956 32050 47012 32060
rect 47180 28084 47236 35532
rect 47292 35522 47348 35532
rect 47180 28018 47236 28028
rect 47292 34916 47348 34926
rect 47292 26404 47348 34860
rect 47404 34692 47460 36540
rect 47628 36372 47684 39200
rect 48076 36596 48132 36606
rect 48076 36502 48132 36540
rect 47516 35028 47572 35038
rect 47516 34802 47572 34972
rect 47516 34750 47518 34802
rect 47570 34750 47572 34802
rect 47516 34738 47572 34750
rect 47404 33460 47460 34636
rect 47516 33460 47572 33470
rect 47404 33458 47572 33460
rect 47404 33406 47518 33458
rect 47570 33406 47572 33458
rect 47404 33404 47572 33406
rect 47516 33394 47572 33404
rect 47628 32786 47684 36316
rect 48412 35924 48468 35934
rect 48412 35830 48468 35868
rect 48300 35028 48356 35038
rect 47852 34916 47908 34926
rect 47852 34822 47908 34860
rect 48188 34692 48244 34702
rect 47628 32734 47630 32786
rect 47682 32734 47684 32786
rect 47628 32722 47684 32734
rect 47852 34690 48244 34692
rect 47852 34638 48190 34690
rect 48242 34638 48244 34690
rect 47852 34636 48244 34638
rect 47292 26338 47348 26348
rect 46508 14354 46564 14364
rect 46732 13412 46788 13422
rect 46620 6020 46676 6030
rect 45836 6018 46676 6020
rect 45836 5966 46622 6018
rect 46674 5966 46676 6018
rect 45836 5964 46676 5966
rect 45276 5794 45332 5806
rect 45276 5742 45278 5794
rect 45330 5742 45332 5794
rect 45276 5012 45332 5742
rect 45276 4946 45332 4956
rect 45612 5012 45668 5022
rect 45612 4918 45668 4956
rect 45052 4162 45108 4172
rect 45276 4340 45332 4350
rect 45276 3444 45332 4284
rect 45836 4338 45892 5964
rect 46620 5954 46676 5964
rect 45836 4286 45838 4338
rect 45890 4286 45892 4338
rect 45836 4274 45892 4286
rect 46732 3668 46788 13356
rect 47068 9268 47124 9278
rect 46956 6020 47012 6030
rect 46956 5926 47012 5964
rect 46956 5236 47012 5246
rect 47068 5236 47124 9212
rect 47852 7476 47908 34636
rect 48188 34626 48244 34636
rect 48188 34356 48244 34366
rect 48188 34130 48244 34300
rect 48188 34078 48190 34130
rect 48242 34078 48244 34130
rect 48188 34066 48244 34078
rect 48300 33908 48356 34972
rect 48524 34244 48580 39200
rect 49420 36932 49476 39200
rect 49420 36876 49812 36932
rect 49532 36708 49588 36718
rect 49196 36484 49252 36494
rect 49196 36390 49252 36428
rect 48748 35700 48804 35710
rect 48804 35644 48916 35700
rect 48748 35606 48804 35644
rect 48748 34356 48804 34366
rect 48748 34262 48804 34300
rect 48524 34178 48580 34188
rect 48188 33852 48356 33908
rect 48860 33908 48916 35644
rect 49532 35252 49588 36652
rect 49644 36370 49700 36382
rect 49644 36318 49646 36370
rect 49698 36318 49700 36370
rect 49644 36260 49700 36318
rect 49644 36194 49700 36204
rect 49756 35812 49812 36876
rect 49980 36260 50036 36270
rect 49980 36166 50036 36204
rect 49756 35810 50036 35812
rect 49756 35758 49758 35810
rect 49810 35758 50036 35810
rect 49756 35756 50036 35758
rect 49756 35746 49812 35756
rect 49532 35196 49812 35252
rect 49756 35138 49812 35196
rect 49756 35086 49758 35138
rect 49810 35086 49812 35138
rect 49532 34916 49588 34926
rect 48972 34802 49028 34814
rect 48972 34750 48974 34802
rect 49026 34750 49028 34802
rect 48972 34692 49028 34750
rect 49532 34802 49588 34860
rect 49532 34750 49534 34802
rect 49586 34750 49588 34802
rect 49532 34738 49588 34750
rect 48972 34626 49028 34636
rect 49644 34244 49700 34254
rect 49644 34150 49700 34188
rect 49756 33908 49812 35086
rect 48860 33852 49028 33908
rect 47964 33572 48020 33582
rect 47964 33234 48020 33516
rect 47964 33182 47966 33234
rect 48018 33182 48020 33234
rect 47964 33170 48020 33182
rect 48188 32786 48244 33852
rect 48860 33348 48916 33358
rect 48188 32734 48190 32786
rect 48242 32734 48244 32786
rect 48188 32722 48244 32734
rect 48300 33234 48356 33246
rect 48300 33182 48302 33234
rect 48354 33182 48356 33234
rect 48300 32564 48356 33182
rect 48860 33234 48916 33292
rect 48860 33182 48862 33234
rect 48914 33182 48916 33234
rect 48860 33170 48916 33182
rect 48524 32564 48580 32574
rect 48300 32508 48524 32564
rect 48524 32470 48580 32508
rect 48972 31554 49028 33852
rect 49756 33842 49812 33852
rect 48972 31502 48974 31554
rect 49026 31502 49028 31554
rect 48972 16884 49028 31502
rect 49196 33236 49252 33246
rect 49196 23492 49252 33180
rect 49420 33236 49476 33246
rect 49420 32786 49476 33180
rect 49868 33124 49924 33134
rect 49868 33030 49924 33068
rect 49420 32734 49422 32786
rect 49474 32734 49476 32786
rect 49420 32722 49476 32734
rect 49868 32788 49924 32798
rect 49980 32788 50036 35756
rect 50204 35476 50260 35486
rect 49868 32786 50036 32788
rect 49868 32734 49870 32786
rect 49922 32734 50036 32786
rect 49868 32732 50036 32734
rect 50092 34690 50148 34702
rect 50092 34638 50094 34690
rect 50146 34638 50148 34690
rect 49868 32722 49924 32732
rect 49196 23426 49252 23436
rect 48972 16818 49028 16828
rect 47852 6914 47908 7420
rect 48748 7476 48804 7486
rect 48748 7382 48804 7420
rect 50092 7476 50148 34638
rect 50204 33346 50260 35420
rect 50316 35028 50372 39200
rect 51212 37380 51268 39200
rect 50988 37324 51268 37380
rect 50988 36484 51044 37324
rect 52108 36708 52164 39200
rect 52108 36652 52388 36708
rect 51996 36596 52052 36606
rect 51996 36594 52164 36596
rect 51996 36542 51998 36594
rect 52050 36542 52164 36594
rect 51996 36540 52164 36542
rect 51996 36530 52052 36540
rect 50988 36370 51044 36428
rect 50988 36318 50990 36370
rect 51042 36318 51044 36370
rect 50988 36306 51044 36318
rect 51548 36260 51604 36270
rect 51100 36036 51156 36046
rect 50316 34962 50372 34972
rect 50428 35588 50484 35598
rect 50204 33294 50206 33346
rect 50258 33294 50260 33346
rect 50204 33282 50260 33294
rect 50428 34916 50484 35532
rect 51100 35586 51156 35980
rect 51100 35534 51102 35586
rect 51154 35534 51156 35586
rect 51100 35522 51156 35534
rect 50876 35028 50932 35038
rect 50876 34934 50932 34972
rect 50428 32788 50484 34860
rect 50764 34244 50820 34254
rect 50764 34130 50820 34188
rect 50764 34078 50766 34130
rect 50818 34078 50820 34130
rect 50764 34066 50820 34078
rect 51436 34242 51492 34254
rect 51436 34190 51438 34242
rect 51490 34190 51492 34242
rect 50764 33908 50820 33918
rect 50764 33458 50820 33852
rect 51436 33796 51492 34190
rect 51436 33730 51492 33740
rect 51324 33572 51380 33582
rect 50764 33406 50766 33458
rect 50818 33406 50820 33458
rect 50764 33394 50820 33406
rect 51212 33460 51268 33470
rect 51212 33234 51268 33404
rect 51212 33182 51214 33234
rect 51266 33182 51268 33234
rect 51212 33170 51268 33182
rect 50540 32788 50596 32798
rect 50428 32786 50596 32788
rect 50428 32734 50542 32786
rect 50594 32734 50596 32786
rect 50428 32732 50596 32734
rect 50540 32722 50596 32732
rect 51324 32450 51380 33516
rect 51548 33460 51604 36204
rect 51660 35476 51716 35486
rect 51996 35476 52052 35486
rect 51660 35382 51716 35420
rect 51884 35474 52052 35476
rect 51884 35422 51998 35474
rect 52050 35422 52052 35474
rect 51884 35420 52052 35422
rect 51772 34130 51828 34142
rect 51772 34078 51774 34130
rect 51826 34078 51828 34130
rect 51772 33796 51828 34078
rect 51772 33730 51828 33740
rect 51548 33404 51716 33460
rect 51548 33234 51604 33246
rect 51548 33182 51550 33234
rect 51602 33182 51604 33234
rect 51548 32900 51604 33182
rect 51548 32834 51604 32844
rect 51324 32398 51326 32450
rect 51378 32398 51380 32450
rect 51324 17668 51380 32398
rect 51660 27972 51716 33404
rect 51884 31780 51940 35420
rect 51996 35410 52052 35420
rect 51996 34914 52052 34926
rect 51996 34862 51998 34914
rect 52050 34862 52052 34914
rect 51996 34804 52052 34862
rect 51996 34738 52052 34748
rect 51996 33122 52052 33134
rect 51996 33070 51998 33122
rect 52050 33070 52052 33122
rect 51996 32900 52052 33070
rect 51996 32834 52052 32844
rect 51884 31714 51940 31724
rect 51660 27906 51716 27916
rect 52108 24612 52164 36540
rect 52220 35812 52276 35822
rect 52220 35718 52276 35756
rect 52332 34244 52388 36652
rect 52892 36372 52948 36382
rect 52780 35924 52836 35934
rect 52668 35812 52724 35822
rect 52668 35586 52724 35756
rect 52668 35534 52670 35586
rect 52722 35534 52724 35586
rect 52668 35476 52724 35534
rect 52556 35420 52724 35476
rect 52556 34802 52612 35420
rect 52668 35140 52724 35150
rect 52780 35140 52836 35868
rect 52668 35138 52836 35140
rect 52668 35086 52670 35138
rect 52722 35086 52836 35138
rect 52668 35084 52836 35086
rect 52668 35074 52724 35084
rect 52556 34750 52558 34802
rect 52610 34750 52612 34802
rect 52444 34244 52500 34254
rect 52332 34242 52500 34244
rect 52332 34190 52446 34242
rect 52498 34190 52500 34242
rect 52332 34188 52500 34190
rect 52444 34178 52500 34188
rect 52108 24546 52164 24556
rect 52444 33796 52500 33806
rect 52444 33458 52500 33740
rect 52556 33572 52612 34750
rect 52892 34580 52948 36316
rect 53004 35812 53060 39200
rect 53116 36484 53172 36494
rect 53116 36390 53172 36428
rect 53788 36482 53844 36494
rect 53788 36430 53790 36482
rect 53842 36430 53844 36482
rect 53564 36258 53620 36270
rect 53564 36206 53566 36258
rect 53618 36206 53620 36258
rect 53340 35812 53396 35822
rect 53004 35810 53396 35812
rect 53004 35758 53342 35810
rect 53394 35758 53396 35810
rect 53004 35756 53396 35758
rect 52892 34514 52948 34524
rect 52556 33506 52612 33516
rect 52444 33406 52446 33458
rect 52498 33406 52500 33458
rect 52444 22932 52500 33406
rect 53340 33460 53396 35756
rect 53564 35140 53620 36206
rect 53564 35074 53620 35084
rect 53676 34692 53732 34702
rect 53788 34692 53844 36430
rect 53900 35028 53956 39200
rect 54796 36484 54852 39200
rect 55692 37156 55748 39200
rect 54796 36370 54852 36428
rect 54796 36318 54798 36370
rect 54850 36318 54852 36370
rect 54796 36306 54852 36318
rect 55580 37100 55748 37156
rect 56252 38164 56308 38174
rect 55580 35810 55636 37100
rect 55580 35758 55582 35810
rect 55634 35758 55636 35810
rect 55580 35746 55636 35758
rect 55692 36594 55748 36606
rect 55692 36542 55694 36594
rect 55746 36542 55748 36594
rect 54572 35700 54628 35710
rect 54460 35588 54516 35598
rect 54348 35586 54516 35588
rect 54348 35534 54462 35586
rect 54514 35534 54516 35586
rect 54348 35532 54516 35534
rect 54236 35028 54292 35038
rect 53900 35026 54292 35028
rect 53900 34974 54238 35026
rect 54290 34974 54292 35026
rect 53900 34972 54292 34974
rect 54236 34962 54292 34972
rect 53676 34690 53844 34692
rect 53676 34638 53678 34690
rect 53730 34638 53844 34690
rect 53676 34636 53844 34638
rect 53564 34130 53620 34142
rect 53564 34078 53566 34130
rect 53618 34078 53620 34130
rect 53452 33460 53508 33470
rect 53340 33458 53508 33460
rect 53340 33406 53454 33458
rect 53506 33406 53508 33458
rect 53340 33404 53508 33406
rect 53452 33394 53508 33404
rect 53564 33460 53620 34078
rect 53564 33394 53620 33404
rect 52556 32450 52612 32462
rect 52556 32398 52558 32450
rect 52610 32398 52612 32450
rect 52556 31780 52612 32398
rect 52556 31714 52612 31724
rect 52444 22866 52500 22876
rect 52892 23492 52948 23502
rect 52892 20188 52948 23436
rect 52892 20132 53060 20188
rect 51324 17602 51380 17612
rect 51436 16884 51492 16894
rect 50316 8484 50372 8494
rect 50316 7588 50372 8428
rect 50316 7494 50372 7532
rect 48412 7364 48468 7374
rect 47852 6862 47854 6914
rect 47906 6862 47908 6914
rect 47852 6850 47908 6862
rect 48300 7362 48468 7364
rect 48300 7310 48414 7362
rect 48466 7310 48468 7362
rect 48300 7308 48468 7310
rect 48300 6692 48356 7308
rect 48412 7298 48468 7308
rect 49756 7362 49812 7374
rect 49756 7310 49758 7362
rect 49810 7310 49812 7362
rect 49756 7252 49812 7310
rect 49756 7186 49812 7196
rect 50092 6916 50148 7420
rect 50540 7474 50596 7486
rect 50540 7422 50542 7474
rect 50594 7422 50596 7474
rect 50540 7252 50596 7422
rect 50540 7186 50596 7196
rect 51100 7362 51156 7374
rect 51100 7310 51102 7362
rect 51154 7310 51156 7362
rect 51100 7252 51156 7310
rect 51156 7196 51268 7252
rect 51100 7186 51156 7196
rect 50204 6916 50260 6926
rect 50092 6914 50260 6916
rect 50092 6862 50206 6914
rect 50258 6862 50260 6914
rect 50092 6860 50260 6862
rect 50204 6850 50260 6860
rect 48076 6580 48132 6590
rect 48300 6580 48356 6636
rect 49532 6692 49588 6702
rect 49588 6636 49812 6692
rect 49532 6598 49588 6636
rect 48076 6578 48356 6580
rect 48076 6526 48078 6578
rect 48130 6526 48356 6578
rect 48076 6524 48356 6526
rect 48412 6578 48468 6590
rect 48412 6526 48414 6578
rect 48466 6526 48468 6578
rect 47516 6466 47572 6478
rect 47516 6414 47518 6466
rect 47570 6414 47572 6466
rect 47516 6020 47572 6414
rect 48076 6468 48132 6524
rect 48076 6402 48132 6412
rect 47516 5954 47572 5964
rect 47628 5796 47684 5806
rect 46956 5234 47124 5236
rect 46956 5182 46958 5234
rect 47010 5182 47124 5234
rect 46956 5180 47124 5182
rect 47404 5794 47684 5796
rect 47404 5742 47630 5794
rect 47682 5742 47684 5794
rect 47404 5740 47684 5742
rect 46956 5170 47012 5180
rect 46732 3602 46788 3612
rect 45276 3378 45332 3388
rect 45836 3444 45892 3454
rect 46396 3444 46452 3454
rect 45836 3442 46452 3444
rect 45836 3390 45838 3442
rect 45890 3390 46398 3442
rect 46450 3390 46452 3442
rect 45836 3388 46452 3390
rect 45836 3378 45892 3388
rect 46060 800 46116 3388
rect 46396 3378 46452 3388
rect 47404 800 47460 5740
rect 47628 5730 47684 5740
rect 48412 5460 48468 6526
rect 49420 6578 49476 6590
rect 49420 6526 49422 6578
rect 49474 6526 49476 6578
rect 48748 5908 48804 5918
rect 48748 5814 48804 5852
rect 49084 5908 49140 5918
rect 48412 5394 48468 5404
rect 48860 5460 48916 5470
rect 48076 5124 48132 5134
rect 48076 5030 48132 5068
rect 48636 5124 48692 5134
rect 48636 5030 48692 5068
rect 48524 4900 48580 4910
rect 48300 4898 48580 4900
rect 48300 4846 48526 4898
rect 48578 4846 48580 4898
rect 48300 4844 48580 4846
rect 48300 4562 48356 4844
rect 48524 4834 48580 4844
rect 48300 4510 48302 4562
rect 48354 4510 48356 4562
rect 48300 4498 48356 4510
rect 48860 4562 48916 5404
rect 49084 5346 49140 5852
rect 49420 5908 49476 6526
rect 49420 5842 49476 5852
rect 49756 6132 49812 6636
rect 51212 6690 51268 7196
rect 51212 6638 51214 6690
rect 51266 6638 51268 6690
rect 51212 6626 51268 6638
rect 50540 6580 50596 6590
rect 50540 6486 50596 6524
rect 49756 5906 49812 6076
rect 50316 6468 50372 6478
rect 50316 6130 50372 6412
rect 50316 6078 50318 6130
rect 50370 6078 50372 6130
rect 50316 6066 50372 6078
rect 51100 6132 51156 6142
rect 51100 6038 51156 6076
rect 49756 5854 49758 5906
rect 49810 5854 49812 5906
rect 49756 5842 49812 5854
rect 49084 5294 49086 5346
rect 49138 5294 49140 5346
rect 49084 5282 49140 5294
rect 49868 5124 49924 5134
rect 49868 5010 49924 5068
rect 49868 4958 49870 5010
rect 49922 4958 49924 5010
rect 49868 4946 49924 4958
rect 48860 4510 48862 4562
rect 48914 4510 48916 4562
rect 48860 4498 48916 4510
rect 49644 4452 49700 4462
rect 49196 4450 49700 4452
rect 49196 4398 49646 4450
rect 49698 4398 49700 4450
rect 49196 4396 49700 4398
rect 47516 3668 47572 3678
rect 47516 3574 47572 3612
rect 48860 3444 48916 3454
rect 48860 3350 48916 3388
rect 49196 3442 49252 4396
rect 49644 4386 49700 4396
rect 50764 4228 50820 4238
rect 50764 4134 50820 4172
rect 51436 3668 51492 16828
rect 51548 7476 51604 7486
rect 51548 7382 51604 7420
rect 52108 6580 52164 6590
rect 52108 6486 52164 6524
rect 51548 6468 51604 6478
rect 52444 6468 52500 6478
rect 51548 4562 51604 6412
rect 52220 6466 52500 6468
rect 52220 6414 52446 6466
rect 52498 6414 52500 6466
rect 52220 6412 52500 6414
rect 51772 5796 51828 5806
rect 51548 4510 51550 4562
rect 51602 4510 51604 4562
rect 51548 4498 51604 4510
rect 51660 5794 51828 5796
rect 51660 5742 51774 5794
rect 51826 5742 51828 5794
rect 51660 5740 51828 5742
rect 51548 3668 51604 3678
rect 51436 3666 51604 3668
rect 51436 3614 51550 3666
rect 51602 3614 51604 3666
rect 51436 3612 51604 3614
rect 51548 3602 51604 3612
rect 49196 3390 49198 3442
rect 49250 3390 49252 3442
rect 49196 2548 49252 3390
rect 49868 3444 49924 3454
rect 50428 3444 50484 3454
rect 49868 3442 50484 3444
rect 49868 3390 49870 3442
rect 49922 3390 50430 3442
rect 50482 3390 50484 3442
rect 49868 3388 50484 3390
rect 49868 3378 49924 3388
rect 48748 2492 49252 2548
rect 48748 800 48804 2492
rect 50092 800 50148 3388
rect 50428 3378 50484 3388
rect 51660 980 51716 5740
rect 51772 5730 51828 5740
rect 52220 5122 52276 6412
rect 52444 6402 52500 6412
rect 52892 5908 52948 5918
rect 52892 5814 52948 5852
rect 52220 5070 52222 5122
rect 52274 5070 52276 5122
rect 52220 5058 52276 5070
rect 52556 5796 52612 5806
rect 52556 5236 52612 5740
rect 52556 5122 52612 5180
rect 52556 5070 52558 5122
rect 52610 5070 52612 5122
rect 52556 5058 52612 5070
rect 53004 5012 53060 20132
rect 53676 12852 53732 34636
rect 54124 34244 54180 34254
rect 54124 34150 54180 34188
rect 53900 33460 53956 33470
rect 53900 33366 53956 33404
rect 53676 12786 53732 12796
rect 54236 32116 54292 32126
rect 53340 5908 53396 5918
rect 53340 5814 53396 5852
rect 53564 5348 53620 5358
rect 53564 5234 53620 5292
rect 53564 5182 53566 5234
rect 53618 5182 53620 5234
rect 53564 5170 53620 5182
rect 54124 5348 54180 5358
rect 54124 5234 54180 5292
rect 54124 5182 54126 5234
rect 54178 5182 54180 5234
rect 53452 5124 53508 5134
rect 53452 5030 53508 5068
rect 54124 5124 54180 5182
rect 54124 5058 54180 5068
rect 53004 4946 53060 4956
rect 53116 4452 53172 4462
rect 52780 4450 53172 4452
rect 52780 4398 53118 4450
rect 53170 4398 53172 4450
rect 52780 4396 53172 4398
rect 52556 4228 52612 4238
rect 52780 4228 52836 4396
rect 53116 4386 53172 4396
rect 52556 4226 52836 4228
rect 52556 4174 52558 4226
rect 52610 4174 52836 4226
rect 52556 4172 52836 4174
rect 52556 4162 52612 4172
rect 51436 924 51716 980
rect 51436 800 51492 924
rect 52780 800 52836 4172
rect 54236 4226 54292 32060
rect 54348 22596 54404 35532
rect 54460 35522 54516 35532
rect 54572 34244 54628 35644
rect 55356 34916 55412 34926
rect 55356 34822 55412 34860
rect 54572 34178 54628 34188
rect 54460 34130 54516 34142
rect 54460 34078 54462 34130
rect 54514 34078 54516 34130
rect 54460 34020 54516 34078
rect 54908 34020 54964 34030
rect 54460 34018 54964 34020
rect 54460 33966 54910 34018
rect 54962 33966 54964 34018
rect 54460 33964 54964 33966
rect 54348 22530 54404 22540
rect 54908 21364 54964 33964
rect 55692 25732 55748 36542
rect 56252 35700 56308 38108
rect 56588 37044 56644 39200
rect 57484 37044 57540 39200
rect 56588 36988 56868 37044
rect 57484 36988 57764 37044
rect 56442 36876 56706 36886
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56442 36810 56706 36820
rect 56812 35812 56868 36988
rect 57484 36372 57540 36382
rect 57148 36370 57540 36372
rect 57148 36318 57486 36370
rect 57538 36318 57540 36370
rect 57148 36316 57540 36318
rect 56476 35700 56532 35710
rect 56140 35698 56532 35700
rect 56140 35646 56478 35698
rect 56530 35646 56532 35698
rect 56140 35644 56532 35646
rect 56140 34356 56196 35644
rect 56476 35634 56532 35644
rect 56442 35308 56706 35318
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56442 35242 56706 35252
rect 56700 34804 56756 34814
rect 56700 34710 56756 34748
rect 56252 34692 56308 34702
rect 56252 34598 56308 34636
rect 56364 34356 56420 34366
rect 56140 34354 56420 34356
rect 56140 34302 56366 34354
rect 56418 34302 56420 34354
rect 56140 34300 56420 34302
rect 56364 34290 56420 34300
rect 56812 34354 56868 35756
rect 57036 36258 57092 36270
rect 57036 36206 57038 36258
rect 57090 36206 57092 36258
rect 57036 35252 57092 36206
rect 57036 35186 57092 35196
rect 56812 34302 56814 34354
rect 56866 34302 56868 34354
rect 56812 34290 56868 34302
rect 57036 34802 57092 34814
rect 57036 34750 57038 34802
rect 57090 34750 57092 34802
rect 57036 34692 57092 34750
rect 56442 33740 56706 33750
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56442 33674 56706 33684
rect 56442 32172 56706 32182
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56442 32106 56706 32116
rect 56442 30604 56706 30614
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56442 30538 56706 30548
rect 56442 29036 56706 29046
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56442 28970 56706 28980
rect 56442 27468 56706 27478
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56442 27402 56706 27412
rect 56442 25900 56706 25910
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56442 25834 56706 25844
rect 55692 25666 55748 25676
rect 56442 24332 56706 24342
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56442 24266 56706 24276
rect 56442 22764 56706 22774
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56442 22698 56706 22708
rect 54908 21298 54964 21308
rect 56442 21196 56706 21206
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56442 21130 56706 21140
rect 56442 19628 56706 19638
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56442 19562 56706 19572
rect 56442 18060 56706 18070
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56442 17994 56706 18004
rect 57036 17668 57092 34636
rect 57148 33458 57204 36316
rect 57484 36306 57540 36316
rect 57596 35812 57652 35822
rect 57596 35718 57652 35756
rect 57708 35026 57764 36988
rect 58380 36372 58436 39200
rect 58492 36372 58548 36382
rect 58380 36370 58548 36372
rect 58380 36318 58494 36370
rect 58546 36318 58548 36370
rect 58380 36316 58548 36318
rect 57820 36260 57876 36270
rect 57820 36258 57988 36260
rect 57820 36206 57822 36258
rect 57874 36206 57988 36258
rect 57820 36204 57988 36206
rect 57820 36194 57876 36204
rect 57708 34974 57710 35026
rect 57762 34974 57764 35026
rect 57708 34962 57764 34974
rect 57484 34356 57540 34366
rect 57484 34262 57540 34300
rect 57148 33406 57150 33458
rect 57202 33406 57204 33458
rect 57148 32788 57204 33406
rect 57148 32722 57204 32732
rect 57820 34130 57876 34142
rect 57820 34078 57822 34130
rect 57874 34078 57876 34130
rect 57820 33122 57876 34078
rect 57820 33070 57822 33122
rect 57874 33070 57876 33122
rect 57036 17602 57092 17612
rect 56442 16492 56706 16502
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56442 16426 56706 16436
rect 56442 14924 56706 14934
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56442 14858 56706 14868
rect 57820 14308 57876 33070
rect 57932 26292 57988 36204
rect 58268 34020 58324 34030
rect 58268 33458 58324 33964
rect 58492 33796 58548 36316
rect 59276 35812 59332 39200
rect 59724 36594 59780 36606
rect 59724 36542 59726 36594
rect 59778 36542 59780 36594
rect 59500 36148 59556 36158
rect 59500 35922 59556 36092
rect 59500 35870 59502 35922
rect 59554 35870 59556 35922
rect 59500 35858 59556 35870
rect 59276 35756 59444 35812
rect 58940 35588 58996 35598
rect 58940 35586 59108 35588
rect 58940 35534 58942 35586
rect 58994 35534 59108 35586
rect 58940 35532 59108 35534
rect 58940 35522 58996 35532
rect 58716 34914 58772 34926
rect 58716 34862 58718 34914
rect 58770 34862 58772 34914
rect 58604 34130 58660 34142
rect 58604 34078 58606 34130
rect 58658 34078 58660 34130
rect 58604 34020 58660 34078
rect 58604 33954 58660 33964
rect 58492 33730 58548 33740
rect 58268 33406 58270 33458
rect 58322 33406 58324 33458
rect 58268 33394 58324 33406
rect 58716 33572 58772 34862
rect 58716 31948 58772 33516
rect 58940 34242 58996 34254
rect 58940 34190 58942 34242
rect 58994 34190 58996 34242
rect 57932 26226 57988 26236
rect 58604 31892 58772 31948
rect 58828 32564 58884 32574
rect 58604 23156 58660 31892
rect 58604 23090 58660 23100
rect 58828 20188 58884 32508
rect 58940 31668 58996 34190
rect 58940 31602 58996 31612
rect 59052 30212 59108 35532
rect 59388 35028 59444 35756
rect 59500 35028 59556 35038
rect 59388 35026 59556 35028
rect 59388 34974 59502 35026
rect 59554 34974 59556 35026
rect 59388 34972 59556 34974
rect 59500 34962 59556 34972
rect 59500 34804 59556 34814
rect 59500 34018 59556 34748
rect 59500 33966 59502 34018
rect 59554 33966 59556 34018
rect 59500 33908 59556 33966
rect 59500 33842 59556 33852
rect 59612 33796 59668 33806
rect 59164 33572 59220 33582
rect 59164 33458 59220 33516
rect 59164 33406 59166 33458
rect 59218 33406 59220 33458
rect 59164 33394 59220 33406
rect 59612 33458 59668 33740
rect 59612 33406 59614 33458
rect 59666 33406 59668 33458
rect 59612 33394 59668 33406
rect 59052 30146 59108 30156
rect 59724 26852 59780 36542
rect 60172 35812 60228 39200
rect 61068 36596 61124 39200
rect 61068 36540 61460 36596
rect 60844 36372 60900 36382
rect 60844 36278 60900 36316
rect 61292 36258 61348 36270
rect 61292 36206 61294 36258
rect 61346 36206 61348 36258
rect 60508 35812 60564 35822
rect 60172 35810 60564 35812
rect 60172 35758 60510 35810
rect 60562 35758 60564 35810
rect 60172 35756 60564 35758
rect 59836 35698 59892 35710
rect 59836 35646 59838 35698
rect 59890 35646 59892 35698
rect 59836 34804 59892 35646
rect 59836 34738 59892 34748
rect 59724 26786 59780 26796
rect 59836 34018 59892 34030
rect 59836 33966 59838 34018
rect 59890 33966 59892 34018
rect 59836 33236 59892 33966
rect 60172 33458 60228 35756
rect 60508 35746 60564 35756
rect 60620 34914 60676 34926
rect 60620 34862 60622 34914
rect 60674 34862 60676 34914
rect 60172 33406 60174 33458
rect 60226 33406 60228 33458
rect 60172 33394 60228 33406
rect 60396 34130 60452 34142
rect 60396 34078 60398 34130
rect 60450 34078 60452 34130
rect 60396 33236 60452 34078
rect 60620 33460 60676 34862
rect 61292 34916 61348 36206
rect 61292 34850 61348 34860
rect 60732 34244 60788 34254
rect 60732 34242 60900 34244
rect 60732 34190 60734 34242
rect 60786 34190 60900 34242
rect 60732 34188 60900 34190
rect 60732 34178 60788 34188
rect 60732 33460 60788 33470
rect 60620 33458 60788 33460
rect 60620 33406 60734 33458
rect 60786 33406 60788 33458
rect 60620 33404 60788 33406
rect 59836 33180 60452 33236
rect 58828 20132 58996 20188
rect 57820 14242 57876 14252
rect 58044 14420 58100 14430
rect 56442 13356 56706 13366
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56442 13290 56706 13300
rect 56442 11788 56706 11798
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56442 11722 56706 11732
rect 56442 10220 56706 10230
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56442 10154 56706 10164
rect 56442 8652 56706 8662
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56442 8586 56706 8596
rect 56442 7084 56706 7094
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56442 7018 56706 7028
rect 56476 5796 56532 5806
rect 56252 5794 56532 5796
rect 56252 5742 56478 5794
rect 56530 5742 56532 5794
rect 56252 5740 56532 5742
rect 54460 5236 54516 5246
rect 54460 5142 54516 5180
rect 55692 5012 55748 5022
rect 55020 4564 55076 4574
rect 55020 4470 55076 4508
rect 55580 4228 55636 4238
rect 54236 4174 54238 4226
rect 54290 4174 54292 4226
rect 54236 4162 54292 4174
rect 55468 4226 55636 4228
rect 55468 4174 55582 4226
rect 55634 4174 55636 4226
rect 55468 4172 55636 4174
rect 53900 3444 53956 3454
rect 54460 3444 54516 3454
rect 53900 3442 54516 3444
rect 53900 3390 53902 3442
rect 53954 3390 54462 3442
rect 54514 3390 54516 3442
rect 53900 3388 54516 3390
rect 53900 3378 53956 3388
rect 54124 800 54180 3388
rect 54460 3378 54516 3388
rect 55468 800 55524 4172
rect 55580 4162 55636 4172
rect 55692 3666 55748 4956
rect 55692 3614 55694 3666
rect 55746 3614 55748 3666
rect 55692 3602 55748 3614
rect 55916 4900 55972 4910
rect 56252 4900 56308 5740
rect 56476 5730 56532 5740
rect 57484 5796 57540 5806
rect 57484 5794 57652 5796
rect 57484 5742 57486 5794
rect 57538 5742 57652 5794
rect 57484 5740 57652 5742
rect 57484 5730 57540 5740
rect 56442 5516 56706 5526
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56442 5450 56706 5460
rect 56476 5010 56532 5022
rect 56476 4958 56478 5010
rect 56530 4958 56532 5010
rect 56476 4900 56532 4958
rect 55916 4898 56532 4900
rect 55916 4846 55918 4898
rect 55970 4846 56532 4898
rect 55916 4844 56532 4846
rect 56812 4900 56868 4910
rect 55916 3332 55972 4844
rect 56812 4806 56868 4844
rect 57260 4900 57316 4910
rect 57260 4806 57316 4844
rect 56476 4564 56532 4574
rect 56476 4338 56532 4508
rect 56476 4286 56478 4338
rect 56530 4286 56532 4338
rect 56476 4274 56532 4286
rect 56812 4452 56868 4462
rect 56442 3948 56706 3958
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56442 3882 56706 3892
rect 55916 3266 55972 3276
rect 56700 3442 56756 3454
rect 56700 3390 56702 3442
rect 56754 3390 56756 3442
rect 56700 3332 56756 3390
rect 56700 3266 56756 3276
rect 56812 800 56868 4396
rect 57596 4452 57652 5740
rect 57820 5124 57876 5134
rect 57820 5010 57876 5068
rect 57820 4958 57822 5010
rect 57874 4958 57876 5010
rect 57820 4946 57876 4958
rect 57596 4358 57652 4396
rect 57036 4004 57092 4014
rect 57036 3330 57092 3948
rect 58044 3668 58100 14364
rect 58156 5010 58212 5022
rect 58156 4958 58158 5010
rect 58210 4958 58212 5010
rect 58156 4900 58212 4958
rect 58156 4834 58212 4844
rect 58828 4898 58884 4910
rect 58828 4846 58830 4898
rect 58882 4846 58884 4898
rect 58828 4004 58884 4846
rect 58940 4226 58996 20132
rect 59836 10948 59892 33180
rect 60396 31108 60452 31118
rect 60396 30324 60452 31052
rect 60732 30996 60788 33404
rect 60732 30930 60788 30940
rect 60844 30884 60900 34188
rect 61404 34242 61460 36540
rect 61628 36372 61684 36382
rect 61964 36372 62020 39200
rect 62524 37716 62580 37726
rect 62300 36372 62356 36382
rect 61628 36370 61908 36372
rect 61628 36318 61630 36370
rect 61682 36318 61908 36370
rect 61628 36316 61908 36318
rect 61964 36370 62356 36372
rect 61964 36318 62302 36370
rect 62354 36318 62356 36370
rect 61964 36316 62356 36318
rect 61628 36306 61684 36316
rect 61404 34190 61406 34242
rect 61458 34190 61460 34242
rect 61404 34178 61460 34190
rect 61628 35586 61684 35598
rect 61628 35534 61630 35586
rect 61682 35534 61684 35586
rect 61516 33346 61572 33358
rect 61516 33294 61518 33346
rect 61570 33294 61572 33346
rect 61516 32676 61572 33294
rect 61516 32610 61572 32620
rect 60844 30818 60900 30828
rect 60396 23268 60452 30268
rect 61628 24164 61684 35534
rect 61740 34914 61796 34926
rect 61740 34862 61742 34914
rect 61794 34862 61796 34914
rect 61740 30324 61796 34862
rect 61852 32450 61908 36316
rect 62300 35252 62356 36316
rect 62300 35186 62356 35196
rect 62412 35476 62468 35486
rect 62188 34914 62244 34926
rect 62188 34862 62190 34914
rect 62242 34862 62244 34914
rect 61964 33908 62020 33918
rect 61964 33124 62020 33852
rect 62076 33348 62132 33358
rect 62188 33348 62244 34862
rect 62412 34468 62468 35420
rect 62412 34402 62468 34412
rect 62524 34132 62580 37660
rect 62636 35588 62692 35598
rect 62636 35494 62692 35532
rect 62860 35028 62916 39200
rect 63644 37828 63700 37838
rect 63644 36594 63700 37772
rect 63644 36542 63646 36594
rect 63698 36542 63700 36594
rect 63644 36530 63700 36542
rect 63644 35812 63700 35822
rect 63756 35812 63812 39200
rect 63532 35810 63812 35812
rect 63532 35758 63646 35810
rect 63698 35758 63812 35810
rect 63532 35756 63812 35758
rect 64092 37492 64148 37502
rect 63084 35588 63140 35598
rect 62972 35028 63028 35038
rect 62860 35026 63028 35028
rect 62860 34974 62974 35026
rect 63026 34974 63028 35026
rect 62860 34972 63028 34974
rect 62972 34962 63028 34972
rect 62524 34130 62916 34132
rect 62524 34078 62526 34130
rect 62578 34078 62916 34130
rect 62524 34076 62916 34078
rect 62524 34066 62580 34076
rect 62636 33348 62692 33358
rect 62076 33346 62692 33348
rect 62076 33294 62078 33346
rect 62130 33294 62638 33346
rect 62690 33294 62692 33346
rect 62076 33292 62692 33294
rect 62076 33282 62132 33292
rect 61964 33068 62244 33124
rect 61852 32398 61854 32450
rect 61906 32398 61908 32450
rect 61852 32228 61908 32398
rect 61852 32162 61908 32172
rect 61740 30258 61796 30268
rect 62188 24388 62244 33068
rect 62300 32788 62356 33292
rect 62636 33282 62692 33292
rect 62300 32656 62356 32732
rect 62860 32786 62916 34076
rect 62860 32734 62862 32786
rect 62914 32734 62916 32786
rect 62860 32722 62916 32734
rect 62972 33236 63028 33246
rect 63084 33236 63140 35532
rect 62972 33234 63140 33236
rect 62972 33182 62974 33234
rect 63026 33182 63140 33234
rect 62972 33180 63140 33182
rect 63308 34130 63364 34142
rect 63308 34078 63310 34130
rect 63362 34078 63364 34130
rect 62972 31780 63028 33180
rect 63308 33124 63364 34078
rect 63420 33124 63476 33134
rect 63308 33068 63420 33124
rect 63196 32788 63252 32798
rect 63308 32788 63364 33068
rect 63420 32992 63476 33068
rect 63252 32732 63364 32788
rect 63196 32694 63252 32732
rect 63532 31948 63588 35756
rect 63644 35746 63700 35756
rect 64092 34914 64148 37436
rect 64652 36820 64708 39200
rect 65436 37492 65492 37502
rect 64652 36764 65044 36820
rect 64764 36594 64820 36606
rect 64764 36542 64766 36594
rect 64818 36542 64820 36594
rect 64092 34862 64094 34914
rect 64146 34862 64148 34914
rect 64092 34850 64148 34862
rect 64652 35586 64708 35598
rect 64652 35534 64654 35586
rect 64706 35534 64708 35586
rect 63644 34242 63700 34254
rect 63644 34190 63646 34242
rect 63698 34190 63700 34242
rect 63644 33908 63700 34190
rect 64540 34242 64596 34254
rect 64540 34190 64542 34242
rect 64594 34190 64596 34242
rect 64316 34130 64372 34142
rect 64316 34078 64318 34130
rect 64370 34078 64372 34130
rect 63644 33842 63700 33852
rect 63980 33908 64036 33918
rect 63308 31892 63588 31948
rect 63868 33124 63924 33134
rect 63308 31826 63364 31836
rect 62972 31714 63028 31724
rect 62188 24322 62244 24332
rect 62636 25172 62692 25182
rect 61628 24098 61684 24108
rect 60396 23202 60452 23212
rect 61740 23044 61796 23054
rect 61740 20188 61796 22988
rect 61740 20132 62020 20188
rect 59836 10882 59892 10892
rect 60844 6468 60900 6478
rect 59948 6356 60004 6366
rect 59948 6130 60004 6300
rect 59948 6078 59950 6130
rect 60002 6078 60004 6130
rect 59948 6066 60004 6078
rect 60396 6356 60452 6366
rect 59612 5234 59668 5246
rect 59612 5182 59614 5234
rect 59666 5182 59668 5234
rect 59500 4452 59556 4462
rect 58940 4174 58942 4226
rect 58994 4174 58996 4226
rect 58940 4162 58996 4174
rect 59388 4450 59556 4452
rect 59388 4398 59502 4450
rect 59554 4398 59556 4450
rect 59388 4396 59556 4398
rect 58828 3938 58884 3948
rect 58044 3602 58100 3612
rect 59388 3556 59444 4396
rect 59500 4386 59556 4396
rect 59612 3892 59668 5182
rect 60396 5122 60452 6300
rect 60844 6132 60900 6412
rect 60844 6000 60900 6076
rect 61852 6466 61908 6478
rect 61852 6414 61854 6466
rect 61906 6414 61908 6466
rect 61516 6020 61572 6030
rect 61180 6018 61572 6020
rect 61180 5966 61518 6018
rect 61570 5966 61572 6018
rect 61180 5964 61572 5966
rect 60396 5070 60398 5122
rect 60450 5070 60452 5122
rect 60396 5058 60452 5070
rect 60508 5794 60564 5806
rect 60508 5742 60510 5794
rect 60562 5742 60564 5794
rect 60508 5682 60564 5742
rect 60508 5630 60510 5682
rect 60562 5630 60564 5682
rect 59836 4338 59892 4350
rect 59836 4286 59838 4338
rect 59890 4286 59892 4338
rect 59836 4004 59892 4286
rect 59836 3938 59892 3948
rect 59388 3490 59444 3500
rect 59500 3836 59668 3892
rect 57932 3444 57988 3454
rect 58492 3444 58548 3454
rect 57932 3442 58548 3444
rect 57932 3390 57934 3442
rect 57986 3390 58494 3442
rect 58546 3390 58548 3442
rect 57932 3388 58548 3390
rect 57932 3378 57988 3388
rect 57036 3278 57038 3330
rect 57090 3278 57092 3330
rect 57036 3266 57092 3278
rect 58156 800 58212 3388
rect 58492 3378 58548 3388
rect 59500 800 59556 3836
rect 59612 3668 59668 3678
rect 59612 3574 59668 3612
rect 60508 3332 60564 5630
rect 61180 5682 61236 5964
rect 61516 5954 61572 5964
rect 61180 5630 61182 5682
rect 61234 5630 61236 5682
rect 61180 5618 61236 5630
rect 60620 5236 60676 5246
rect 60620 4564 60676 5180
rect 61740 5124 61796 5134
rect 60620 4562 61124 4564
rect 60620 4510 60622 4562
rect 60674 4510 61124 4562
rect 60620 4508 61124 4510
rect 60620 4498 60676 4508
rect 61068 4338 61124 4508
rect 61068 4286 61070 4338
rect 61122 4286 61124 4338
rect 61068 4274 61124 4286
rect 61740 4338 61796 5068
rect 61740 4286 61742 4338
rect 61794 4286 61796 4338
rect 61740 4274 61796 4286
rect 60844 3556 60900 3566
rect 60844 3462 60900 3500
rect 61740 3444 61796 3454
rect 61852 3444 61908 6414
rect 61964 3892 62020 20132
rect 62524 7586 62580 7598
rect 62524 7534 62526 7586
rect 62578 7534 62580 7586
rect 62300 6690 62356 6702
rect 62300 6638 62302 6690
rect 62354 6638 62356 6690
rect 61964 3826 62020 3836
rect 62188 5234 62244 5246
rect 62188 5182 62190 5234
rect 62242 5182 62244 5234
rect 62188 5012 62244 5182
rect 62300 5236 62356 6638
rect 62300 5170 62356 5180
rect 62524 5124 62580 7534
rect 62636 5794 62692 25116
rect 63868 20188 63924 33068
rect 63980 32786 64036 33852
rect 63980 32734 63982 32786
rect 64034 32734 64036 32786
rect 63980 32722 64036 32734
rect 64316 33122 64372 34078
rect 64316 33070 64318 33122
rect 64370 33070 64372 33122
rect 64316 27748 64372 33070
rect 64428 33572 64484 33582
rect 64428 32450 64484 33516
rect 64540 32788 64596 34190
rect 64652 33236 64708 35534
rect 64764 35476 64820 36542
rect 64876 35476 64932 35486
rect 64764 35420 64876 35476
rect 64876 34914 64932 35420
rect 64876 34862 64878 34914
rect 64930 34862 64932 34914
rect 64876 34850 64932 34862
rect 64764 34802 64820 34814
rect 64764 34750 64766 34802
rect 64818 34750 64820 34802
rect 64764 33572 64820 34750
rect 64764 33506 64820 33516
rect 64988 33458 65044 36764
rect 65100 36482 65156 36494
rect 65100 36430 65102 36482
rect 65154 36430 65156 36482
rect 65100 33908 65156 36430
rect 65100 33842 65156 33852
rect 64988 33406 64990 33458
rect 65042 33406 65044 33458
rect 64988 33394 65044 33406
rect 64652 33180 65044 33236
rect 64540 32722 64596 32732
rect 64428 32398 64430 32450
rect 64482 32398 64484 32450
rect 64428 32004 64484 32398
rect 64428 31938 64484 31948
rect 64876 31892 64932 31902
rect 64876 31798 64932 31836
rect 64988 29540 65044 33180
rect 65436 32786 65492 37436
rect 65548 36372 65604 39200
rect 65548 36306 65604 36316
rect 65660 37940 65716 37950
rect 65660 35810 65716 37884
rect 65884 36372 65940 36382
rect 65884 36278 65940 36316
rect 65660 35758 65662 35810
rect 65714 35758 65716 35810
rect 65548 35698 65604 35710
rect 65548 35646 65550 35698
rect 65602 35646 65604 35698
rect 65548 35476 65604 35646
rect 65548 35410 65604 35420
rect 65660 35364 65716 35758
rect 66332 35476 66388 35486
rect 66332 35382 66388 35420
rect 66220 35364 66276 35374
rect 65660 35308 65828 35364
rect 65548 34916 65604 34926
rect 65548 34914 65716 34916
rect 65548 34862 65550 34914
rect 65602 34862 65716 34914
rect 65548 34860 65716 34862
rect 65548 34850 65604 34860
rect 65660 34020 65716 34860
rect 65660 33926 65716 33964
rect 65436 32734 65438 32786
rect 65490 32734 65492 32786
rect 65436 32722 65492 32734
rect 65772 32786 65828 35308
rect 65884 34690 65940 34702
rect 65884 34638 65886 34690
rect 65938 34638 65940 34690
rect 65884 34356 65940 34638
rect 65884 34300 66164 34356
rect 65884 33346 65940 33358
rect 65884 33294 65886 33346
rect 65938 33294 65940 33346
rect 65884 33124 65940 33294
rect 65884 33058 65940 33068
rect 65996 33348 66052 33358
rect 65772 32734 65774 32786
rect 65826 32734 65828 32786
rect 65772 32722 65828 32734
rect 65996 31948 66052 33292
rect 64988 29474 65044 29484
rect 65884 31892 66052 31948
rect 64316 27682 64372 27692
rect 65884 20188 65940 31892
rect 66108 20188 66164 34300
rect 66220 32786 66276 35308
rect 66444 34018 66500 39200
rect 67228 38388 67284 38398
rect 66556 36932 66612 36942
rect 66556 34356 66612 36876
rect 67228 36594 67284 38332
rect 67228 36542 67230 36594
rect 67282 36542 67284 36594
rect 67228 36530 67284 36542
rect 67340 36596 67396 39200
rect 68012 37604 68068 37614
rect 67676 36596 67732 36606
rect 67340 36594 67732 36596
rect 67340 36542 67678 36594
rect 67730 36542 67732 36594
rect 67340 36540 67732 36542
rect 67676 35810 67732 36540
rect 67676 35758 67678 35810
rect 67730 35758 67732 35810
rect 67676 35746 67732 35758
rect 66556 34290 66612 34300
rect 66668 35474 66724 35486
rect 66668 35422 66670 35474
rect 66722 35422 66724 35474
rect 66444 33966 66446 34018
rect 66498 33966 66500 34018
rect 66444 33954 66500 33966
rect 66668 33348 66724 35422
rect 67004 35476 67060 35486
rect 66780 34692 66836 34702
rect 66780 34598 66836 34636
rect 66668 33282 66724 33292
rect 66220 32734 66222 32786
rect 66274 32734 66276 32786
rect 66220 32722 66276 32734
rect 66668 33124 66724 33134
rect 66668 32004 66724 33068
rect 67004 32788 67060 35420
rect 67116 34804 67172 34814
rect 67116 33458 67172 34748
rect 67340 34804 67396 34814
rect 67340 34710 67396 34748
rect 67900 34802 67956 34814
rect 67900 34750 67902 34802
rect 67954 34750 67956 34802
rect 67900 34692 67956 34750
rect 68012 34692 68068 37548
rect 68124 35140 68180 35150
rect 68124 35046 68180 35084
rect 68012 34636 68180 34692
rect 67900 34626 67956 34636
rect 68124 34242 68180 34636
rect 68236 34356 68292 39200
rect 69020 37604 69076 37614
rect 68460 36596 68516 36606
rect 68460 36502 68516 36540
rect 68908 36372 68964 36382
rect 68908 35588 68964 36316
rect 68908 35522 68964 35532
rect 69020 35586 69076 37548
rect 69132 36596 69188 39200
rect 69916 38500 69972 38510
rect 69132 36372 69188 36540
rect 69804 37940 69860 37950
rect 69468 36372 69524 36382
rect 69132 36370 69524 36372
rect 69132 36318 69470 36370
rect 69522 36318 69524 36370
rect 69132 36316 69524 36318
rect 69468 36306 69524 36316
rect 69692 36260 69748 36270
rect 69692 35924 69748 36204
rect 69692 35792 69748 35868
rect 69020 35534 69022 35586
rect 69074 35534 69076 35586
rect 69020 35522 69076 35534
rect 69356 35140 69412 35150
rect 68236 34290 68292 34300
rect 68460 34690 68516 34702
rect 68460 34638 68462 34690
rect 68514 34638 68516 34690
rect 68124 34190 68126 34242
rect 68178 34190 68180 34242
rect 67340 34132 67396 34142
rect 67340 34038 67396 34076
rect 68124 33908 68180 34190
rect 67116 33406 67118 33458
rect 67170 33406 67172 33458
rect 67116 33394 67172 33406
rect 67676 33852 68180 33908
rect 68236 34132 68292 34142
rect 67676 33458 67732 33852
rect 67676 33406 67678 33458
rect 67730 33406 67732 33458
rect 67676 33394 67732 33406
rect 68124 33460 68180 33470
rect 68236 33460 68292 34076
rect 68124 33458 68292 33460
rect 68124 33406 68126 33458
rect 68178 33406 68292 33458
rect 68124 33404 68292 33406
rect 68124 33394 68180 33404
rect 67340 33012 67396 33022
rect 67116 32788 67172 32798
rect 67004 32786 67172 32788
rect 67004 32734 67118 32786
rect 67170 32734 67172 32786
rect 67004 32732 67172 32734
rect 67116 32722 67172 32732
rect 67228 32788 67284 32798
rect 67340 32788 67396 32956
rect 67284 32732 67396 32788
rect 67228 32722 67284 32732
rect 66668 31938 66724 31948
rect 63868 20132 64036 20188
rect 62860 8820 62916 8830
rect 62860 7586 62916 8764
rect 63644 8258 63700 8270
rect 63644 8206 63646 8258
rect 63698 8206 63700 8258
rect 63196 8036 63252 8046
rect 63644 8036 63700 8206
rect 63196 8034 63700 8036
rect 63196 7982 63198 8034
rect 63250 7982 63700 8034
rect 63196 7980 63700 7982
rect 63084 7588 63140 7598
rect 62860 7534 62862 7586
rect 62914 7534 62916 7586
rect 62860 7522 62916 7534
rect 62972 7586 63140 7588
rect 62972 7534 63086 7586
rect 63138 7534 63140 7586
rect 62972 7532 63140 7534
rect 62860 6692 62916 6702
rect 62972 6692 63028 7532
rect 63084 7522 63140 7532
rect 62860 6690 63028 6692
rect 62860 6638 62862 6690
rect 62914 6638 63028 6690
rect 62860 6636 63028 6638
rect 62860 6626 62916 6636
rect 62636 5742 62638 5794
rect 62690 5742 62692 5794
rect 62636 5730 62692 5742
rect 62524 5058 62580 5068
rect 62188 3444 62244 4956
rect 63196 5012 63252 7980
rect 63308 7588 63364 7598
rect 63532 7588 63588 7598
rect 63308 7586 63588 7588
rect 63308 7534 63310 7586
rect 63362 7534 63534 7586
rect 63586 7534 63588 7586
rect 63308 7532 63588 7534
rect 63308 7522 63364 7532
rect 63532 7522 63588 7532
rect 63868 7476 63924 7486
rect 63868 7382 63924 7420
rect 63196 4946 63252 4956
rect 63532 5794 63588 5806
rect 63532 5742 63534 5794
rect 63586 5742 63588 5794
rect 61740 3442 62132 3444
rect 61740 3390 61742 3442
rect 61794 3390 62132 3442
rect 61740 3388 62132 3390
rect 61740 3378 61796 3388
rect 60508 3276 60900 3332
rect 60844 800 60900 3276
rect 62076 3220 62132 3388
rect 62188 3378 62244 3388
rect 62076 3164 62244 3220
rect 62188 800 62244 3164
rect 63532 800 63588 5742
rect 63868 3780 63924 3790
rect 63980 3780 64036 20132
rect 65772 20132 65940 20188
rect 65996 20132 66164 20188
rect 64652 9156 64708 9166
rect 64652 9062 64708 9100
rect 64876 9156 64932 9166
rect 64316 8930 64372 8942
rect 64316 8878 64318 8930
rect 64370 8878 64372 8930
rect 64316 8428 64372 8878
rect 64316 8372 64708 8428
rect 64204 8260 64260 8270
rect 64092 8258 64260 8260
rect 64092 8206 64206 8258
rect 64258 8206 64260 8258
rect 64092 8204 64260 8206
rect 64092 6580 64148 8204
rect 64204 8194 64260 8204
rect 64652 7364 64708 8372
rect 64652 7362 64820 7364
rect 64652 7310 64654 7362
rect 64706 7310 64820 7362
rect 64652 7308 64820 7310
rect 64652 7298 64708 7308
rect 64540 7252 64596 7262
rect 64092 6514 64148 6524
rect 64204 7250 64596 7252
rect 64204 7198 64542 7250
rect 64594 7198 64596 7250
rect 64204 7196 64596 7198
rect 64204 4562 64260 7196
rect 64540 7186 64596 7196
rect 64652 6692 64708 6702
rect 64652 5906 64708 6636
rect 64652 5854 64654 5906
rect 64706 5854 64708 5906
rect 64652 5842 64708 5854
rect 64764 5684 64820 7308
rect 64204 4510 64206 4562
rect 64258 4510 64260 4562
rect 64204 4498 64260 4510
rect 64652 5628 64820 5684
rect 64876 5796 64932 9100
rect 65548 8820 65604 8830
rect 65548 8726 65604 8764
rect 65772 8372 65828 20132
rect 65996 9268 66052 20132
rect 65884 9044 65940 9054
rect 65996 9044 66052 9212
rect 67228 9268 67284 9278
rect 67228 9174 67284 9212
rect 65884 9042 66052 9044
rect 65884 8990 65886 9042
rect 65938 8990 66052 9042
rect 65884 8988 66052 8990
rect 66108 9154 66164 9166
rect 66108 9102 66110 9154
rect 66162 9102 66164 9154
rect 65884 8978 65940 8988
rect 65548 7476 65604 7486
rect 65772 7476 65828 8316
rect 66108 7586 66164 9102
rect 66444 9156 66500 9166
rect 66444 9062 66500 9100
rect 68460 8428 68516 34638
rect 68572 34692 68628 34702
rect 68572 34242 68628 34636
rect 68572 34190 68574 34242
rect 68626 34190 68628 34242
rect 68572 34178 68628 34190
rect 68796 34132 68852 34142
rect 68796 34130 69300 34132
rect 68796 34078 68798 34130
rect 68850 34078 69300 34130
rect 68796 34076 69300 34078
rect 68796 34066 68852 34076
rect 69132 33906 69188 33918
rect 69132 33854 69134 33906
rect 69186 33854 69188 33906
rect 69132 20188 69188 33854
rect 69244 33570 69300 34076
rect 69244 33518 69246 33570
rect 69298 33518 69300 33570
rect 69244 33506 69300 33518
rect 69356 33458 69412 35084
rect 69468 34692 69524 34702
rect 69468 34598 69524 34636
rect 69356 33406 69358 33458
rect 69410 33406 69412 33458
rect 69356 33394 69412 33406
rect 69468 34020 69524 34030
rect 69468 30100 69524 33964
rect 69804 33570 69860 37884
rect 69916 35140 69972 38444
rect 70028 37044 70084 39200
rect 70924 38836 70980 39200
rect 70924 38780 71316 38836
rect 71148 38612 71204 38622
rect 70812 38276 70868 38286
rect 70028 36988 70420 37044
rect 69916 35074 69972 35084
rect 70252 35810 70308 35822
rect 70252 35758 70254 35810
rect 70306 35758 70308 35810
rect 69916 34356 69972 34366
rect 69916 34242 69972 34300
rect 69916 34190 69918 34242
rect 69970 34190 69972 34242
rect 69916 34178 69972 34190
rect 69804 33518 69806 33570
rect 69858 33518 69860 33570
rect 69804 33458 69860 33518
rect 69804 33406 69806 33458
rect 69858 33406 69860 33458
rect 69804 33394 69860 33406
rect 70252 33460 70308 35758
rect 70364 35026 70420 36988
rect 70812 36594 70868 38220
rect 70812 36542 70814 36594
rect 70866 36542 70868 36594
rect 70812 36530 70868 36542
rect 70364 34974 70366 35026
rect 70418 34974 70420 35026
rect 70364 34962 70420 34974
rect 70588 35698 70644 35710
rect 70588 35646 70590 35698
rect 70642 35646 70644 35698
rect 70252 33394 70308 33404
rect 70588 33124 70644 35646
rect 71036 34130 71092 34142
rect 71036 34078 71038 34130
rect 71090 34078 71092 34130
rect 71036 34018 71092 34078
rect 71148 34132 71204 38556
rect 71148 34066 71204 34076
rect 71260 35810 71316 38780
rect 71820 37044 71876 39200
rect 72716 39060 72772 39200
rect 73052 39060 73108 39228
rect 72716 39004 73108 39060
rect 73164 37268 73220 37278
rect 71820 36988 72212 37044
rect 71708 36596 71764 36606
rect 71708 36502 71764 36540
rect 71260 35758 71262 35810
rect 71314 35758 71316 35810
rect 71036 33966 71038 34018
rect 71090 33966 71092 34018
rect 71036 33954 71092 33966
rect 71260 33460 71316 35758
rect 72156 35028 72212 36988
rect 72380 36372 72436 36382
rect 72380 36278 72436 36316
rect 73164 36370 73220 37212
rect 73164 36318 73166 36370
rect 73218 36318 73220 36370
rect 73164 36306 73220 36318
rect 72492 36260 72548 36270
rect 72492 36166 72548 36204
rect 72716 36258 72772 36270
rect 72716 36206 72718 36258
rect 72770 36206 72772 36258
rect 72716 35700 72772 36206
rect 73388 35812 73444 39228
rect 73584 39200 73696 40000
rect 74480 39200 74592 40000
rect 75376 39200 75488 40000
rect 76272 39200 76384 40000
rect 77168 39200 77280 40000
rect 78064 39200 78176 40000
rect 78960 39200 79072 40000
rect 79856 39200 79968 40000
rect 80220 39228 80612 39284
rect 73500 37380 73556 37390
rect 73500 36482 73556 37324
rect 73500 36430 73502 36482
rect 73554 36430 73556 36482
rect 73500 36418 73556 36430
rect 73500 35812 73556 35822
rect 72716 35634 72772 35644
rect 72828 35810 73556 35812
rect 72828 35758 73502 35810
rect 73554 35758 73556 35810
rect 72828 35756 73556 35758
rect 72380 35586 72436 35598
rect 72380 35534 72382 35586
rect 72434 35534 72436 35586
rect 72268 35028 72324 35038
rect 72156 35026 72324 35028
rect 72156 34974 72270 35026
rect 72322 34974 72324 35026
rect 72156 34972 72324 34974
rect 72268 34962 72324 34972
rect 71484 34916 71540 34926
rect 71484 34914 71988 34916
rect 71484 34862 71486 34914
rect 71538 34862 71988 34914
rect 71484 34860 71988 34862
rect 71484 34850 71540 34860
rect 71484 34018 71540 34030
rect 71484 33966 71486 34018
rect 71538 33966 71540 34018
rect 71484 33906 71540 33966
rect 71484 33854 71486 33906
rect 71538 33854 71540 33906
rect 71372 33460 71428 33470
rect 71260 33458 71428 33460
rect 71260 33406 71374 33458
rect 71426 33406 71428 33458
rect 71260 33404 71428 33406
rect 71372 33394 71428 33404
rect 70812 33124 70868 33134
rect 70588 33122 70868 33124
rect 70588 33070 70814 33122
rect 70866 33070 70868 33122
rect 70588 33068 70868 33070
rect 70812 32004 70868 33068
rect 70812 31938 70868 31948
rect 69468 30034 69524 30044
rect 71484 28420 71540 33854
rect 71932 34018 71988 34860
rect 71932 33966 71934 34018
rect 71986 33966 71988 34018
rect 71932 31892 71988 33966
rect 71932 31826 71988 31836
rect 72380 28532 72436 35534
rect 72716 34356 72772 34366
rect 72828 34356 72884 35756
rect 73500 35746 73556 35756
rect 73612 35028 73668 39200
rect 73612 34962 73668 34972
rect 73724 37380 73780 37390
rect 73276 34914 73332 34926
rect 73276 34862 73278 34914
rect 73330 34862 73332 34914
rect 73276 34804 73332 34862
rect 73276 34738 73332 34748
rect 73724 34580 73780 37324
rect 74508 36596 74564 39200
rect 74508 36370 74564 36540
rect 74508 36318 74510 36370
rect 74562 36318 74564 36370
rect 74508 36306 74564 36318
rect 75292 38724 75348 38734
rect 74852 36092 75116 36102
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 74852 36026 75116 36036
rect 74732 35812 74788 35822
rect 74508 35028 74564 35038
rect 74508 34934 74564 34972
rect 72716 34354 72884 34356
rect 72716 34302 72718 34354
rect 72770 34302 72884 34354
rect 72716 34300 72884 34302
rect 73612 34524 73780 34580
rect 73836 34914 73892 34926
rect 73836 34862 73838 34914
rect 73890 34862 73892 34914
rect 72716 34290 72772 34300
rect 73500 34132 73556 34142
rect 73500 34038 73556 34076
rect 73612 33460 73668 34524
rect 73724 34356 73780 34366
rect 73836 34356 73892 34862
rect 73724 34354 73892 34356
rect 73724 34302 73726 34354
rect 73778 34302 73892 34354
rect 73724 34300 73892 34302
rect 74172 34916 74228 34926
rect 74172 34354 74228 34860
rect 74172 34302 74174 34354
rect 74226 34302 74228 34354
rect 73724 34290 73780 34300
rect 74172 34132 74228 34302
rect 74732 34354 74788 35756
rect 75292 35812 75348 38668
rect 75292 35746 75348 35756
rect 74844 35588 74900 35598
rect 74844 35494 74900 35532
rect 74852 34524 75116 34534
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 74852 34458 75116 34468
rect 74732 34302 74734 34354
rect 74786 34302 74788 34354
rect 74732 34290 74788 34302
rect 75404 34356 75460 39200
rect 75628 37044 75684 37054
rect 75516 36596 75572 36606
rect 75628 36596 75684 36988
rect 75516 36594 75684 36596
rect 75516 36542 75518 36594
rect 75570 36542 75684 36594
rect 75516 36540 75684 36542
rect 75516 36530 75572 36540
rect 75628 35812 75684 35822
rect 75628 35718 75684 35756
rect 76076 35810 76132 35822
rect 76076 35758 76078 35810
rect 76130 35758 76132 35810
rect 75740 34914 75796 34926
rect 75740 34862 75742 34914
rect 75794 34862 75796 34914
rect 75740 34468 75796 34862
rect 75628 34356 75684 34366
rect 75404 34354 75684 34356
rect 75404 34302 75630 34354
rect 75682 34302 75684 34354
rect 75404 34300 75684 34302
rect 75628 34290 75684 34300
rect 74172 34066 74228 34076
rect 75068 34018 75124 34030
rect 75068 33966 75070 34018
rect 75122 33966 75124 34018
rect 75068 33908 75124 33966
rect 75068 33842 75124 33852
rect 75740 33908 75796 34412
rect 75740 33842 75796 33852
rect 76076 34916 76132 35758
rect 76300 35812 76356 39200
rect 76300 35746 76356 35756
rect 76412 38052 76468 38062
rect 76412 36370 76468 37996
rect 77196 36820 77252 39200
rect 77196 36754 77252 36764
rect 77308 38052 77364 38062
rect 77196 36596 77252 36606
rect 77308 36596 77364 37996
rect 78092 36820 78148 39200
rect 78764 38724 78820 38734
rect 78652 38052 78708 38062
rect 78092 36764 78484 36820
rect 77532 36708 77588 36718
rect 77532 36706 78372 36708
rect 77532 36654 77534 36706
rect 77586 36654 78372 36706
rect 77532 36652 78372 36654
rect 77532 36642 77588 36652
rect 77196 36594 77364 36596
rect 77196 36542 77198 36594
rect 77250 36542 77364 36594
rect 77196 36540 77364 36542
rect 77196 36530 77252 36540
rect 78204 36484 78260 36494
rect 77980 36482 78260 36484
rect 77980 36430 78206 36482
rect 78258 36430 78260 36482
rect 77980 36428 78260 36430
rect 76412 36318 76414 36370
rect 76466 36318 76468 36370
rect 76300 35476 76356 35486
rect 76300 35382 76356 35420
rect 76188 34916 76244 34926
rect 76076 34914 76244 34916
rect 76076 34862 76190 34914
rect 76242 34862 76244 34914
rect 76076 34860 76244 34862
rect 76076 34692 76132 34860
rect 73724 33460 73780 33470
rect 73612 33458 73780 33460
rect 73612 33406 73726 33458
rect 73778 33406 73780 33458
rect 73612 33404 73780 33406
rect 72380 28466 72436 28476
rect 71484 28354 71540 28364
rect 71708 22932 71764 22942
rect 69132 20132 69524 20188
rect 67676 8372 67732 8382
rect 67676 8278 67732 8316
rect 67900 8372 68516 8428
rect 66780 8034 66836 8046
rect 66780 7982 66782 8034
rect 66834 7982 66836 8034
rect 66108 7534 66110 7586
rect 66162 7534 66164 7586
rect 65884 7476 65940 7486
rect 65772 7474 65940 7476
rect 65772 7422 65886 7474
rect 65938 7422 65940 7474
rect 65772 7420 65940 7422
rect 65548 7382 65604 7420
rect 65884 7410 65940 7420
rect 65884 7252 65940 7262
rect 65324 6468 65380 6478
rect 65324 6374 65380 6412
rect 65884 6466 65940 7196
rect 65884 6414 65886 6466
rect 65938 6414 65940 6466
rect 65548 6132 65604 6142
rect 65548 6038 65604 6076
rect 63868 3778 64036 3780
rect 63868 3726 63870 3778
rect 63922 3726 64036 3778
rect 63868 3724 64036 3726
rect 63868 3714 63924 3724
rect 64652 3668 64708 5628
rect 64764 4564 64820 4574
rect 64876 4564 64932 5740
rect 64764 4562 64932 4564
rect 64764 4510 64766 4562
rect 64818 4510 64932 4562
rect 64764 4508 64932 4510
rect 65884 4564 65940 6414
rect 66108 5908 66164 7534
rect 66444 7586 66500 7598
rect 66444 7534 66446 7586
rect 66498 7534 66500 7586
rect 66444 7252 66500 7534
rect 66444 7186 66500 7196
rect 66332 6580 66388 6590
rect 66332 6486 66388 6524
rect 66668 6578 66724 6590
rect 66668 6526 66670 6578
rect 66722 6526 66724 6578
rect 66668 6020 66724 6526
rect 66668 5954 66724 5964
rect 66108 5814 66164 5852
rect 66668 5794 66724 5806
rect 66668 5742 66670 5794
rect 66722 5742 66724 5794
rect 66668 5684 66724 5742
rect 66668 5618 66724 5628
rect 66780 5572 66836 7982
rect 67340 8034 67396 8046
rect 67340 7982 67342 8034
rect 67394 7982 67396 8034
rect 67228 7362 67284 7374
rect 67228 7310 67230 7362
rect 67282 7310 67284 7362
rect 67228 7252 67284 7310
rect 67228 7186 67284 7196
rect 67340 6804 67396 7982
rect 67788 7588 67844 7598
rect 67340 6738 67396 6748
rect 67676 7586 67844 7588
rect 67676 7534 67790 7586
rect 67842 7534 67844 7586
rect 67676 7532 67844 7534
rect 67564 6580 67620 6590
rect 67564 6356 67620 6524
rect 67564 6290 67620 6300
rect 67340 6020 67396 6030
rect 66780 5506 66836 5516
rect 67004 5906 67060 5918
rect 67004 5854 67006 5906
rect 67058 5854 67060 5906
rect 67004 5796 67060 5854
rect 67116 5796 67172 5806
rect 67004 5740 67116 5796
rect 67004 5236 67060 5740
rect 67116 5730 67172 5740
rect 67340 5346 67396 5964
rect 67676 5906 67732 7532
rect 67788 7522 67844 7532
rect 67900 6804 67956 8372
rect 68236 8036 68292 8046
rect 68236 8034 68628 8036
rect 68236 7982 68238 8034
rect 68290 7982 68628 8034
rect 68236 7980 68628 7982
rect 68236 7970 68292 7980
rect 68124 7476 68180 7486
rect 68124 7474 68516 7476
rect 68124 7422 68126 7474
rect 68178 7422 68516 7474
rect 68124 7420 68516 7422
rect 68124 7410 68180 7420
rect 68124 6916 68180 6926
rect 68124 6822 68180 6860
rect 68460 6914 68516 7420
rect 68460 6862 68462 6914
rect 68514 6862 68516 6914
rect 68460 6850 68516 6862
rect 67676 5854 67678 5906
rect 67730 5854 67732 5906
rect 67676 5842 67732 5854
rect 67788 6748 67956 6804
rect 67788 5684 67844 6748
rect 68236 6692 68292 6702
rect 67340 5294 67342 5346
rect 67394 5294 67396 5346
rect 67340 5282 67396 5294
rect 67676 5348 67732 5358
rect 67788 5348 67844 5628
rect 67676 5346 67844 5348
rect 67676 5294 67678 5346
rect 67730 5294 67844 5346
rect 67676 5292 67844 5294
rect 67900 6578 67956 6590
rect 67900 6526 67902 6578
rect 67954 6526 67956 6578
rect 67900 5908 67956 6526
rect 67676 5282 67732 5292
rect 67004 5170 67060 5180
rect 64764 4498 64820 4508
rect 65884 4498 65940 4508
rect 66668 5122 66724 5134
rect 66668 5070 66670 5122
rect 66722 5070 66724 5122
rect 66668 4340 66724 5070
rect 66668 4274 66724 4284
rect 67564 5124 67620 5134
rect 64652 3574 64708 3612
rect 64876 3556 64932 3566
rect 64876 800 64932 3500
rect 65212 3556 65268 3566
rect 65212 3442 65268 3500
rect 65212 3390 65214 3442
rect 65266 3390 65268 3442
rect 65212 3378 65268 3390
rect 67564 800 67620 5068
rect 67900 5010 67956 5852
rect 67900 4958 67902 5010
rect 67954 4958 67956 5010
rect 67900 4946 67956 4958
rect 68236 5010 68292 6636
rect 68236 4958 68238 5010
rect 68290 4958 68292 5010
rect 68236 4946 68292 4958
rect 68460 5572 68516 5582
rect 67676 3892 67732 3902
rect 67676 3778 67732 3836
rect 67676 3726 67678 3778
rect 67730 3726 67732 3778
rect 67676 3714 67732 3726
rect 68460 3778 68516 5516
rect 68572 4340 68628 7980
rect 68684 7362 68740 7374
rect 68684 7310 68686 7362
rect 68738 7310 68740 7362
rect 68684 6132 68740 7310
rect 68684 5796 68740 6076
rect 69132 7362 69188 7374
rect 69132 7310 69134 7362
rect 69186 7310 69188 7362
rect 69132 6580 69188 7310
rect 69468 7362 69524 20132
rect 71708 12740 71764 22876
rect 71708 8428 71764 12684
rect 73724 11732 73780 33404
rect 76076 33458 76132 34636
rect 76188 34580 76244 34860
rect 76188 34514 76244 34524
rect 76300 34356 76356 34366
rect 76300 34262 76356 34300
rect 76076 33406 76078 33458
rect 76130 33406 76132 33458
rect 76076 33394 76132 33406
rect 76412 33460 76468 36318
rect 76860 36370 76916 36382
rect 76860 36318 76862 36370
rect 76914 36318 76916 36370
rect 76636 35474 76692 35486
rect 76636 35422 76638 35474
rect 76690 35422 76692 35474
rect 76524 33460 76580 33470
rect 76412 33458 76580 33460
rect 76412 33406 76526 33458
rect 76578 33406 76580 33458
rect 76412 33404 76580 33406
rect 76524 33394 76580 33404
rect 74852 32956 75116 32966
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 74852 32890 75116 32900
rect 74852 31388 75116 31398
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 74852 31322 75116 31332
rect 74852 29820 75116 29830
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 74852 29754 75116 29764
rect 74852 28252 75116 28262
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 74852 28186 75116 28196
rect 75516 26964 75572 26974
rect 74852 26684 75116 26694
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 74852 26618 75116 26628
rect 74852 25116 75116 25126
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 74852 25050 75116 25060
rect 74852 23548 75116 23558
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 74852 23482 75116 23492
rect 74852 21980 75116 21990
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 74852 21914 75116 21924
rect 74852 20412 75116 20422
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 74852 20346 75116 20356
rect 74852 18844 75116 18854
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 74852 18778 75116 18788
rect 74852 17276 75116 17286
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 74852 17210 75116 17220
rect 74852 15708 75116 15718
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 74852 15642 75116 15652
rect 74852 14140 75116 14150
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 74852 14074 75116 14084
rect 74852 12572 75116 12582
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 74852 12506 75116 12516
rect 73724 11666 73780 11676
rect 74852 11004 75116 11014
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 74852 10938 75116 10948
rect 74852 9436 75116 9446
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 74852 9370 75116 9380
rect 71708 8372 71876 8428
rect 69468 7310 69470 7362
rect 69522 7310 69524 7362
rect 69468 6916 69524 7310
rect 69916 7364 69972 7374
rect 69916 7362 70084 7364
rect 69916 7310 69918 7362
rect 69970 7310 70084 7362
rect 69916 7308 70084 7310
rect 69916 7298 69972 7308
rect 69468 6850 69524 6860
rect 69132 5908 69188 6524
rect 69468 6578 69524 6590
rect 69468 6526 69470 6578
rect 69522 6526 69524 6578
rect 69356 6468 69412 6478
rect 69356 6374 69412 6412
rect 69468 6468 69524 6526
rect 69916 6468 69972 6478
rect 69468 6466 69972 6468
rect 69468 6414 69918 6466
rect 69970 6414 69972 6466
rect 69468 6412 69972 6414
rect 69132 5842 69188 5852
rect 68684 4450 68740 5740
rect 69468 5348 69524 6412
rect 69916 6402 69972 6412
rect 68684 4398 68686 4450
rect 68738 4398 68740 4450
rect 68684 4386 68740 4398
rect 69356 5292 69524 5348
rect 69356 4900 69412 5292
rect 69468 5124 69524 5134
rect 69468 5030 69524 5068
rect 68572 4274 68628 4284
rect 69244 4340 69300 4350
rect 69244 4246 69300 4284
rect 68460 3726 68462 3778
rect 68514 3726 68516 3778
rect 68460 3714 68516 3726
rect 68572 3668 68628 3678
rect 68572 3574 68628 3612
rect 69356 3668 69412 4844
rect 69356 3602 69412 3612
rect 69580 3444 69636 3454
rect 70028 3444 70084 7308
rect 71260 6692 71316 6702
rect 70700 6690 71316 6692
rect 70700 6638 71262 6690
rect 71314 6638 71316 6690
rect 70700 6636 71316 6638
rect 70700 6468 70756 6636
rect 71260 6626 71316 6636
rect 70588 6466 70756 6468
rect 70588 6414 70702 6466
rect 70754 6414 70756 6466
rect 70588 6412 70756 6414
rect 70140 6130 70196 6142
rect 70140 6078 70142 6130
rect 70194 6078 70196 6130
rect 70140 6020 70196 6078
rect 70140 5954 70196 5964
rect 70476 5684 70532 5694
rect 70476 5122 70532 5628
rect 70476 5070 70478 5122
rect 70530 5070 70532 5122
rect 70476 5058 70532 5070
rect 69580 3442 70084 3444
rect 69580 3390 69582 3442
rect 69634 3390 70084 3442
rect 69580 3388 70084 3390
rect 68908 924 69300 980
rect 68908 800 68964 924
rect 4368 0 4480 800
rect 5712 0 5824 800
rect 7056 0 7168 800
rect 8400 0 8512 800
rect 9744 0 9856 800
rect 11088 0 11200 800
rect 12432 0 12544 800
rect 13776 0 13888 800
rect 15120 0 15232 800
rect 16464 0 16576 800
rect 17808 0 17920 800
rect 19152 0 19264 800
rect 20496 0 20608 800
rect 21840 0 21952 800
rect 23184 0 23296 800
rect 24528 0 24640 800
rect 25872 0 25984 800
rect 27216 0 27328 800
rect 28560 0 28672 800
rect 29904 0 30016 800
rect 31248 0 31360 800
rect 32592 0 32704 800
rect 33936 0 34048 800
rect 35280 0 35392 800
rect 36624 0 36736 800
rect 37968 0 38080 800
rect 39312 0 39424 800
rect 40656 0 40768 800
rect 42000 0 42112 800
rect 43344 0 43456 800
rect 44688 0 44800 800
rect 46032 0 46144 800
rect 47376 0 47488 800
rect 48720 0 48832 800
rect 50064 0 50176 800
rect 51408 0 51520 800
rect 52752 0 52864 800
rect 54096 0 54208 800
rect 55440 0 55552 800
rect 56784 0 56896 800
rect 58128 0 58240 800
rect 59472 0 59584 800
rect 60816 0 60928 800
rect 62160 0 62272 800
rect 63504 0 63616 800
rect 64848 0 64960 800
rect 66192 0 66304 800
rect 67536 0 67648 800
rect 68880 0 68992 800
rect 69244 756 69300 924
rect 69580 756 69636 3388
rect 70588 2548 70644 6412
rect 70700 6402 70756 6412
rect 71148 6020 71204 6030
rect 71148 5926 71204 5964
rect 70700 5908 70756 5918
rect 70700 5814 70756 5852
rect 71260 5796 71316 5806
rect 71708 5796 71764 5806
rect 71148 5794 71764 5796
rect 71148 5742 71262 5794
rect 71314 5742 71710 5794
rect 71762 5742 71764 5794
rect 71148 5740 71764 5742
rect 71148 4900 71204 5740
rect 71260 5730 71316 5740
rect 71708 5730 71764 5740
rect 71484 5012 71540 5022
rect 71484 4918 71540 4956
rect 71148 4806 71204 4844
rect 70588 2482 70644 2492
rect 71596 4226 71652 4238
rect 71596 4174 71598 4226
rect 71650 4174 71652 4226
rect 71596 800 71652 4174
rect 71708 3780 71764 3790
rect 71820 3780 71876 8372
rect 74852 7868 75116 7878
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 74852 7802 75116 7812
rect 74620 7364 74676 7374
rect 74060 7252 74116 7262
rect 72604 6580 72660 6590
rect 72156 6132 72212 6142
rect 72156 6038 72212 6076
rect 72604 5796 72660 6524
rect 73276 6580 73332 6590
rect 73276 6132 73332 6524
rect 73500 6132 73556 6142
rect 73276 6130 73556 6132
rect 73276 6078 73502 6130
rect 73554 6078 73556 6130
rect 73276 6076 73556 6078
rect 73500 6066 73556 6076
rect 74060 6130 74116 7196
rect 74060 6078 74062 6130
rect 74114 6078 74116 6130
rect 74060 6066 74116 6078
rect 72492 5794 72660 5796
rect 72492 5742 72606 5794
rect 72658 5742 72660 5794
rect 72492 5740 72660 5742
rect 72380 5348 72436 5358
rect 71932 5012 71988 5022
rect 71932 4918 71988 4956
rect 72380 4338 72436 5292
rect 72380 4286 72382 4338
rect 72434 4286 72436 4338
rect 72380 4274 72436 4286
rect 72492 5124 72548 5740
rect 72604 5730 72660 5740
rect 72940 6020 72996 6030
rect 72940 5348 72996 5964
rect 72940 5216 72996 5292
rect 72492 4340 72548 5068
rect 72604 4900 72660 4910
rect 73724 4900 73780 4910
rect 72604 4898 72772 4900
rect 72604 4846 72606 4898
rect 72658 4846 72772 4898
rect 72604 4844 72772 4846
rect 72604 4834 72660 4844
rect 72492 4274 72548 4284
rect 71708 3778 71876 3780
rect 71708 3726 71710 3778
rect 71762 3726 71876 3778
rect 71708 3724 71876 3726
rect 71708 3714 71764 3724
rect 72604 3556 72660 3566
rect 72604 3462 72660 3500
rect 72716 3444 72772 4844
rect 73724 4806 73780 4844
rect 74620 4338 74676 7308
rect 75068 7364 75124 7374
rect 75516 7364 75572 26908
rect 76636 26964 76692 35422
rect 76860 34580 76916 36318
rect 77308 35700 77364 35710
rect 77308 35606 77364 35644
rect 76860 34514 76916 34524
rect 77420 34914 77476 34926
rect 77420 34862 77422 34914
rect 77474 34862 77476 34914
rect 76860 34356 76916 34366
rect 76860 34242 76916 34300
rect 76860 34190 76862 34242
rect 76914 34190 76916 34242
rect 76860 34178 76916 34190
rect 77196 34242 77252 34254
rect 77196 34190 77198 34242
rect 77250 34190 77252 34242
rect 77196 31332 77252 34190
rect 77420 34020 77476 34862
rect 77644 34692 77700 34702
rect 77644 34690 77812 34692
rect 77644 34638 77646 34690
rect 77698 34638 77812 34690
rect 77644 34636 77812 34638
rect 77644 34626 77700 34636
rect 77644 34020 77700 34030
rect 77420 34018 77700 34020
rect 77420 33966 77646 34018
rect 77698 33966 77700 34018
rect 77420 33964 77700 33966
rect 77644 33124 77700 33964
rect 77756 33460 77812 34636
rect 77756 33394 77812 33404
rect 77980 33458 78036 36428
rect 78204 36418 78260 36428
rect 78092 35812 78148 35822
rect 78092 35586 78148 35756
rect 78092 35534 78094 35586
rect 78146 35534 78148 35586
rect 78092 35522 78148 35534
rect 78204 34804 78260 34814
rect 78204 34710 78260 34748
rect 78204 34018 78260 34030
rect 78204 33966 78206 34018
rect 78258 33966 78260 34018
rect 78204 33906 78260 33966
rect 78204 33854 78206 33906
rect 78258 33854 78260 33906
rect 78204 33842 78260 33854
rect 77980 33406 77982 33458
rect 78034 33406 78036 33458
rect 77644 33058 77700 33068
rect 77196 31266 77252 31276
rect 76636 26898 76692 26908
rect 77980 24724 78036 33406
rect 77980 24658 78036 24668
rect 75068 7270 75124 7308
rect 75404 7362 75572 7364
rect 75404 7310 75518 7362
rect 75570 7310 75572 7362
rect 75404 7308 75572 7310
rect 75180 7252 75236 7262
rect 74852 6300 75116 6310
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 74852 6234 75116 6244
rect 74732 6020 74788 6030
rect 74732 5926 74788 5964
rect 75180 6018 75236 7196
rect 75180 5966 75182 6018
rect 75234 5966 75236 6018
rect 75180 5954 75236 5966
rect 75404 5906 75460 7308
rect 75516 7298 75572 7308
rect 75852 12852 75908 12862
rect 75740 6580 75796 6590
rect 75740 6130 75796 6524
rect 75740 6078 75742 6130
rect 75794 6078 75796 6130
rect 75740 6066 75796 6078
rect 75404 5854 75406 5906
rect 75458 5854 75460 5906
rect 75404 5842 75460 5854
rect 75628 5124 75684 5134
rect 74852 4732 75116 4742
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 74852 4666 75116 4676
rect 74620 4286 74622 4338
rect 74674 4286 74676 4338
rect 74620 4274 74676 4286
rect 75628 4338 75684 5068
rect 75628 4286 75630 4338
rect 75682 4286 75684 4338
rect 75628 4274 75684 4286
rect 73836 4226 73892 4238
rect 73836 4174 73838 4226
rect 73890 4174 73892 4226
rect 73164 3444 73220 3454
rect 72716 3442 73220 3444
rect 72716 3390 73166 3442
rect 73218 3390 73220 3442
rect 72716 3388 73220 3390
rect 72940 800 72996 3388
rect 73164 3378 73220 3388
rect 73836 3444 73892 4174
rect 75628 3780 75684 3790
rect 75852 3780 75908 12796
rect 76972 12852 77028 12862
rect 76972 11844 77028 12796
rect 76972 11778 77028 11788
rect 78316 7698 78372 36652
rect 78428 35588 78484 36764
rect 78428 35522 78484 35532
rect 78540 34804 78596 34814
rect 78540 34710 78596 34748
rect 78652 34354 78708 37996
rect 78652 34302 78654 34354
rect 78706 34302 78708 34354
rect 78652 34290 78708 34302
rect 78764 35476 78820 38668
rect 78988 37044 79044 39200
rect 79884 39060 79940 39200
rect 80220 39060 80276 39228
rect 79884 39004 80276 39060
rect 78988 36988 79156 37044
rect 78988 36820 79044 36830
rect 78988 36594 79044 36764
rect 78988 36542 78990 36594
rect 79042 36542 79044 36594
rect 78988 36530 79044 36542
rect 79100 36372 79156 36988
rect 80220 36596 80276 36606
rect 79100 36306 79156 36316
rect 79660 36594 80276 36596
rect 79660 36542 80222 36594
rect 80274 36542 80276 36594
rect 79660 36540 80276 36542
rect 78764 33906 78820 35420
rect 79100 35698 79156 35710
rect 79100 35646 79102 35698
rect 79154 35646 79156 35698
rect 78988 34690 79044 34702
rect 78988 34638 78990 34690
rect 79042 34638 79044 34690
rect 78988 34580 79044 34638
rect 78988 34514 79044 34524
rect 78764 33854 78766 33906
rect 78818 33854 78820 33906
rect 78764 33842 78820 33854
rect 79100 34018 79156 35646
rect 79436 34804 79492 34814
rect 79436 34710 79492 34748
rect 79100 33966 79102 34018
rect 79154 33966 79156 34018
rect 79100 29652 79156 33966
rect 79100 29586 79156 29596
rect 79660 27636 79716 36540
rect 80220 36530 80276 36540
rect 79772 35588 79828 35598
rect 79772 35494 79828 35532
rect 80556 35252 80612 39228
rect 80752 39200 80864 40000
rect 81648 39200 81760 40000
rect 82544 39200 82656 40000
rect 83440 39200 83552 40000
rect 84336 39200 84448 40000
rect 85232 39200 85344 40000
rect 86128 39200 86240 40000
rect 87024 39200 87136 40000
rect 87920 39200 88032 40000
rect 88816 39200 88928 40000
rect 89712 39200 89824 40000
rect 90608 39200 90720 40000
rect 91504 39200 91616 40000
rect 92400 39200 92512 40000
rect 93296 39200 93408 40000
rect 94192 39200 94304 40000
rect 95088 39200 95200 40000
rect 95984 39200 96096 40000
rect 96880 39200 96992 40000
rect 97776 39200 97888 40000
rect 98672 39200 98784 40000
rect 99568 39200 99680 40000
rect 100464 39200 100576 40000
rect 101360 39200 101472 40000
rect 102256 39200 102368 40000
rect 103152 39200 103264 40000
rect 104048 39200 104160 40000
rect 104944 39200 105056 40000
rect 105840 39200 105952 40000
rect 106736 39200 106848 40000
rect 107632 39200 107744 40000
rect 108528 39200 108640 40000
rect 109424 39200 109536 40000
rect 110320 39200 110432 40000
rect 111216 39200 111328 40000
rect 112112 39200 112224 40000
rect 113008 39200 113120 40000
rect 113904 39200 114016 40000
rect 114800 39200 114912 40000
rect 115696 39200 115808 40000
rect 116592 39200 116704 40000
rect 117488 39200 117600 40000
rect 118384 39200 118496 40000
rect 119280 39200 119392 40000
rect 120176 39200 120288 40000
rect 121072 39200 121184 40000
rect 121968 39200 122080 40000
rect 122864 39200 122976 40000
rect 123760 39200 123872 40000
rect 124656 39200 124768 40000
rect 125552 39200 125664 40000
rect 126448 39200 126560 40000
rect 127344 39200 127456 40000
rect 128240 39200 128352 40000
rect 129136 39200 129248 40000
rect 130032 39200 130144 40000
rect 130928 39200 131040 40000
rect 131824 39200 131936 40000
rect 132720 39200 132832 40000
rect 133616 39200 133728 40000
rect 134512 39200 134624 40000
rect 135408 39200 135520 40000
rect 136304 39200 136416 40000
rect 137200 39200 137312 40000
rect 138096 39200 138208 40000
rect 138992 39200 139104 40000
rect 139888 39200 140000 40000
rect 140784 39200 140896 40000
rect 141680 39200 141792 40000
rect 142044 39228 142436 39284
rect 80780 35700 80836 39200
rect 81564 37268 81620 37278
rect 81228 36372 81284 36382
rect 81228 36278 81284 36316
rect 81564 35812 81620 37212
rect 81676 36036 81732 39200
rect 82572 37378 82628 39200
rect 82572 37326 82574 37378
rect 82626 37326 82628 37378
rect 82572 37314 82628 37326
rect 82796 38948 82852 38958
rect 82572 37156 82628 37166
rect 82236 36370 82292 36382
rect 82236 36318 82238 36370
rect 82290 36318 82292 36370
rect 82236 36260 82292 36318
rect 82572 36370 82628 37100
rect 82572 36318 82574 36370
rect 82626 36318 82628 36370
rect 82572 36306 82628 36318
rect 81676 35980 81844 36036
rect 81676 35812 81732 35822
rect 81564 35810 81732 35812
rect 81564 35758 81678 35810
rect 81730 35758 81732 35810
rect 81564 35756 81732 35758
rect 81676 35746 81732 35756
rect 80780 35644 80948 35700
rect 80556 35196 80836 35252
rect 80780 35026 80836 35196
rect 80892 35140 80948 35644
rect 80892 35074 80948 35084
rect 81340 35698 81396 35710
rect 81340 35646 81342 35698
rect 81394 35646 81396 35698
rect 80780 34974 80782 35026
rect 80834 34974 80836 35026
rect 80780 34962 80836 34974
rect 80108 34916 80164 34926
rect 79772 34914 80164 34916
rect 79772 34862 80110 34914
rect 80162 34862 80164 34914
rect 79772 34860 80164 34862
rect 79772 34018 79828 34860
rect 80108 34850 80164 34860
rect 79772 33966 79774 34018
rect 79826 33966 79828 34018
rect 79772 27860 79828 33966
rect 80444 34804 80500 34814
rect 80444 33908 80500 34748
rect 80444 33842 80500 33852
rect 80556 34018 80612 34030
rect 80556 33966 80558 34018
rect 80610 33966 80612 34018
rect 80556 33236 80612 33966
rect 80556 33170 80612 33180
rect 81340 33236 81396 35646
rect 81788 34356 81844 35980
rect 82124 35588 82180 35598
rect 81788 34290 81844 34300
rect 82012 35586 82180 35588
rect 82012 35534 82126 35586
rect 82178 35534 82180 35586
rect 82012 35532 82180 35534
rect 82012 34914 82068 35532
rect 82124 35522 82180 35532
rect 82012 34862 82014 34914
rect 82066 34862 82068 34914
rect 81900 34130 81956 34142
rect 81900 34078 81902 34130
rect 81954 34078 81956 34130
rect 81340 33170 81396 33180
rect 81452 34020 81508 34030
rect 81900 34020 81956 34078
rect 81452 34018 81956 34020
rect 81452 33966 81454 34018
rect 81506 33966 81956 34018
rect 81452 33964 81956 33966
rect 81452 29988 81508 33964
rect 82012 31220 82068 34862
rect 82236 32676 82292 36204
rect 82796 35586 82852 38892
rect 83020 36372 83076 36382
rect 83020 36278 83076 36316
rect 83468 35812 83524 39200
rect 84028 38164 84084 38174
rect 83468 35746 83524 35756
rect 83804 37378 83860 37390
rect 83804 37326 83806 37378
rect 83858 37326 83860 37378
rect 83804 35810 83860 37326
rect 83804 35758 83806 35810
rect 83858 35758 83860 35810
rect 82796 35534 82798 35586
rect 82850 35534 82852 35586
rect 82796 35522 82852 35534
rect 82572 35140 82628 35150
rect 82572 35026 82628 35084
rect 82572 34974 82574 35026
rect 82626 34974 82628 35026
rect 82572 34962 82628 34974
rect 82572 34804 82628 34814
rect 82572 33458 82628 34748
rect 83804 34804 83860 35758
rect 83804 34738 83860 34748
rect 84028 34802 84084 38108
rect 84028 34750 84030 34802
rect 84082 34750 84084 34802
rect 84028 34738 84084 34750
rect 84140 36370 84196 36382
rect 84140 36318 84142 36370
rect 84194 36318 84196 36370
rect 82684 34356 82740 34366
rect 82684 34018 82740 34300
rect 83804 34132 83860 34142
rect 83804 34038 83860 34076
rect 84140 34132 84196 36318
rect 84364 35140 84420 39200
rect 84476 36258 84532 36270
rect 84476 36206 84478 36258
rect 84530 36206 84532 36258
rect 84476 36148 84532 36206
rect 84924 36260 84980 36270
rect 84924 36166 84980 36204
rect 84476 36082 84532 36092
rect 84924 35812 84980 35822
rect 84924 35718 84980 35756
rect 85260 35812 85316 39200
rect 85820 38836 85876 38846
rect 85820 36594 85876 38780
rect 85820 36542 85822 36594
rect 85874 36542 85876 36594
rect 85820 36530 85876 36542
rect 86156 36484 86212 39200
rect 86156 36418 86212 36428
rect 86828 36484 86884 36494
rect 86828 36370 86884 36428
rect 86828 36318 86830 36370
rect 86882 36318 86884 36370
rect 86828 36306 86884 36318
rect 85260 35746 85316 35756
rect 86716 35812 86772 35822
rect 86716 35718 86772 35756
rect 84364 35074 84420 35084
rect 85820 35698 85876 35710
rect 85820 35646 85822 35698
rect 85874 35646 85876 35698
rect 85260 34916 85316 34926
rect 85148 34914 85316 34916
rect 85148 34862 85262 34914
rect 85314 34862 85316 34914
rect 85148 34860 85316 34862
rect 84140 34066 84196 34076
rect 84364 34802 84420 34814
rect 84364 34750 84366 34802
rect 84418 34750 84420 34802
rect 82684 33966 82686 34018
rect 82738 33966 82740 34018
rect 82684 33954 82740 33966
rect 84364 34020 84420 34750
rect 84588 34020 84644 34030
rect 84364 34018 84644 34020
rect 84364 33966 84590 34018
rect 84642 33966 84644 34018
rect 84364 33964 84644 33966
rect 82572 33406 82574 33458
rect 82626 33406 82628 33458
rect 82572 33394 82628 33406
rect 84588 33012 84644 33964
rect 84588 32946 84644 32956
rect 85148 34018 85204 34860
rect 85260 34850 85316 34860
rect 85820 34468 85876 35646
rect 85932 35140 85988 35150
rect 85932 35026 85988 35084
rect 87052 35140 87108 39200
rect 87612 35700 87668 35710
rect 87052 35074 87108 35084
rect 87500 35698 87668 35700
rect 87500 35646 87614 35698
rect 87666 35646 87668 35698
rect 87500 35644 87668 35646
rect 85932 34974 85934 35026
rect 85986 34974 85988 35026
rect 85932 34962 85988 34974
rect 87276 34916 87332 34926
rect 85148 33966 85150 34018
rect 85202 33966 85204 34018
rect 82236 32610 82292 32620
rect 82012 31154 82068 31164
rect 81452 29922 81508 29932
rect 85148 27972 85204 33966
rect 85148 27906 85204 27916
rect 85484 34412 85876 34468
rect 87052 34914 87332 34916
rect 87052 34862 87278 34914
rect 87330 34862 87332 34914
rect 87052 34860 87332 34862
rect 85484 34354 85540 34412
rect 85484 34302 85486 34354
rect 85538 34302 85540 34354
rect 79772 27794 79828 27804
rect 79660 27570 79716 27580
rect 85484 26180 85540 34302
rect 87052 34018 87108 34860
rect 87276 34850 87332 34860
rect 87052 33966 87054 34018
rect 87106 33966 87108 34018
rect 87052 26516 87108 33966
rect 87500 27300 87556 35644
rect 87612 35588 87668 35644
rect 87836 35588 87892 35598
rect 87612 35586 87892 35588
rect 87612 35534 87838 35586
rect 87890 35534 87892 35586
rect 87612 35532 87892 35534
rect 87836 35522 87892 35532
rect 87948 35364 88004 39200
rect 88396 36482 88452 36494
rect 88396 36430 88398 36482
rect 88450 36430 88452 36482
rect 88284 35698 88340 35710
rect 88284 35646 88286 35698
rect 88338 35646 88340 35698
rect 88172 35588 88228 35598
rect 88284 35588 88340 35646
rect 88172 35586 88340 35588
rect 88172 35534 88174 35586
rect 88226 35534 88340 35586
rect 88172 35532 88340 35534
rect 88172 35522 88228 35532
rect 87948 35308 88116 35364
rect 87948 35140 88004 35150
rect 87948 35026 88004 35084
rect 87948 34974 87950 35026
rect 88002 34974 88004 35026
rect 87948 34962 88004 34974
rect 87612 34356 87668 34366
rect 87612 33684 87668 34300
rect 87612 33618 87668 33628
rect 88060 33460 88116 35308
rect 88396 34356 88452 36430
rect 88620 36258 88676 36270
rect 88620 36206 88622 36258
rect 88674 36206 88676 36258
rect 88620 34804 88676 36206
rect 88620 34738 88676 34748
rect 88396 34290 88452 34300
rect 88508 34692 88564 34702
rect 88172 34020 88228 34030
rect 88172 33926 88228 33964
rect 88060 33394 88116 33404
rect 88172 33346 88228 33358
rect 88172 33294 88174 33346
rect 88226 33294 88228 33346
rect 87724 33124 87780 33134
rect 88172 33124 88228 33294
rect 87724 33122 88228 33124
rect 87724 33070 87726 33122
rect 87778 33070 88228 33122
rect 87724 33068 88228 33070
rect 87724 30884 87780 33068
rect 87724 30818 87780 30828
rect 87500 27234 87556 27244
rect 87052 26450 87108 26460
rect 85484 26114 85540 26124
rect 80668 24388 80724 24398
rect 79772 23044 79828 23054
rect 79772 11844 79828 22988
rect 80668 20188 80724 24332
rect 86492 22932 86548 22942
rect 84924 21364 84980 21374
rect 83132 21028 83188 21038
rect 80668 20132 80836 20188
rect 79772 11778 79828 11788
rect 78316 7646 78318 7698
rect 78370 7646 78372 7698
rect 76300 7586 76356 7598
rect 76300 7534 76302 7586
rect 76354 7534 76356 7586
rect 76076 6468 76132 6478
rect 76076 5122 76132 6412
rect 76300 5684 76356 7534
rect 76748 7586 76804 7598
rect 76748 7534 76750 7586
rect 76802 7534 76804 7586
rect 76748 7252 76804 7534
rect 76972 7476 77028 7486
rect 76972 7382 77028 7420
rect 78316 7476 78372 7646
rect 78316 7410 78372 7420
rect 78428 11732 78484 11742
rect 77868 7362 77924 7374
rect 77868 7310 77870 7362
rect 77922 7310 77924 7362
rect 76748 7186 76804 7196
rect 77308 7252 77364 7262
rect 77644 7252 77700 7262
rect 77308 7250 77700 7252
rect 77308 7198 77310 7250
rect 77362 7198 77646 7250
rect 77698 7198 77700 7250
rect 77308 7196 77700 7198
rect 77308 7186 77364 7196
rect 77644 7186 77700 7196
rect 77868 7252 77924 7310
rect 77868 7186 77924 7196
rect 78204 7250 78260 7262
rect 78204 7198 78206 7250
rect 78258 7198 78260 7250
rect 78204 6690 78260 7198
rect 78204 6638 78206 6690
rect 78258 6638 78260 6690
rect 78204 6626 78260 6638
rect 77644 6580 77700 6590
rect 77644 6486 77700 6524
rect 77308 6468 77364 6478
rect 77308 6374 77364 6412
rect 76300 5590 76356 5628
rect 77084 6018 77140 6030
rect 77084 5966 77086 6018
rect 77138 5966 77140 6018
rect 76076 5070 76078 5122
rect 76130 5070 76132 5122
rect 76076 5058 76132 5070
rect 76300 5124 76356 5134
rect 75628 3778 75908 3780
rect 75628 3726 75630 3778
rect 75682 3726 75908 3778
rect 75628 3724 75908 3726
rect 75628 3714 75684 3724
rect 76300 3666 76356 5068
rect 76300 3614 76302 3666
rect 76354 3614 76356 3666
rect 76300 3602 76356 3614
rect 76636 5124 76692 5134
rect 76636 3668 76692 5068
rect 77084 3780 77140 5966
rect 77308 5236 77364 5246
rect 77308 5122 77364 5180
rect 77308 5070 77310 5122
rect 77362 5070 77364 5122
rect 77308 5058 77364 5070
rect 77084 3714 77140 3724
rect 76748 3668 76804 3678
rect 76636 3666 76804 3668
rect 76636 3614 76750 3666
rect 76802 3614 76804 3666
rect 76636 3612 76804 3614
rect 76748 3602 76804 3612
rect 78428 3666 78484 11676
rect 80780 8372 80836 20132
rect 79996 6580 80052 6590
rect 79660 6578 80052 6580
rect 79660 6526 79998 6578
rect 80050 6526 80052 6578
rect 79660 6524 80052 6526
rect 78540 6468 78596 6478
rect 78540 6374 78596 6412
rect 79324 6468 79380 6478
rect 79324 5906 79380 6412
rect 79324 5854 79326 5906
rect 79378 5854 79380 5906
rect 79324 5842 79380 5854
rect 79212 3780 79268 3790
rect 79212 3686 79268 3724
rect 78428 3614 78430 3666
rect 78482 3614 78484 3666
rect 78428 3602 78484 3614
rect 79324 3668 79380 3678
rect 79324 3574 79380 3612
rect 76972 3556 77028 3566
rect 73836 3378 73892 3388
rect 75628 3444 75684 3454
rect 74852 3164 75116 3174
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 74852 3098 75116 3108
rect 75628 800 75684 3388
rect 76972 800 77028 3500
rect 77308 3556 77364 3566
rect 77308 3442 77364 3500
rect 77308 3390 77310 3442
rect 77362 3390 77364 3442
rect 77308 3378 77364 3390
rect 79660 800 79716 6524
rect 79996 6514 80052 6524
rect 79996 5906 80052 5918
rect 79996 5854 79998 5906
rect 80050 5854 80052 5906
rect 79996 5796 80052 5854
rect 80444 5796 80500 5806
rect 79996 5794 80500 5796
rect 79996 5742 80446 5794
rect 80498 5742 80500 5794
rect 79996 5740 80500 5742
rect 80444 5124 80500 5740
rect 80332 5068 80444 5124
rect 80220 4900 80276 4910
rect 80220 3778 80276 4844
rect 80332 4450 80388 5068
rect 80444 5058 80500 5068
rect 80332 4398 80334 4450
rect 80386 4398 80388 4450
rect 80332 4386 80388 4398
rect 80444 4676 80500 4686
rect 80220 3726 80222 3778
rect 80274 3726 80276 3778
rect 80220 3714 80276 3726
rect 80332 3668 80388 3678
rect 80444 3668 80500 4620
rect 80780 3778 80836 8316
rect 83132 8372 83188 20972
rect 84924 15988 84980 21308
rect 84924 15922 84980 15932
rect 83132 8306 83188 8316
rect 84700 14308 84756 14318
rect 81788 7588 81844 7598
rect 81116 6690 81172 6702
rect 81116 6638 81118 6690
rect 81170 6638 81172 6690
rect 81116 6580 81172 6638
rect 81116 6514 81172 6524
rect 81564 6580 81620 6590
rect 81564 6486 81620 6524
rect 81228 4676 81284 4686
rect 81228 4562 81284 4620
rect 81228 4510 81230 4562
rect 81282 4510 81284 4562
rect 81228 4498 81284 4510
rect 81676 4676 81732 4686
rect 81676 4562 81732 4620
rect 81676 4510 81678 4562
rect 81730 4510 81732 4562
rect 81676 4498 81732 4510
rect 81788 3892 81844 7532
rect 84476 5124 84532 5134
rect 84476 5030 84532 5068
rect 82236 5012 82292 5022
rect 82236 4918 82292 4956
rect 84028 4228 84084 4238
rect 81788 3826 81844 3836
rect 83692 4226 84084 4228
rect 83692 4174 84030 4226
rect 84082 4174 84084 4226
rect 83692 4172 84084 4174
rect 80780 3726 80782 3778
rect 80834 3726 80836 3778
rect 80780 3714 80836 3726
rect 80388 3612 80500 3668
rect 80332 3536 80388 3612
rect 81004 3444 81060 3454
rect 81004 800 81060 3388
rect 82908 3444 82964 3454
rect 82908 3350 82964 3388
rect 83692 800 83748 4172
rect 84028 4162 84084 4172
rect 84700 3778 84756 14252
rect 86492 14308 86548 22876
rect 86492 14242 86548 14252
rect 88508 7476 88564 34636
rect 88620 34244 88676 34254
rect 88620 34150 88676 34188
rect 88844 33572 88900 39200
rect 89740 36820 89796 39200
rect 89740 36764 89908 36820
rect 89740 36594 89796 36606
rect 89740 36542 89742 36594
rect 89794 36542 89796 36594
rect 89068 36484 89124 36494
rect 89068 36390 89124 36428
rect 89180 36372 89236 36382
rect 88956 35252 89012 35262
rect 88956 35026 89012 35196
rect 88956 34974 88958 35026
rect 89010 34974 89012 35026
rect 88956 34962 89012 34974
rect 88844 33506 88900 33516
rect 88956 34580 89012 34590
rect 88956 28084 89012 34524
rect 89068 33460 89124 33470
rect 89068 33366 89124 33404
rect 89180 32788 89236 36316
rect 89516 36372 89572 36382
rect 89516 35810 89572 36316
rect 89516 35758 89518 35810
rect 89570 35758 89572 35810
rect 89516 35746 89572 35758
rect 89628 34692 89684 34702
rect 89628 34598 89684 34636
rect 89740 34356 89796 36542
rect 89852 36372 89908 36764
rect 89852 36306 89908 36316
rect 90188 36260 90244 36270
rect 89964 35810 90020 35822
rect 89964 35758 89966 35810
rect 90018 35758 90020 35810
rect 89964 35700 90020 35758
rect 89964 35634 90020 35644
rect 90188 35698 90244 36204
rect 90188 35646 90190 35698
rect 90242 35646 90244 35698
rect 90188 35634 90244 35646
rect 90412 35700 90468 35710
rect 90300 35252 90356 35262
rect 89964 34916 90020 34926
rect 89964 34914 90132 34916
rect 89964 34862 89966 34914
rect 90018 34862 90132 34914
rect 89964 34860 90132 34862
rect 89964 34850 90020 34860
rect 89516 34300 89796 34356
rect 89292 34244 89348 34254
rect 89292 34242 89460 34244
rect 89292 34190 89294 34242
rect 89346 34190 89460 34242
rect 89292 34188 89460 34190
rect 89292 34178 89348 34188
rect 89292 32788 89348 32798
rect 89180 32786 89348 32788
rect 89180 32734 89294 32786
rect 89346 32734 89348 32786
rect 89180 32732 89348 32734
rect 89292 32722 89348 32732
rect 88956 28018 89012 28028
rect 89404 23156 89460 34188
rect 89516 24948 89572 34300
rect 89516 24882 89572 24892
rect 89628 34130 89684 34142
rect 89628 34078 89630 34130
rect 89682 34078 89684 34130
rect 89628 34020 89684 34078
rect 89628 24500 89684 33964
rect 89964 33346 90020 33358
rect 89964 33294 89966 33346
rect 90018 33294 90020 33346
rect 89740 32452 89796 32462
rect 89964 32452 90020 33294
rect 90076 32676 90132 34860
rect 90300 34356 90356 35196
rect 90412 34914 90468 35644
rect 90636 35588 90692 39200
rect 91420 37044 91476 37054
rect 90748 36372 90804 36382
rect 90804 36316 90916 36372
rect 90748 36278 90804 36316
rect 90636 35532 90804 35588
rect 90524 35476 90580 35486
rect 90524 35474 90692 35476
rect 90524 35422 90526 35474
rect 90578 35422 90692 35474
rect 90524 35420 90692 35422
rect 90524 35410 90580 35420
rect 90412 34862 90414 34914
rect 90466 34862 90468 34914
rect 90412 34850 90468 34862
rect 90524 34802 90580 34814
rect 90524 34750 90526 34802
rect 90578 34750 90580 34802
rect 90524 34580 90580 34750
rect 90524 34514 90580 34524
rect 90300 34130 90356 34300
rect 90412 34244 90468 34254
rect 90412 34150 90468 34188
rect 90300 34078 90302 34130
rect 90354 34078 90356 34130
rect 90300 34066 90356 34078
rect 90076 32610 90132 32620
rect 89740 32450 90020 32452
rect 89740 32398 89742 32450
rect 89794 32398 90020 32450
rect 89740 32396 90020 32398
rect 89740 27188 89796 32396
rect 89740 27122 89796 27132
rect 90636 26908 90692 35420
rect 90748 35252 90804 35532
rect 90748 35186 90804 35196
rect 90860 34132 90916 36316
rect 91420 35810 91476 36988
rect 91420 35758 91422 35810
rect 91474 35758 91476 35810
rect 91420 35746 91476 35758
rect 90860 34066 90916 34076
rect 91196 35700 91252 35710
rect 91084 34020 91140 34030
rect 91084 33926 91140 33964
rect 90748 33572 90804 33582
rect 90748 33458 90804 33516
rect 90748 33406 90750 33458
rect 90802 33406 90804 33458
rect 90748 33394 90804 33406
rect 90748 32788 90804 32798
rect 91196 32788 91252 35644
rect 91308 35698 91364 35710
rect 91308 35646 91310 35698
rect 91362 35646 91364 35698
rect 91308 35140 91364 35646
rect 91308 35074 91364 35084
rect 91532 35140 91588 39200
rect 91980 36370 92036 36382
rect 91980 36318 91982 36370
rect 92034 36318 92036 36370
rect 91980 36148 92036 36318
rect 91532 35074 91588 35084
rect 91756 36092 92036 36148
rect 92316 36258 92372 36270
rect 92316 36206 92318 36258
rect 92370 36206 92372 36258
rect 91308 34690 91364 34702
rect 91308 34638 91310 34690
rect 91362 34638 91364 34690
rect 91308 34580 91364 34638
rect 91308 34514 91364 34524
rect 90748 32786 91252 32788
rect 90748 32734 90750 32786
rect 90802 32734 91198 32786
rect 91250 32734 91252 32786
rect 90748 32732 91252 32734
rect 90748 32722 90804 32732
rect 91196 32722 91252 32732
rect 91420 33906 91476 33918
rect 91420 33854 91422 33906
rect 91474 33854 91476 33906
rect 89628 24434 89684 24444
rect 90524 26852 90692 26908
rect 89404 23090 89460 23100
rect 87500 7474 88564 7476
rect 87500 7422 88510 7474
rect 88562 7422 88564 7474
rect 87500 7420 88564 7422
rect 87500 7252 87556 7420
rect 88508 7410 88564 7420
rect 88620 15988 88676 15998
rect 87388 7196 87556 7252
rect 87612 7252 87668 7262
rect 87388 6914 87444 7196
rect 87388 6862 87390 6914
rect 87442 6862 87444 6914
rect 87388 6850 87444 6862
rect 87612 6580 87668 7196
rect 88172 6580 88228 6590
rect 87612 6578 88004 6580
rect 87612 6526 87614 6578
rect 87666 6526 88004 6578
rect 87612 6524 88004 6526
rect 87612 6514 87668 6524
rect 85596 6468 85652 6478
rect 87052 6468 87108 6478
rect 85484 5124 85540 5134
rect 85484 5030 85540 5068
rect 85596 4564 85652 6412
rect 86492 6466 87108 6468
rect 86492 6414 87054 6466
rect 87106 6414 87108 6466
rect 86492 6412 87108 6414
rect 86156 6020 86212 6030
rect 85932 6018 86212 6020
rect 85932 5966 86158 6018
rect 86210 5966 86212 6018
rect 85932 5964 86212 5966
rect 85932 5122 85988 5964
rect 86156 5954 86212 5964
rect 86492 6018 86548 6412
rect 87052 6402 87108 6412
rect 87388 6132 87444 6142
rect 87388 6038 87444 6076
rect 86492 5966 86494 6018
rect 86546 5966 86548 6018
rect 86492 5954 86548 5966
rect 87948 5906 88004 6524
rect 88172 6486 88228 6524
rect 88508 6132 88564 6142
rect 88508 6038 88564 6076
rect 87948 5854 87950 5906
rect 88002 5854 88004 5906
rect 87948 5842 88004 5854
rect 85932 5070 85934 5122
rect 85986 5070 85988 5122
rect 85932 5058 85988 5070
rect 88396 5236 88452 5246
rect 85148 4562 85652 4564
rect 85148 4510 85598 4562
rect 85650 4510 85652 4562
rect 85148 4508 85652 4510
rect 85148 4338 85204 4508
rect 85596 4498 85652 4508
rect 86268 5012 86324 5022
rect 86268 4562 86324 4956
rect 88396 4898 88452 5180
rect 88396 4846 88398 4898
rect 88450 4846 88452 4898
rect 88396 4834 88452 4846
rect 86268 4510 86270 4562
rect 86322 4510 86324 4562
rect 85148 4286 85150 4338
rect 85202 4286 85204 4338
rect 85148 4274 85204 4286
rect 86268 4340 86324 4510
rect 86828 4452 86884 4462
rect 86828 4358 86884 4396
rect 88508 4452 88564 4462
rect 86268 4274 86324 4284
rect 88508 4338 88564 4396
rect 88508 4286 88510 4338
rect 88562 4286 88564 4338
rect 88508 4274 88564 4286
rect 84700 3726 84702 3778
rect 84754 3726 84756 3778
rect 84700 3714 84756 3726
rect 87724 4226 87780 4238
rect 87724 4174 87726 4226
rect 87778 4174 87780 4226
rect 84028 3444 84084 3454
rect 84028 3350 84084 3388
rect 85036 3444 85092 3454
rect 85036 800 85092 3388
rect 86828 3444 86884 3454
rect 86828 3350 86884 3388
rect 87724 800 87780 4174
rect 88620 3778 88676 15932
rect 90524 8428 90580 26852
rect 91420 11172 91476 33854
rect 91644 32676 91700 32686
rect 91644 32582 91700 32620
rect 91756 32452 91812 36092
rect 92092 35588 92148 35598
rect 92092 35494 92148 35532
rect 92092 34804 92148 34814
rect 91980 34802 92148 34804
rect 91980 34750 92094 34802
rect 92146 34750 92148 34802
rect 91980 34748 92148 34750
rect 91868 34020 91924 34030
rect 91868 33458 91924 33964
rect 91868 33406 91870 33458
rect 91922 33406 91924 33458
rect 91868 33394 91924 33406
rect 91980 32564 92036 34748
rect 92092 34738 92148 34748
rect 92316 34244 92372 36206
rect 92428 35924 92484 39200
rect 92764 37044 92820 37054
rect 92764 36594 92820 36988
rect 93324 37044 93380 39200
rect 93324 36978 93380 36988
rect 93262 36876 93526 36886
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93262 36810 93526 36820
rect 93660 36820 93716 36830
rect 93548 36596 93604 36606
rect 92764 36542 92766 36594
rect 92818 36542 92820 36594
rect 92764 36530 92820 36542
rect 93212 36594 93604 36596
rect 93212 36542 93550 36594
rect 93602 36542 93604 36594
rect 93212 36540 93604 36542
rect 93212 36148 93268 36540
rect 93548 36530 93604 36540
rect 92428 35858 92484 35868
rect 92876 36092 93268 36148
rect 93660 36260 93716 36764
rect 92428 35476 92484 35486
rect 92428 35474 92708 35476
rect 92428 35422 92430 35474
rect 92482 35422 92708 35474
rect 92428 35420 92708 35422
rect 92428 35410 92484 35420
rect 92428 34690 92484 34702
rect 92428 34638 92430 34690
rect 92482 34638 92484 34690
rect 92428 34580 92484 34638
rect 92428 34514 92484 34524
rect 92316 34178 92372 34188
rect 91980 32470 92036 32508
rect 92204 34130 92260 34142
rect 92204 34078 92206 34130
rect 92258 34078 92260 34130
rect 92204 33122 92260 34078
rect 92204 33070 92206 33122
rect 92258 33070 92260 33122
rect 91756 32386 91812 32396
rect 92204 29316 92260 33070
rect 92428 34132 92484 34142
rect 92428 32786 92484 34076
rect 92428 32734 92430 32786
rect 92482 32734 92484 32786
rect 92428 32722 92484 32734
rect 92204 29250 92260 29260
rect 92652 27748 92708 35420
rect 92764 35252 92820 35262
rect 92764 34018 92820 35196
rect 92764 33966 92766 34018
rect 92818 33966 92820 34018
rect 92764 33954 92820 33966
rect 92652 27682 92708 27692
rect 92876 24836 92932 36092
rect 92988 35924 93044 35934
rect 92988 34916 93044 35868
rect 93324 35810 93380 35822
rect 93324 35758 93326 35810
rect 93378 35758 93380 35810
rect 93324 35476 93380 35758
rect 92988 34850 93044 34860
rect 93100 35420 93380 35476
rect 92876 24770 92932 24780
rect 92988 32452 93044 32462
rect 93100 32452 93156 35420
rect 93262 35308 93526 35318
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93262 35242 93526 35252
rect 93324 35140 93380 35150
rect 93324 35026 93380 35084
rect 93324 34974 93326 35026
rect 93378 34974 93380 35026
rect 93324 34962 93380 34974
rect 93262 33740 93526 33750
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93262 33674 93526 33684
rect 93660 33572 93716 36204
rect 93772 35810 93828 35822
rect 93772 35758 93774 35810
rect 93826 35758 93828 35810
rect 93772 35700 93828 35758
rect 93772 35634 93828 35644
rect 93996 35474 94052 35486
rect 93996 35422 93998 35474
rect 94050 35422 94052 35474
rect 93772 34356 93828 34366
rect 93772 34262 93828 34300
rect 93212 33516 93716 33572
rect 93212 33458 93268 33516
rect 93212 33406 93214 33458
rect 93266 33406 93268 33458
rect 93212 33394 93268 33406
rect 93996 33460 94052 35422
rect 94220 35140 94276 39200
rect 94332 37380 94388 37390
rect 94332 35924 94388 37324
rect 94332 35858 94388 35868
rect 94556 36932 94612 36942
rect 94556 36370 94612 36876
rect 94556 36318 94558 36370
rect 94610 36318 94612 36370
rect 94220 35074 94276 35084
rect 94332 35474 94388 35486
rect 94332 35422 94334 35474
rect 94386 35422 94388 35474
rect 94220 34914 94276 34926
rect 94220 34862 94222 34914
rect 94274 34862 94276 34914
rect 94220 34018 94276 34862
rect 94220 33966 94222 34018
rect 94274 33966 94276 34018
rect 93996 33394 94052 33404
rect 94108 33684 94164 33694
rect 94108 33458 94164 33628
rect 94108 33406 94110 33458
rect 94162 33406 94164 33458
rect 94108 33394 94164 33406
rect 92988 32450 93156 32452
rect 92988 32398 92990 32450
rect 93042 32398 93156 32450
rect 92988 32396 93156 32398
rect 93548 33122 93604 33134
rect 93548 33070 93550 33122
rect 93602 33070 93604 33122
rect 93548 32452 93604 33070
rect 92988 20132 93044 32396
rect 93548 32386 93604 32396
rect 93996 33124 94052 33134
rect 93262 32172 93526 32182
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93262 32106 93526 32116
rect 93996 31668 94052 33068
rect 93996 31602 94052 31612
rect 93262 30604 93526 30614
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93262 30538 93526 30548
rect 93262 29036 93526 29046
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93262 28970 93526 28980
rect 93262 27468 93526 27478
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93262 27402 93526 27412
rect 94220 26292 94276 33966
rect 94220 26226 94276 26236
rect 93262 25900 93526 25910
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93262 25834 93526 25844
rect 93262 24332 93526 24342
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93262 24266 93526 24276
rect 93262 22764 93526 22774
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93262 22698 93526 22708
rect 93262 21196 93526 21206
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93262 21130 93526 21140
rect 92988 20066 93044 20076
rect 93262 19628 93526 19638
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93262 19562 93526 19572
rect 93262 18060 93526 18070
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93262 17994 93526 18004
rect 91420 11106 91476 11116
rect 92428 17668 92484 17678
rect 90412 8372 90580 8428
rect 92428 8428 92484 17612
rect 93262 16492 93526 16502
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93262 16426 93526 16436
rect 93262 14924 93526 14934
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93262 14858 93526 14868
rect 93262 13356 93526 13366
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93262 13290 93526 13300
rect 93262 11788 93526 11798
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93262 11722 93526 11732
rect 93262 10220 93526 10230
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93262 10154 93526 10164
rect 93262 8652 93526 8662
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93262 8586 93526 8596
rect 92428 8372 92596 8428
rect 88956 8034 89012 8046
rect 88956 7982 88958 8034
rect 89010 7982 89012 8034
rect 88956 6580 89012 7982
rect 89740 7476 89796 7486
rect 88956 5346 89012 6524
rect 89068 7364 89124 7374
rect 89068 6578 89124 7308
rect 89180 7362 89236 7374
rect 89180 7310 89182 7362
rect 89234 7310 89236 7362
rect 89180 7252 89236 7310
rect 89180 6690 89236 7196
rect 89628 7362 89684 7374
rect 89628 7310 89630 7362
rect 89682 7310 89684 7362
rect 89628 7252 89684 7310
rect 89628 7186 89684 7196
rect 89740 6914 89796 7420
rect 89740 6862 89742 6914
rect 89794 6862 89796 6914
rect 89740 6850 89796 6862
rect 90412 7362 90468 8372
rect 90860 7700 90916 7710
rect 90860 7476 90916 7644
rect 90860 7410 90916 7420
rect 90412 7310 90414 7362
rect 90466 7310 90468 7362
rect 90412 6916 90468 7310
rect 91420 7364 91476 7374
rect 91420 7270 91476 7308
rect 90412 6850 90468 6860
rect 91196 6916 91252 6926
rect 91196 6822 91252 6860
rect 89180 6638 89182 6690
rect 89234 6638 89236 6690
rect 89180 6626 89236 6638
rect 91980 6692 92036 6702
rect 89068 6526 89070 6578
rect 89122 6526 89124 6578
rect 89068 6514 89124 6526
rect 91868 6580 91924 6590
rect 91868 6486 91924 6524
rect 90076 6468 90132 6478
rect 89516 6466 90132 6468
rect 89516 6414 90078 6466
rect 90130 6414 90132 6466
rect 89516 6412 90132 6414
rect 89404 5908 89460 5918
rect 89516 5908 89572 6412
rect 90076 6402 90132 6412
rect 90860 6468 90916 6478
rect 90860 6466 91364 6468
rect 90860 6414 90862 6466
rect 90914 6414 91364 6466
rect 90860 6412 91364 6414
rect 90860 6402 90916 6412
rect 90076 6132 90132 6142
rect 89628 6020 89684 6030
rect 89628 6018 89796 6020
rect 89628 5966 89630 6018
rect 89682 5966 89796 6018
rect 89628 5964 89796 5966
rect 89628 5954 89684 5964
rect 89404 5906 89572 5908
rect 89404 5854 89406 5906
rect 89458 5854 89572 5906
rect 89404 5852 89572 5854
rect 89404 5842 89460 5852
rect 88956 5294 88958 5346
rect 89010 5294 89012 5346
rect 88956 5282 89012 5294
rect 89404 5236 89460 5246
rect 89404 5142 89460 5180
rect 89516 5122 89572 5134
rect 89516 5070 89518 5122
rect 89570 5070 89572 5122
rect 89516 4676 89572 5070
rect 89516 4610 89572 4620
rect 89180 4340 89236 4350
rect 89180 4246 89236 4284
rect 89740 4338 89796 5964
rect 90076 5234 90132 6076
rect 90412 6132 90468 6142
rect 91308 6132 91364 6412
rect 91308 6076 91588 6132
rect 90412 6038 90468 6076
rect 91532 6018 91588 6076
rect 91532 5966 91534 6018
rect 91586 5966 91588 6018
rect 91532 5954 91588 5966
rect 91868 6020 91924 6030
rect 91868 5926 91924 5964
rect 90972 5908 91028 5918
rect 90972 5814 91028 5852
rect 91980 5908 92036 6636
rect 91980 5842 92036 5852
rect 92428 5794 92484 5806
rect 92428 5742 92430 5794
rect 92482 5742 92484 5794
rect 90076 5182 90078 5234
rect 90130 5182 90132 5234
rect 90076 5170 90132 5182
rect 90748 5236 90804 5246
rect 90748 5010 90804 5180
rect 91644 5236 91700 5246
rect 91644 5142 91700 5180
rect 92204 5236 92260 5246
rect 92204 5142 92260 5180
rect 90748 4958 90750 5010
rect 90802 4958 90804 5010
rect 90748 4676 90804 4958
rect 91084 5012 91140 5022
rect 91084 4918 91140 4956
rect 92428 5012 92484 5742
rect 92428 4946 92484 4956
rect 91756 4900 91812 4910
rect 91756 4898 92148 4900
rect 91756 4846 91758 4898
rect 91810 4846 92148 4898
rect 91756 4844 92148 4846
rect 91756 4834 91812 4844
rect 90748 4610 90804 4620
rect 92092 4562 92148 4844
rect 92092 4510 92094 4562
rect 92146 4510 92148 4562
rect 92092 4498 92148 4510
rect 89740 4286 89742 4338
rect 89794 4286 89796 4338
rect 89740 4274 89796 4286
rect 88620 3726 88622 3778
rect 88674 3726 88676 3778
rect 88620 3714 88676 3726
rect 91756 4228 91812 4238
rect 87948 3444 88004 3454
rect 87948 3350 88004 3388
rect 89068 3444 89124 3454
rect 89068 800 89124 3388
rect 91084 3444 91140 3454
rect 91084 3350 91140 3388
rect 91756 800 91812 4172
rect 92540 3778 92596 8316
rect 94332 7700 94388 35422
rect 94556 33684 94612 36318
rect 95004 35698 95060 35710
rect 95004 35646 95006 35698
rect 95058 35646 95060 35698
rect 94780 35588 94836 35598
rect 94780 34020 94836 35532
rect 94780 34018 94948 34020
rect 94780 33966 94782 34018
rect 94834 33966 94948 34018
rect 94780 33964 94948 33966
rect 94780 33954 94836 33964
rect 94556 33618 94612 33628
rect 94780 33124 94836 33134
rect 94780 33030 94836 33068
rect 94892 31668 94948 33964
rect 95004 33124 95060 35646
rect 95116 35252 95172 39200
rect 96012 36372 96068 39200
rect 96236 36708 96292 36718
rect 96236 36594 96292 36652
rect 96236 36542 96238 36594
rect 96290 36542 96292 36594
rect 96236 36530 96292 36542
rect 96012 36306 96068 36316
rect 96460 36148 96516 36158
rect 95116 35186 95172 35196
rect 95564 35700 95620 35710
rect 95116 34914 95172 34926
rect 95116 34862 95118 34914
rect 95170 34862 95172 34914
rect 95116 34018 95172 34862
rect 95564 34354 95620 35644
rect 95900 35586 95956 35598
rect 95900 35534 95902 35586
rect 95954 35534 95956 35586
rect 95788 35140 95844 35150
rect 95788 35026 95844 35084
rect 95788 34974 95790 35026
rect 95842 34974 95844 35026
rect 95788 34962 95844 34974
rect 95900 34916 95956 35534
rect 95900 34850 95956 34860
rect 96460 35364 96516 36092
rect 95564 34302 95566 34354
rect 95618 34302 95620 34354
rect 95564 34290 95620 34302
rect 96460 34354 96516 35308
rect 96460 34302 96462 34354
rect 96514 34302 96516 34354
rect 96460 34290 96516 34302
rect 96796 34914 96852 34926
rect 96796 34862 96798 34914
rect 96850 34862 96852 34914
rect 95116 33966 95118 34018
rect 95170 33966 95172 34018
rect 95116 33348 95172 33966
rect 96012 34018 96068 34030
rect 96012 33966 96014 34018
rect 96066 33966 96068 34018
rect 96012 33906 96068 33966
rect 96012 33854 96014 33906
rect 96066 33854 96068 33906
rect 95116 33282 95172 33292
rect 95228 33460 95284 33470
rect 95004 33058 95060 33068
rect 95228 32564 95284 33404
rect 96012 32788 96068 33854
rect 96684 33908 96740 33918
rect 96796 33908 96852 34862
rect 96908 34020 96964 39200
rect 97468 36372 97524 36382
rect 97468 36278 97524 36316
rect 97580 35700 97636 35710
rect 97468 35698 97636 35700
rect 97468 35646 97582 35698
rect 97634 35646 97636 35698
rect 97468 35644 97636 35646
rect 97244 35364 97300 35374
rect 97244 34130 97300 35308
rect 97244 34078 97246 34130
rect 97298 34078 97300 34130
rect 97244 34066 97300 34078
rect 96908 33954 96964 33964
rect 96684 33906 96852 33908
rect 96684 33854 96686 33906
rect 96738 33854 96852 33906
rect 96684 33852 96852 33854
rect 96684 33842 96740 33852
rect 97468 33460 97524 35644
rect 97580 35634 97636 35644
rect 97580 35252 97636 35262
rect 97580 35026 97636 35196
rect 97804 35140 97860 39200
rect 98364 36484 98420 36494
rect 98700 36484 98756 39200
rect 98364 36482 98532 36484
rect 98364 36430 98366 36482
rect 98418 36430 98532 36482
rect 98364 36428 98532 36430
rect 98364 36418 98420 36428
rect 97916 35812 97972 35822
rect 98252 35812 98308 35822
rect 97916 35810 98084 35812
rect 97916 35758 97918 35810
rect 97970 35758 98084 35810
rect 97916 35756 98084 35758
rect 97916 35746 97972 35756
rect 97804 35074 97860 35084
rect 97580 34974 97582 35026
rect 97634 34974 97636 35026
rect 97580 34962 97636 34974
rect 98028 34132 98084 35756
rect 98028 34066 98084 34076
rect 97916 34020 97972 34030
rect 97916 33926 97972 33964
rect 96012 32722 96068 32732
rect 97244 33404 97524 33460
rect 98252 33458 98308 35756
rect 98252 33406 98254 33458
rect 98306 33406 98308 33458
rect 97244 33122 97300 33404
rect 98252 33394 98308 33406
rect 98476 33460 98532 36428
rect 98700 36418 98756 36428
rect 99036 36372 99092 36382
rect 99036 36278 99092 36316
rect 98588 36258 98644 36270
rect 98588 36206 98590 36258
rect 98642 36206 98644 36258
rect 98588 36036 98644 36206
rect 98588 35980 98868 36036
rect 98700 35812 98756 35822
rect 98700 35718 98756 35756
rect 98588 35700 98644 35710
rect 98588 35606 98644 35644
rect 98588 34914 98644 34926
rect 98588 34862 98590 34914
rect 98642 34862 98644 34914
rect 98588 34804 98644 34862
rect 98812 34916 98868 35980
rect 99596 35588 99652 39200
rect 100156 37268 100212 37278
rect 99484 35532 99652 35588
rect 99820 36594 99876 36606
rect 99820 36542 99822 36594
rect 99874 36542 99876 36594
rect 99372 35476 99428 35486
rect 99372 35382 99428 35420
rect 99260 35140 99316 35150
rect 99260 35026 99316 35084
rect 99260 34974 99262 35026
rect 99314 34974 99316 35026
rect 99260 34962 99316 34974
rect 98812 34850 98868 34860
rect 98588 34738 98644 34748
rect 98924 34804 98980 34814
rect 98924 34354 98980 34748
rect 98924 34302 98926 34354
rect 98978 34302 98980 34354
rect 98924 34290 98980 34302
rect 99484 34020 99540 35532
rect 99708 35476 99764 35486
rect 99484 33954 99540 33964
rect 99596 35474 99764 35476
rect 99596 35422 99710 35474
rect 99762 35422 99764 35474
rect 99596 35420 99764 35422
rect 98588 33460 98644 33470
rect 98476 33458 98644 33460
rect 98476 33406 98590 33458
rect 98642 33406 98644 33458
rect 98476 33404 98644 33406
rect 97244 33070 97246 33122
rect 97298 33070 97300 33122
rect 95228 32498 95284 32508
rect 94892 31602 94948 31612
rect 94332 7634 94388 7644
rect 97244 7588 97300 33070
rect 98252 26292 98308 26302
rect 98252 8372 98308 26236
rect 98588 23380 98644 33404
rect 99484 33122 99540 33134
rect 99484 33070 99486 33122
rect 99538 33070 99540 33122
rect 99484 31948 99540 33070
rect 99036 31892 99540 31948
rect 99036 30996 99092 31892
rect 99036 30930 99092 30940
rect 98588 23314 98644 23324
rect 99596 8428 99652 35420
rect 99708 35410 99764 35420
rect 99820 34356 99876 36542
rect 99708 34300 99876 34356
rect 100156 35028 100212 37212
rect 100380 36036 100436 36046
rect 100380 35922 100436 35980
rect 100380 35870 100382 35922
rect 100434 35870 100436 35922
rect 100380 35858 100436 35870
rect 100492 35140 100548 39200
rect 100828 36484 100884 36494
rect 100828 36370 100884 36428
rect 100828 36318 100830 36370
rect 100882 36318 100884 36370
rect 100828 36306 100884 36318
rect 100492 35074 100548 35084
rect 100940 35700 100996 35710
rect 100268 35028 100324 35038
rect 100156 35026 100324 35028
rect 100156 34974 100270 35026
rect 100322 34974 100324 35026
rect 100156 34972 100324 34974
rect 99708 26404 99764 34300
rect 100044 34132 100100 34142
rect 100156 34132 100212 34972
rect 100268 34962 100324 34972
rect 100044 34130 100212 34132
rect 100044 34078 100046 34130
rect 100098 34078 100212 34130
rect 100044 34076 100212 34078
rect 100044 34066 100100 34076
rect 100492 34020 100548 34030
rect 100492 33926 100548 33964
rect 100940 33460 100996 35644
rect 101388 35252 101444 39200
rect 101612 36596 101668 36606
rect 101388 35186 101444 35196
rect 101500 36036 101556 36046
rect 101164 34916 101220 34926
rect 101164 34822 101220 34860
rect 101500 34354 101556 35980
rect 101612 35586 101668 36540
rect 102172 36258 102228 36270
rect 102172 36206 102174 36258
rect 102226 36206 102228 36258
rect 102172 36036 102228 36206
rect 102172 35970 102228 35980
rect 101612 35534 101614 35586
rect 101666 35534 101668 35586
rect 101612 35522 101668 35534
rect 102060 35476 102116 35486
rect 101500 34302 101502 34354
rect 101554 34302 101556 34354
rect 101500 34290 101556 34302
rect 101612 35252 101668 35262
rect 101052 33460 101108 33470
rect 100940 33458 101108 33460
rect 100940 33406 101054 33458
rect 101106 33406 101108 33458
rect 100940 33404 101108 33406
rect 101052 33394 101108 33404
rect 101612 33458 101668 35196
rect 101836 35140 101892 35150
rect 101836 35026 101892 35084
rect 101836 34974 101838 35026
rect 101890 34974 101892 35026
rect 101836 34962 101892 34974
rect 102060 34354 102116 35420
rect 102284 34804 102340 39200
rect 102732 36482 102788 36494
rect 102732 36430 102734 36482
rect 102786 36430 102788 36482
rect 102620 35810 102676 35822
rect 102620 35758 102622 35810
rect 102674 35758 102676 35810
rect 102396 35476 102452 35486
rect 102396 35252 102452 35420
rect 102620 35476 102676 35758
rect 102620 35410 102676 35420
rect 102396 35186 102452 35196
rect 102732 35252 102788 36430
rect 102732 35186 102788 35196
rect 102956 34916 103012 34926
rect 102284 34738 102340 34748
rect 102732 34914 103012 34916
rect 102732 34862 102958 34914
rect 103010 34862 103012 34914
rect 102732 34860 103012 34862
rect 102060 34302 102062 34354
rect 102114 34302 102116 34354
rect 102060 34290 102116 34302
rect 102620 34244 102676 34254
rect 102620 34150 102676 34188
rect 101612 33406 101614 33458
rect 101666 33406 101668 33458
rect 101612 33394 101668 33406
rect 102732 33458 102788 34860
rect 102956 34850 103012 34860
rect 103180 34468 103236 39200
rect 103628 36484 103684 36494
rect 103628 36390 103684 36428
rect 104076 36372 104132 39200
rect 104748 37828 104804 37838
rect 103964 36316 104076 36372
rect 103740 35700 103796 35710
rect 103628 35026 103684 35038
rect 103628 34974 103630 35026
rect 103682 34974 103684 35026
rect 103628 34804 103684 34974
rect 103628 34738 103684 34748
rect 103180 34402 103236 34412
rect 103180 34244 103236 34254
rect 103180 34130 103236 34188
rect 103180 34078 103182 34130
rect 103234 34078 103236 34130
rect 103180 34066 103236 34078
rect 102732 33406 102734 33458
rect 102786 33406 102788 33458
rect 99820 33236 99876 33246
rect 100268 33236 100324 33246
rect 99820 33234 100324 33236
rect 99820 33182 99822 33234
rect 99874 33182 100270 33234
rect 100322 33182 100324 33234
rect 99820 33180 100324 33182
rect 99820 33170 99876 33180
rect 100268 32788 100324 33180
rect 100268 32722 100324 32732
rect 102396 32788 102452 32798
rect 99708 26338 99764 26348
rect 98252 8306 98308 8316
rect 99484 8372 99652 8428
rect 101836 24388 101892 24398
rect 97244 7522 97300 7532
rect 99260 7474 99316 7486
rect 99260 7422 99262 7474
rect 99314 7422 99316 7474
rect 92876 7364 92932 7374
rect 92876 4562 92932 7308
rect 93262 7084 93526 7094
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93262 7018 93526 7028
rect 99148 6916 99204 6926
rect 99260 6916 99316 7422
rect 99148 6914 99316 6916
rect 99148 6862 99150 6914
rect 99202 6862 99316 6914
rect 99148 6860 99316 6862
rect 99484 6916 99540 8372
rect 101724 7700 101780 7710
rect 99148 6850 99204 6860
rect 97132 6804 97188 6814
rect 99484 6784 99540 6860
rect 99596 7586 99652 7598
rect 99596 7534 99598 7586
rect 99650 7534 99652 7586
rect 93100 6692 93156 6702
rect 93100 6598 93156 6636
rect 93660 6580 93716 6590
rect 93660 6466 93716 6524
rect 93660 6414 93662 6466
rect 93714 6414 93716 6466
rect 93262 5516 93526 5526
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93262 5450 93526 5460
rect 93660 5348 93716 6414
rect 95564 6020 95620 6030
rect 93660 5282 93716 5292
rect 94892 5794 94948 5806
rect 94892 5742 94894 5794
rect 94946 5742 94948 5794
rect 93100 5236 93156 5246
rect 93100 5142 93156 5180
rect 94556 5236 94612 5246
rect 93660 5122 93716 5134
rect 93660 5070 93662 5122
rect 93714 5070 93716 5122
rect 93660 5012 93716 5070
rect 93660 4946 93716 4956
rect 94220 5012 94276 5022
rect 94220 4918 94276 4956
rect 94556 5010 94612 5180
rect 94892 5124 94948 5742
rect 94892 5058 94948 5068
rect 95228 5124 95284 5134
rect 95228 5030 95284 5068
rect 95564 5122 95620 5964
rect 95564 5070 95566 5122
rect 95618 5070 95620 5122
rect 95564 5058 95620 5070
rect 94556 4958 94558 5010
rect 94610 4958 94612 5010
rect 94556 4946 94612 4958
rect 97132 4564 97188 6748
rect 98476 6692 98532 6702
rect 98476 6598 98532 6636
rect 98700 5348 98756 5358
rect 98700 5254 98756 5292
rect 92876 4510 92878 4562
rect 92930 4510 92932 4562
rect 92876 4498 92932 4510
rect 96460 4562 97188 4564
rect 96460 4510 97134 4562
rect 97186 4510 97188 4562
rect 96460 4508 97188 4510
rect 94556 4338 94612 4350
rect 94556 4286 94558 4338
rect 94610 4286 94612 4338
rect 93436 4228 93492 4238
rect 93436 4134 93492 4172
rect 93262 3948 93526 3958
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93262 3882 93526 3892
rect 94556 3892 94612 4286
rect 96460 4338 96516 4508
rect 97132 4498 97188 4508
rect 97804 5236 97860 5246
rect 97804 4450 97860 5180
rect 98364 5236 98420 5246
rect 97916 4898 97972 4910
rect 97916 4846 97918 4898
rect 97970 4846 97972 4898
rect 97916 4562 97972 4846
rect 97916 4510 97918 4562
rect 97970 4510 97972 4562
rect 97916 4498 97972 4510
rect 98364 4562 98420 5180
rect 98364 4510 98366 4562
rect 98418 4510 98420 4562
rect 98364 4498 98420 4510
rect 97804 4398 97806 4450
rect 97858 4398 97860 4450
rect 97804 4386 97860 4398
rect 96460 4286 96462 4338
rect 96514 4286 96516 4338
rect 96460 4274 96516 4286
rect 99036 4340 99092 4350
rect 99036 4246 99092 4284
rect 99484 4340 99540 4350
rect 99596 4340 99652 7534
rect 100268 7364 100324 7374
rect 100268 6692 100324 7308
rect 100044 6578 100100 6590
rect 100044 6526 100046 6578
rect 100098 6526 100100 6578
rect 100268 6560 100324 6636
rect 101052 6916 101108 6926
rect 101052 6690 101108 6860
rect 101724 6692 101780 7644
rect 101052 6638 101054 6690
rect 101106 6638 101108 6690
rect 101052 6626 101108 6638
rect 101276 6636 101780 6692
rect 100044 4564 100100 6526
rect 101276 5906 101332 6636
rect 101276 5854 101278 5906
rect 101330 5854 101332 5906
rect 101276 5842 101332 5854
rect 101612 6466 101668 6478
rect 101612 6414 101614 6466
rect 101666 6414 101668 6466
rect 100044 4498 100100 4508
rect 100156 5794 100212 5806
rect 100156 5742 100158 5794
rect 100210 5742 100212 5794
rect 100044 4340 100100 4350
rect 99596 4338 100100 4340
rect 99596 4286 100046 4338
rect 100098 4286 100100 4338
rect 99596 4284 100100 4286
rect 99484 4246 99540 4284
rect 100044 4274 100100 4284
rect 94556 3826 94612 3836
rect 95788 4226 95844 4238
rect 95788 4174 95790 4226
rect 95842 4174 95844 4226
rect 92540 3726 92542 3778
rect 92594 3726 92596 3778
rect 92540 3714 92596 3726
rect 91868 3444 91924 3454
rect 91868 3350 91924 3388
rect 93100 3444 93156 3454
rect 93100 800 93156 3388
rect 94668 3444 94724 3454
rect 94668 3350 94724 3388
rect 95788 800 95844 4174
rect 95900 3892 95956 3902
rect 95900 3666 95956 3836
rect 95900 3614 95902 3666
rect 95954 3614 95956 3666
rect 95900 3602 95956 3614
rect 98812 3668 98868 3678
rect 98812 3574 98868 3612
rect 96236 3444 96292 3454
rect 96236 3350 96292 3388
rect 96908 3444 96964 3454
rect 97468 3444 97524 3454
rect 96908 3442 97524 3444
rect 96908 3390 96910 3442
rect 96962 3390 97470 3442
rect 97522 3390 97524 3442
rect 96908 3388 97524 3390
rect 96908 3378 96964 3388
rect 97132 800 97188 3388
rect 97468 3378 97524 3388
rect 100156 2884 100212 5742
rect 101612 4452 101668 6414
rect 101724 6130 101780 6636
rect 101724 6078 101726 6130
rect 101778 6078 101780 6130
rect 101724 6066 101780 6078
rect 101612 4386 101668 4396
rect 101836 3668 101892 24332
rect 102396 22708 102452 32732
rect 102732 31332 102788 33406
rect 102732 31266 102788 31276
rect 102396 22642 102452 22652
rect 103740 12740 103796 35644
rect 103852 34468 103908 34478
rect 103852 34018 103908 34412
rect 103852 33966 103854 34018
rect 103906 33966 103908 34018
rect 103852 33954 103908 33966
rect 103964 33460 104020 36316
rect 104076 36306 104132 36316
rect 104412 36594 104468 36606
rect 104412 36542 104414 36594
rect 104466 36542 104468 36594
rect 104076 35810 104132 35822
rect 104076 35758 104078 35810
rect 104130 35758 104132 35810
rect 104076 35476 104132 35758
rect 104076 35410 104132 35420
rect 104076 33460 104132 33470
rect 103964 33458 104132 33460
rect 103964 33406 104078 33458
rect 104130 33406 104132 33458
rect 103964 33404 104132 33406
rect 104076 33394 104132 33404
rect 104412 31948 104468 36542
rect 104748 34804 104804 37772
rect 104748 34738 104804 34748
rect 104860 36260 104916 36270
rect 104860 34914 104916 36204
rect 104860 34862 104862 34914
rect 104914 34862 104916 34914
rect 104860 33570 104916 34862
rect 104972 34020 105028 39200
rect 105756 37716 105812 37726
rect 105644 37268 105700 37278
rect 105308 36372 105364 36382
rect 105308 36278 105364 36316
rect 105084 36036 105140 36046
rect 105084 35922 105140 35980
rect 105084 35870 105086 35922
rect 105138 35870 105140 35922
rect 105084 35858 105140 35870
rect 105532 35700 105588 35710
rect 105532 35606 105588 35644
rect 105420 34914 105476 34926
rect 105420 34862 105422 34914
rect 105474 34862 105476 34914
rect 104972 33954 105028 33964
rect 105196 34580 105252 34590
rect 105196 34130 105252 34524
rect 105420 34244 105476 34862
rect 105420 34178 105476 34188
rect 105196 34078 105198 34130
rect 105250 34078 105252 34130
rect 104860 33518 104862 33570
rect 104914 33518 104916 33570
rect 104860 33506 104916 33518
rect 104972 33460 105028 33470
rect 105196 33460 105252 34078
rect 105644 33796 105700 37212
rect 105756 36484 105812 37660
rect 105756 36418 105812 36428
rect 105868 35812 105924 39200
rect 106316 36260 106372 36270
rect 106316 36166 106372 36204
rect 105868 35746 105924 35756
rect 106092 35586 106148 35598
rect 106092 35534 106094 35586
rect 106146 35534 106148 35586
rect 106092 35364 106148 35534
rect 106092 35298 106148 35308
rect 106092 34804 106148 34814
rect 105868 34020 105924 34030
rect 105868 33926 105924 33964
rect 105644 33730 105700 33740
rect 104972 33458 105252 33460
rect 104972 33406 104974 33458
rect 105026 33406 105252 33458
rect 104972 33404 105252 33406
rect 105420 33570 105476 33582
rect 105420 33518 105422 33570
rect 105474 33518 105476 33570
rect 105420 33458 105476 33518
rect 105420 33406 105422 33458
rect 105474 33406 105476 33458
rect 104972 33394 105028 33404
rect 104300 31892 104468 31948
rect 104300 30100 104356 31892
rect 104300 30034 104356 30044
rect 103740 12674 103796 12684
rect 104972 28644 105028 28654
rect 101948 5236 102004 5246
rect 101948 5142 102004 5180
rect 102508 5236 102564 5246
rect 102508 5142 102564 5180
rect 104188 5124 104244 5134
rect 103852 5122 104244 5124
rect 103852 5070 104190 5122
rect 104242 5070 104244 5122
rect 103852 5068 104244 5070
rect 102060 4898 102116 4910
rect 102060 4846 102062 4898
rect 102114 4846 102116 4898
rect 102060 4564 102116 4846
rect 102060 4498 102116 4508
rect 102508 4564 102564 4574
rect 102508 4470 102564 4508
rect 103180 4452 103236 4462
rect 103180 4358 103236 4396
rect 101836 3602 101892 3612
rect 102844 3668 102900 3678
rect 102844 3574 102900 3612
rect 100940 3444 100996 3454
rect 101500 3444 101556 3454
rect 100940 3442 101556 3444
rect 100940 3390 100942 3442
rect 100994 3390 101502 3442
rect 101554 3390 101556 3442
rect 100940 3388 101556 3390
rect 100940 3378 100996 3388
rect 99820 2828 100212 2884
rect 99820 800 99876 2828
rect 101164 800 101220 3388
rect 101500 3378 101556 3388
rect 103852 800 103908 5068
rect 104188 5058 104244 5068
rect 104972 3668 105028 28588
rect 105420 23268 105476 33406
rect 105868 33460 105924 33470
rect 106092 33460 106148 34748
rect 106652 34802 106708 34814
rect 106652 34750 106654 34802
rect 106706 34750 106708 34802
rect 105868 33458 106148 33460
rect 105868 33406 105870 33458
rect 105922 33406 106148 33458
rect 105868 33404 106148 33406
rect 106316 34244 106372 34254
rect 106316 33458 106372 34188
rect 106652 34244 106708 34750
rect 106652 34178 106708 34188
rect 106764 34020 106820 39200
rect 106988 37156 107044 37166
rect 106876 36482 106932 36494
rect 106876 36430 106878 36482
rect 106930 36430 106932 36482
rect 106876 35140 106932 36430
rect 106876 35074 106932 35084
rect 106764 33954 106820 33964
rect 106876 34914 106932 34926
rect 106876 34862 106878 34914
rect 106930 34862 106932 34914
rect 106876 33572 106932 34862
rect 106876 33506 106932 33516
rect 106988 34130 107044 37100
rect 107660 36372 107716 39200
rect 107884 37940 107940 37950
rect 107884 36594 107940 37884
rect 107884 36542 107886 36594
rect 107938 36542 107940 36594
rect 107884 36530 107940 36542
rect 107660 36306 107716 36316
rect 107100 35812 107156 35822
rect 107100 35718 107156 35756
rect 108444 35810 108500 35822
rect 108444 35758 108446 35810
rect 108498 35758 108500 35810
rect 108108 35698 108164 35710
rect 108108 35646 108110 35698
rect 108162 35646 108164 35698
rect 107436 35140 107492 35150
rect 106988 34078 106990 34130
rect 107042 34078 107044 34130
rect 106316 33406 106318 33458
rect 106370 33406 106372 33458
rect 105868 33394 105924 33404
rect 106316 33394 106372 33406
rect 106764 33348 106820 33358
rect 106988 33348 107044 34078
rect 106764 33346 107044 33348
rect 106764 33294 106766 33346
rect 106818 33294 107044 33346
rect 106764 33292 107044 33294
rect 107212 34690 107268 34702
rect 107212 34638 107214 34690
rect 107266 34638 107268 34690
rect 106764 33282 106820 33292
rect 106652 33012 106708 33022
rect 105756 32340 105812 32350
rect 105756 28644 105812 32284
rect 105756 28578 105812 28588
rect 105420 23202 105476 23212
rect 106652 26180 106708 32956
rect 105756 7140 105812 7150
rect 105756 5236 105812 7084
rect 105308 5234 105812 5236
rect 105308 5182 105758 5234
rect 105810 5182 105812 5234
rect 105308 5180 105812 5182
rect 105308 5122 105364 5180
rect 105756 5170 105812 5180
rect 105308 5070 105310 5122
rect 105362 5070 105364 5122
rect 105308 5058 105364 5070
rect 104972 3602 105028 3612
rect 106652 3666 106708 26124
rect 107212 6132 107268 34638
rect 107436 34468 107492 35084
rect 107436 34402 107492 34412
rect 107884 34802 107940 34814
rect 107884 34750 107886 34802
rect 107938 34750 107940 34802
rect 107660 34020 107716 34030
rect 107660 33926 107716 33964
rect 107884 34020 107940 34750
rect 107660 33572 107716 33582
rect 107660 33458 107716 33516
rect 107660 33406 107662 33458
rect 107714 33406 107716 33458
rect 107660 33394 107716 33406
rect 107548 31556 107604 31566
rect 107548 24388 107604 31500
rect 107548 24322 107604 24332
rect 107884 23044 107940 33964
rect 107996 33460 108052 33470
rect 108108 33460 108164 35646
rect 108444 35364 108500 35758
rect 108444 35298 108500 35308
rect 108556 35140 108612 39200
rect 108892 36372 108948 36382
rect 108948 36316 109060 36372
rect 108892 36278 108948 36316
rect 108892 35812 108948 35822
rect 108892 35718 108948 35756
rect 108556 35074 108612 35084
rect 107996 33458 108164 33460
rect 107996 33406 107998 33458
rect 108050 33406 108164 33458
rect 107996 33404 108164 33406
rect 108220 34690 108276 34702
rect 108220 34638 108222 34690
rect 108274 34638 108276 34690
rect 107996 32004 108052 33404
rect 108220 33348 108276 34638
rect 109004 34356 109060 36316
rect 109452 35812 109508 39200
rect 109452 35746 109508 35756
rect 109676 38500 109732 38510
rect 109676 35586 109732 38444
rect 109900 36484 109956 36494
rect 109900 36370 109956 36428
rect 109900 36318 109902 36370
rect 109954 36318 109956 36370
rect 109900 36306 109956 36318
rect 110236 36370 110292 36382
rect 110236 36318 110238 36370
rect 110290 36318 110292 36370
rect 109676 35534 109678 35586
rect 109730 35534 109732 35586
rect 109676 35522 109732 35534
rect 110124 35812 110180 35822
rect 109788 35140 109844 35150
rect 109788 35026 109844 35084
rect 109788 34974 109790 35026
rect 109842 34974 109844 35026
rect 109788 34962 109844 34974
rect 109004 34290 109060 34300
rect 109228 34914 109284 34926
rect 109228 34862 109230 34914
rect 109282 34862 109284 34914
rect 109228 34354 109284 34862
rect 109228 34302 109230 34354
rect 109282 34302 109284 34354
rect 109228 34132 109284 34302
rect 109564 34356 109620 34366
rect 109564 34262 109620 34300
rect 110124 34354 110180 35756
rect 110124 34302 110126 34354
rect 110178 34302 110180 34354
rect 110124 34290 110180 34302
rect 109228 34066 109284 34076
rect 110236 34132 110292 36318
rect 110348 35140 110404 39200
rect 110348 35074 110404 35084
rect 110572 37044 110628 37054
rect 110236 34066 110292 34076
rect 110460 34132 110516 34142
rect 108668 34020 108724 34030
rect 108668 33926 108724 33964
rect 108220 33282 108276 33292
rect 107996 31938 108052 31948
rect 107884 22978 107940 22988
rect 108556 24500 108612 24510
rect 108556 12740 108612 24444
rect 108556 8428 108612 12684
rect 110460 8708 110516 34076
rect 110572 33908 110628 36988
rect 111244 36372 111300 39200
rect 111580 38052 111636 38062
rect 111580 36594 111636 37996
rect 111580 36542 111582 36594
rect 111634 36542 111636 36594
rect 111580 36530 111636 36542
rect 111244 36306 111300 36316
rect 110684 36260 110740 36270
rect 110684 36166 110740 36204
rect 111672 36092 111936 36102
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111672 36026 111936 36036
rect 111356 35924 111412 35934
rect 110908 35812 110964 35822
rect 110908 35718 110964 35756
rect 110908 35476 110964 35486
rect 110908 34914 110964 35420
rect 110908 34862 110910 34914
rect 110962 34862 110964 34914
rect 110908 34850 110964 34862
rect 110908 34356 110964 34366
rect 110908 34262 110964 34300
rect 111356 34354 111412 35868
rect 111692 35924 111748 35934
rect 111692 35810 111748 35868
rect 111692 35758 111694 35810
rect 111746 35758 111748 35810
rect 111692 35746 111748 35758
rect 112028 35810 112084 35822
rect 112028 35758 112030 35810
rect 112082 35758 112084 35810
rect 112028 35252 112084 35758
rect 112028 35186 112084 35196
rect 111580 35140 111636 35150
rect 111580 35026 111636 35084
rect 111580 34974 111582 35026
rect 111634 34974 111636 35026
rect 111580 34962 111636 34974
rect 111672 34524 111936 34534
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111672 34458 111936 34468
rect 111356 34302 111358 34354
rect 111410 34302 111412 34354
rect 111356 34290 111412 34302
rect 111916 34244 111972 34254
rect 111916 34132 111972 34188
rect 111916 34130 112084 34132
rect 111916 34078 111918 34130
rect 111970 34078 112084 34130
rect 111916 34076 112084 34078
rect 111916 34066 111972 34076
rect 110572 33842 110628 33852
rect 111916 33908 111972 33918
rect 111916 33458 111972 33852
rect 112028 33796 112084 34076
rect 112028 33730 112084 33740
rect 112140 33572 112196 39200
rect 112588 36372 112644 36382
rect 112588 36278 112644 36316
rect 113036 35812 113092 39200
rect 113260 38724 113316 38734
rect 113036 35746 113092 35756
rect 113148 37604 113204 37614
rect 113148 34802 113204 37548
rect 113260 35586 113316 38668
rect 113932 36932 113988 39200
rect 113932 36876 114100 36932
rect 113260 35534 113262 35586
rect 113314 35534 113316 35586
rect 113260 35522 113316 35534
rect 113596 36370 113652 36382
rect 113596 36318 113598 36370
rect 113650 36318 113652 36370
rect 113148 34750 113150 34802
rect 113202 34750 113204 34802
rect 112140 33506 112196 33516
rect 112476 34020 112532 34030
rect 111916 33406 111918 33458
rect 111970 33406 111972 33458
rect 111916 33394 111972 33406
rect 112364 33348 112420 33358
rect 112364 33254 112420 33292
rect 111672 32956 111936 32966
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111672 32890 111936 32900
rect 111672 31388 111936 31398
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111672 31322 111936 31332
rect 111672 29820 111936 29830
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111672 29754 111936 29764
rect 112476 29540 112532 33964
rect 113148 33908 113204 34750
rect 113484 34802 113540 34814
rect 113484 34750 113486 34802
rect 113538 34750 113540 34802
rect 113484 34580 113540 34750
rect 113484 34514 113540 34524
rect 113372 34242 113428 34254
rect 113372 34190 113374 34242
rect 113426 34190 113428 34242
rect 113372 34020 113428 34190
rect 113372 33954 113428 33964
rect 113148 33842 113204 33852
rect 113036 33572 113092 33582
rect 113036 33458 113092 33516
rect 113036 33406 113038 33458
rect 113090 33406 113092 33458
rect 113036 33394 113092 33406
rect 113596 32340 113652 36318
rect 113932 36258 113988 36270
rect 113932 36206 113934 36258
rect 113986 36206 113988 36258
rect 113932 35924 113988 36206
rect 113932 35858 113988 35868
rect 114044 35140 114100 36876
rect 114380 36372 114436 36382
rect 114380 36278 114436 36316
rect 114828 36372 114884 39200
rect 114828 36306 114884 36316
rect 115500 36594 115556 36606
rect 115500 36542 115502 36594
rect 115554 36542 115556 36594
rect 115052 36148 115108 36158
rect 114268 35812 114324 35822
rect 114268 35718 114324 35756
rect 114044 35074 114100 35084
rect 114828 35252 114884 35262
rect 113820 34916 113876 34926
rect 113820 34822 113876 34860
rect 114604 34916 114660 34926
rect 114156 34692 114212 34702
rect 113932 34690 114212 34692
rect 113932 34638 114158 34690
rect 114210 34638 114212 34690
rect 113932 34636 114212 34638
rect 113820 34244 113876 34254
rect 113820 33796 113876 34188
rect 113820 33730 113876 33740
rect 113596 32274 113652 32284
rect 112476 29474 112532 29484
rect 111672 28252 111936 28262
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111672 28186 111936 28196
rect 111672 26684 111936 26694
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111672 26618 111936 26628
rect 111672 25116 111936 25126
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111672 25050 111936 25060
rect 111672 23548 111936 23558
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111672 23482 111936 23492
rect 113260 22708 113316 22718
rect 111672 21980 111936 21990
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111672 21914 111936 21924
rect 111672 20412 111936 20422
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111672 20346 111936 20356
rect 111672 18844 111936 18854
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111672 18778 111936 18788
rect 111672 17276 111936 17286
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111672 17210 111936 17220
rect 111672 15708 111936 15718
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111672 15642 111936 15652
rect 111672 14140 111936 14150
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111672 14074 111936 14084
rect 111672 12572 111936 12582
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111672 12506 111936 12516
rect 111672 11004 111936 11014
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111672 10938 111936 10948
rect 111672 9436 111936 9446
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111672 9370 111936 9380
rect 110460 8642 110516 8652
rect 110460 8484 110516 8494
rect 108556 8372 108836 8428
rect 107212 6066 107268 6076
rect 107884 6132 107940 6142
rect 107884 6038 107940 6076
rect 108556 6020 108612 6030
rect 108108 6018 108612 6020
rect 108108 5966 108558 6018
rect 108610 5966 108612 6018
rect 108108 5964 108612 5966
rect 107548 5236 107604 5246
rect 107548 4562 107604 5180
rect 107548 4510 107550 4562
rect 107602 4510 107604 4562
rect 107548 4498 107604 4510
rect 107884 5124 107940 5134
rect 106652 3614 106654 3666
rect 106706 3614 106708 3666
rect 106652 3602 106708 3614
rect 104972 3444 105028 3454
rect 105532 3444 105588 3454
rect 104972 3442 105588 3444
rect 104972 3390 104974 3442
rect 105026 3390 105534 3442
rect 105586 3390 105588 3442
rect 104972 3388 105588 3390
rect 104972 3378 105028 3388
rect 105196 800 105252 3388
rect 105532 3378 105588 3388
rect 107884 800 107940 5068
rect 108108 5122 108164 5964
rect 108556 5954 108612 5964
rect 108108 5070 108110 5122
rect 108162 5070 108164 5122
rect 108108 5058 108164 5070
rect 108220 5796 108276 5806
rect 108220 5236 108276 5740
rect 108220 4338 108276 5180
rect 108220 4286 108222 4338
rect 108274 4286 108276 4338
rect 108220 4274 108276 4286
rect 108332 4898 108388 4910
rect 108332 4846 108334 4898
rect 108386 4846 108388 4898
rect 108332 4340 108388 4846
rect 108556 4340 108612 4350
rect 108332 4338 108612 4340
rect 108332 4286 108558 4338
rect 108610 4286 108612 4338
rect 108332 4284 108612 4286
rect 108556 4274 108612 4284
rect 108332 4116 108388 4126
rect 108332 3666 108388 4060
rect 108332 3614 108334 3666
rect 108386 3614 108388 3666
rect 108332 3602 108388 3614
rect 108780 3668 108836 8372
rect 110348 6580 110404 6590
rect 108892 6132 108948 6142
rect 108892 5906 108948 6076
rect 110348 6130 110404 6524
rect 110348 6078 110350 6130
rect 110402 6078 110404 6130
rect 109676 6018 109732 6030
rect 109676 5966 109678 6018
rect 109730 5966 109732 6018
rect 108892 5854 108894 5906
rect 108946 5854 108948 5906
rect 108892 5842 108948 5854
rect 109564 5908 109620 5918
rect 109564 5814 109620 5852
rect 109228 5124 109284 5134
rect 109228 5030 109284 5068
rect 109676 5012 109732 5966
rect 110348 5908 110404 6078
rect 110460 6466 110516 8428
rect 111672 7868 111936 7878
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111672 7802 111936 7812
rect 113036 7362 113092 7374
rect 113036 7310 113038 7362
rect 113090 7310 113092 7362
rect 111580 6690 111636 6702
rect 111580 6638 111582 6690
rect 111634 6638 111636 6690
rect 111580 6580 111636 6638
rect 113036 6692 113092 7310
rect 112252 6580 112308 6590
rect 111580 6514 111636 6524
rect 112140 6578 112308 6580
rect 112140 6526 112254 6578
rect 112306 6526 112308 6578
rect 112140 6524 112308 6526
rect 110460 6414 110462 6466
rect 110514 6414 110516 6466
rect 110460 6132 110516 6414
rect 110460 6066 110516 6076
rect 111020 6466 111076 6478
rect 111020 6414 111022 6466
rect 111074 6414 111076 6466
rect 111020 6132 111076 6414
rect 111672 6300 111936 6310
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111672 6234 111936 6244
rect 111020 6066 111076 6076
rect 112028 6020 112084 6030
rect 112028 5926 112084 5964
rect 110348 5842 110404 5852
rect 110684 5794 110740 5806
rect 110684 5742 110686 5794
rect 110738 5742 110740 5794
rect 110348 5572 110404 5582
rect 110348 5122 110404 5516
rect 110348 5070 110350 5122
rect 110402 5070 110404 5122
rect 110348 5058 110404 5070
rect 109676 4946 109732 4956
rect 110684 5012 110740 5742
rect 111132 5794 111188 5806
rect 111132 5742 111134 5794
rect 111186 5742 111188 5794
rect 110684 4228 110740 4956
rect 111020 5684 111076 5694
rect 111020 5010 111076 5628
rect 111132 5572 111188 5742
rect 111132 5506 111188 5516
rect 111020 4958 111022 5010
rect 111074 4958 111076 5010
rect 111020 4946 111076 4958
rect 112028 5122 112084 5134
rect 112028 5070 112030 5122
rect 112082 5070 112084 5122
rect 111356 4900 111412 4910
rect 111356 4806 111412 4844
rect 111672 4732 111936 4742
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111672 4666 111936 4676
rect 111132 4564 111188 4574
rect 111132 4562 111636 4564
rect 111132 4510 111134 4562
rect 111186 4510 111636 4562
rect 111132 4508 111636 4510
rect 111132 4498 111188 4508
rect 110684 4162 110740 4172
rect 111580 3780 111636 4508
rect 112028 4340 112084 5070
rect 112028 4246 112084 4284
rect 111692 4228 111748 4238
rect 111692 4134 111748 4172
rect 111692 3780 111748 3790
rect 111580 3778 111748 3780
rect 111580 3726 111694 3778
rect 111746 3726 111748 3778
rect 111580 3724 111748 3726
rect 111692 3714 111748 3724
rect 108780 3602 108836 3612
rect 110572 3668 110628 3678
rect 110572 3574 110628 3612
rect 111804 3556 111860 3566
rect 111804 3462 111860 3500
rect 108892 3444 108948 3454
rect 109452 3444 109508 3454
rect 108892 3442 109508 3444
rect 108892 3390 108894 3442
rect 108946 3390 109454 3442
rect 109506 3390 109508 3442
rect 108892 3388 109508 3390
rect 108892 3378 108948 3388
rect 109228 800 109284 3388
rect 109452 3378 109508 3388
rect 111672 3164 111936 3174
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111672 3098 111936 3108
rect 112140 980 112196 6524
rect 112252 6514 112308 6524
rect 112364 6018 112420 6030
rect 112364 5966 112366 6018
rect 112418 5966 112420 6018
rect 112364 5122 112420 5966
rect 112364 5070 112366 5122
rect 112418 5070 112420 5122
rect 112364 5058 112420 5070
rect 113036 4340 113092 6636
rect 113036 4246 113092 4284
rect 112588 4116 112644 4126
rect 112588 3780 112644 4060
rect 112364 3556 112420 3566
rect 112364 3442 112420 3500
rect 112588 3554 112644 3724
rect 113260 3666 113316 22652
rect 113932 13412 113988 34636
rect 114156 34626 114212 34636
rect 114156 34132 114212 34142
rect 114156 34038 114212 34076
rect 114492 33906 114548 33918
rect 114492 33854 114494 33906
rect 114546 33854 114548 33906
rect 114044 33122 114100 33134
rect 114044 33070 114046 33122
rect 114098 33070 114100 33122
rect 114044 32340 114100 33070
rect 114044 32274 114100 32284
rect 113932 13346 113988 13356
rect 114492 8428 114548 33854
rect 114604 33458 114660 34860
rect 114828 34914 114884 35196
rect 114828 34862 114830 34914
rect 114882 34862 114884 34914
rect 114828 34850 114884 34862
rect 115052 34354 115108 36092
rect 115388 36036 115444 36046
rect 115052 34302 115054 34354
rect 115106 34302 115108 34354
rect 115052 34132 115108 34302
rect 115052 34066 115108 34076
rect 115276 35698 115332 35710
rect 115276 35646 115278 35698
rect 115330 35646 115332 35698
rect 115276 34692 115332 35646
rect 115388 34916 115444 35980
rect 115500 35364 115556 36542
rect 115612 35810 115668 35822
rect 115612 35758 115614 35810
rect 115666 35758 115668 35810
rect 115612 35700 115668 35758
rect 115612 35634 115668 35644
rect 115500 35308 115668 35364
rect 115500 35140 115556 35150
rect 115500 35026 115556 35084
rect 115500 34974 115502 35026
rect 115554 34974 115556 35026
rect 115500 34962 115556 34974
rect 115388 34850 115444 34860
rect 114604 33406 114606 33458
rect 114658 33406 114660 33458
rect 114604 33394 114660 33406
rect 115276 21028 115332 34636
rect 115612 32564 115668 35308
rect 115724 34020 115780 39200
rect 116508 36372 116564 36382
rect 116508 36278 116564 36316
rect 116060 35812 116116 35822
rect 116060 35718 116116 35756
rect 115948 35700 116004 35710
rect 115948 34130 116004 35644
rect 116620 35140 116676 39200
rect 117180 37492 117236 37502
rect 116620 35074 116676 35084
rect 116844 35586 116900 35598
rect 116844 35534 116846 35586
rect 116898 35534 116900 35586
rect 115948 34078 115950 34130
rect 116002 34078 116004 34130
rect 115948 34066 116004 34078
rect 115724 33954 115780 33964
rect 116620 34020 116676 34030
rect 116620 33926 116676 33964
rect 116844 32676 116900 35534
rect 117068 35140 117124 35150
rect 116956 34692 117012 34702
rect 116956 34598 117012 34636
rect 117068 33458 117124 35084
rect 117180 34356 117236 37436
rect 117516 37156 117572 39200
rect 117292 37100 117572 37156
rect 117628 38388 117684 38398
rect 117628 37156 117684 38332
rect 117292 35252 117348 37100
rect 117628 37090 117684 37100
rect 118412 36708 118468 39200
rect 118412 36642 118468 36652
rect 119196 37156 119252 37166
rect 117516 36372 117572 36382
rect 117292 35186 117348 35196
rect 117404 36370 117572 36372
rect 117404 36318 117518 36370
rect 117570 36318 117572 36370
rect 117404 36316 117572 36318
rect 117180 34290 117236 34300
rect 117068 33406 117070 33458
rect 117122 33406 117124 33458
rect 117068 33394 117124 33406
rect 116844 32610 116900 32620
rect 117404 33122 117460 36316
rect 117516 36306 117572 36316
rect 118300 36372 118356 36382
rect 118300 36278 118356 36316
rect 117852 36260 117908 36270
rect 117740 36258 117908 36260
rect 117740 36206 117854 36258
rect 117906 36206 117908 36258
rect 117740 36204 117908 36206
rect 117740 34914 117796 36204
rect 117852 36194 117908 36204
rect 117852 35810 117908 35822
rect 117852 35758 117854 35810
rect 117906 35758 117908 35810
rect 117852 35140 117908 35758
rect 119196 35810 119252 37100
rect 119196 35758 119198 35810
rect 119250 35758 119252 35810
rect 119196 35746 119252 35758
rect 119084 35698 119140 35710
rect 119084 35646 119086 35698
rect 119138 35646 119140 35698
rect 117852 35074 117908 35084
rect 118412 35252 118468 35262
rect 118412 35026 118468 35196
rect 118412 34974 118414 35026
rect 118466 34974 118468 35026
rect 118412 34962 118468 34974
rect 117740 34862 117742 34914
rect 117794 34862 117796 34914
rect 117740 34850 117796 34862
rect 119084 34580 119140 35646
rect 117740 34356 117796 34366
rect 117740 34262 117796 34300
rect 118076 34130 118132 34142
rect 118076 34078 118078 34130
rect 118130 34078 118132 34130
rect 118076 34020 118132 34078
rect 118524 34020 118580 34030
rect 119084 34020 119140 34524
rect 118076 34018 118580 34020
rect 118076 33966 118526 34018
rect 118578 33966 118580 34018
rect 118076 33964 118580 33966
rect 118524 33572 118580 33964
rect 118524 33506 118580 33516
rect 118972 33964 119140 34020
rect 119308 34018 119364 39200
rect 119420 36596 119476 36606
rect 119420 36502 119476 36540
rect 120092 36260 120148 36270
rect 119868 35476 119924 35486
rect 119868 35382 119924 35420
rect 119420 35140 119476 35150
rect 119420 34804 119476 35084
rect 119980 35140 120036 35150
rect 119980 34914 120036 35084
rect 119980 34862 119982 34914
rect 120034 34862 120036 34914
rect 119868 34804 119924 34814
rect 119420 34738 119476 34748
rect 119532 34802 119924 34804
rect 119532 34750 119870 34802
rect 119922 34750 119924 34802
rect 119532 34748 119924 34750
rect 119308 33966 119310 34018
rect 119362 33966 119364 34018
rect 117404 33070 117406 33122
rect 117458 33070 117460 33122
rect 115612 32498 115668 32508
rect 117404 22932 117460 33070
rect 117852 33236 117908 33246
rect 117852 33122 117908 33180
rect 118412 33236 118468 33246
rect 118412 33142 118468 33180
rect 118748 33236 118804 33246
rect 118748 33142 118804 33180
rect 117852 33070 117854 33122
rect 117906 33070 117908 33122
rect 117852 26908 117908 33070
rect 118748 32452 118804 32462
rect 118748 32358 118804 32396
rect 118972 32452 119028 33964
rect 119308 33954 119364 33966
rect 118972 32386 119028 32396
rect 119084 33572 119140 33582
rect 119084 33348 119140 33516
rect 117628 26852 117908 26908
rect 119084 26908 119140 33292
rect 119308 33122 119364 33134
rect 119308 33070 119310 33122
rect 119362 33070 119364 33122
rect 119308 32676 119364 33070
rect 119196 32620 119364 32676
rect 119196 31780 119252 32620
rect 119196 31714 119252 31724
rect 119308 32452 119364 32462
rect 119532 32452 119588 34748
rect 119868 34738 119924 34748
rect 119644 33234 119700 33246
rect 119644 33182 119646 33234
rect 119698 33182 119700 33234
rect 119644 33124 119700 33182
rect 119644 33058 119700 33068
rect 119980 33012 120036 34862
rect 120092 34130 120148 36204
rect 120204 35700 120260 39200
rect 120428 36708 120484 36718
rect 120428 36370 120484 36652
rect 120428 36318 120430 36370
rect 120482 36318 120484 36370
rect 120428 36306 120484 36318
rect 120652 36596 120708 36606
rect 120204 35644 120372 35700
rect 120092 34078 120094 34130
rect 120146 34078 120148 34130
rect 120092 34066 120148 34078
rect 120204 35474 120260 35486
rect 120204 35422 120206 35474
rect 120258 35422 120260 35474
rect 119756 32956 120036 33012
rect 120092 33124 120148 33134
rect 119756 32786 119812 32956
rect 119756 32734 119758 32786
rect 119810 32734 119812 32786
rect 119756 32722 119812 32734
rect 119308 32450 119588 32452
rect 119308 32398 119310 32450
rect 119362 32398 119588 32450
rect 119308 32396 119588 32398
rect 119084 26852 119252 26908
rect 117628 26180 117684 26852
rect 117628 26114 117684 26124
rect 117404 22866 117460 22876
rect 115276 20962 115332 20972
rect 114268 8372 114548 8428
rect 115724 13412 115780 13422
rect 113596 8148 113652 8158
rect 113596 7700 113652 8092
rect 113484 7698 113652 7700
rect 113484 7646 113598 7698
rect 113650 7646 113652 7698
rect 113484 7644 113652 7646
rect 113372 7250 113428 7262
rect 113372 7198 113374 7250
rect 113426 7198 113428 7250
rect 113372 6690 113428 7198
rect 113372 6638 113374 6690
rect 113426 6638 113428 6690
rect 113372 6626 113428 6638
rect 113484 6580 113540 7644
rect 113596 7634 113652 7644
rect 113372 6132 113428 6142
rect 113484 6132 113540 6524
rect 114156 7362 114212 7374
rect 114156 7310 114158 7362
rect 114210 7310 114212 7362
rect 114156 7250 114212 7310
rect 114156 7198 114158 7250
rect 114210 7198 114212 7250
rect 113372 6130 113540 6132
rect 113372 6078 113374 6130
rect 113426 6078 113540 6130
rect 113372 6076 113540 6078
rect 114044 6466 114100 6478
rect 114044 6414 114046 6466
rect 114098 6414 114100 6466
rect 113372 6066 113428 6076
rect 114044 6020 114100 6414
rect 114156 6244 114212 7198
rect 114156 6178 114212 6188
rect 114044 5954 114100 5964
rect 114268 6020 114324 8372
rect 115164 8148 115220 8158
rect 114380 6804 114436 6814
rect 114380 6710 114436 6748
rect 115164 6690 115220 8092
rect 115724 6804 115780 13356
rect 119196 10052 119252 26852
rect 119308 24612 119364 32396
rect 120092 26180 120148 33068
rect 120204 26908 120260 35422
rect 120316 35252 120372 35644
rect 120316 35186 120372 35196
rect 120540 35476 120596 35486
rect 120540 33460 120596 35420
rect 120652 35138 120708 36540
rect 121100 36036 121156 39200
rect 121548 37156 121604 37166
rect 121436 36260 121492 36270
rect 121436 36166 121492 36204
rect 121100 35980 121492 36036
rect 121100 35588 121156 35598
rect 121100 35494 121156 35532
rect 120652 35086 120654 35138
rect 120706 35086 120708 35138
rect 120652 35074 120708 35086
rect 121100 35252 121156 35262
rect 120988 34690 121044 34702
rect 120988 34638 120990 34690
rect 121042 34638 121044 34690
rect 120652 33460 120708 33470
rect 120540 33458 120708 33460
rect 120540 33406 120654 33458
rect 120706 33406 120708 33458
rect 120540 33404 120708 33406
rect 120652 33394 120708 33404
rect 120204 26852 120484 26908
rect 120092 26114 120148 26124
rect 119308 24546 119364 24556
rect 120428 20188 120484 26852
rect 120988 26068 121044 34638
rect 121100 33458 121156 35196
rect 121436 34242 121492 35980
rect 121548 35026 121604 37100
rect 121772 36372 121828 36382
rect 121996 36372 122052 39200
rect 122220 36708 122276 36718
rect 122220 36594 122276 36652
rect 122220 36542 122222 36594
rect 122274 36542 122276 36594
rect 122220 36530 122276 36542
rect 121772 36370 121940 36372
rect 121772 36318 121774 36370
rect 121826 36318 121940 36370
rect 121772 36316 121940 36318
rect 121772 36306 121828 36316
rect 121548 34974 121550 35026
rect 121602 34974 121604 35026
rect 121548 34962 121604 34974
rect 121436 34190 121438 34242
rect 121490 34190 121492 34242
rect 121436 34178 121492 34190
rect 121100 33406 121102 33458
rect 121154 33406 121156 33458
rect 121100 33394 121156 33406
rect 121772 33570 121828 33582
rect 121772 33518 121774 33570
rect 121826 33518 121828 33570
rect 120988 26002 121044 26012
rect 121772 33122 121828 33518
rect 121772 33070 121774 33122
rect 121826 33070 121828 33122
rect 121772 22596 121828 33070
rect 121884 33124 121940 36316
rect 121996 36306 122052 36316
rect 122108 35810 122164 35822
rect 122108 35758 122110 35810
rect 122162 35758 122164 35810
rect 122108 35252 122164 35758
rect 122108 35186 122164 35196
rect 122556 35812 122612 35822
rect 122332 34804 122388 34814
rect 122220 34802 122388 34804
rect 122220 34750 122334 34802
rect 122386 34750 122388 34802
rect 122220 34748 122388 34750
rect 122220 33570 122276 34748
rect 122332 34738 122388 34748
rect 122556 34130 122612 35756
rect 122668 35140 122724 35150
rect 122668 34914 122724 35084
rect 122668 34862 122670 34914
rect 122722 34862 122724 34914
rect 122668 34850 122724 34862
rect 122556 34078 122558 34130
rect 122610 34078 122612 34130
rect 122556 34066 122612 34078
rect 122892 34020 122948 39200
rect 123340 36596 123396 36606
rect 123340 36502 123396 36540
rect 123116 35812 123172 35822
rect 123788 35812 123844 39200
rect 124684 37156 124740 39200
rect 125356 38612 125412 38622
rect 124684 37100 125188 37156
rect 124348 36372 124404 36382
rect 124348 36278 124404 36316
rect 125020 35812 125076 35822
rect 123788 35810 125076 35812
rect 123788 35758 125022 35810
rect 125074 35758 125076 35810
rect 123788 35756 125076 35758
rect 123116 35718 123172 35756
rect 123452 35698 123508 35710
rect 123452 35646 123454 35698
rect 123506 35646 123508 35698
rect 123452 35588 123508 35646
rect 124012 35588 124068 35598
rect 123452 35522 123508 35532
rect 123564 35586 124068 35588
rect 123564 35534 124014 35586
rect 124066 35534 124068 35586
rect 123564 35532 124068 35534
rect 122892 33954 122948 33964
rect 123004 35364 123060 35374
rect 123564 35364 123620 35532
rect 124012 35522 124068 35532
rect 124796 35588 124852 35598
rect 123004 34132 123060 35308
rect 123116 35308 123620 35364
rect 123116 35138 123172 35308
rect 123116 35086 123118 35138
rect 123170 35086 123172 35138
rect 123116 35074 123172 35086
rect 124012 35140 124068 35150
rect 124012 35026 124068 35084
rect 124012 34974 124014 35026
rect 124066 34974 124068 35026
rect 124012 34916 124068 34974
rect 124012 34850 124068 34860
rect 123452 34690 123508 34702
rect 123452 34638 123454 34690
rect 123506 34638 123508 34690
rect 123116 34132 123172 34142
rect 123004 34130 123172 34132
rect 123004 34078 123118 34130
rect 123170 34078 123172 34130
rect 123004 34076 123172 34078
rect 122220 33518 122222 33570
rect 122274 33518 122276 33570
rect 122220 33506 122276 33518
rect 122892 33460 122948 33470
rect 123004 33460 123060 34076
rect 123116 34066 123172 34076
rect 122892 33458 123060 33460
rect 122892 33406 122894 33458
rect 122946 33406 123060 33458
rect 122892 33404 123060 33406
rect 122892 33394 122948 33404
rect 122108 33124 122164 33134
rect 121884 33122 122164 33124
rect 121884 33070 122110 33122
rect 122162 33070 122164 33122
rect 121884 33068 122164 33070
rect 121772 22530 121828 22540
rect 120428 20132 120596 20188
rect 119196 9986 119252 9996
rect 115724 6738 115780 6748
rect 115836 8708 115892 8718
rect 115164 6638 115166 6690
rect 115218 6638 115220 6690
rect 115052 6580 115108 6590
rect 115052 6486 115108 6524
rect 115164 6356 115220 6638
rect 114940 6300 115220 6356
rect 115724 6580 115780 6590
rect 114380 6020 114436 6030
rect 114268 5964 114380 6020
rect 114268 5906 114324 5964
rect 114380 5954 114436 5964
rect 114268 5854 114270 5906
rect 114322 5854 114324 5906
rect 114268 5842 114324 5854
rect 114940 5906 114996 6300
rect 114940 5854 114942 5906
rect 114994 5854 114996 5906
rect 114940 5842 114996 5854
rect 115052 6018 115108 6030
rect 115052 5966 115054 6018
rect 115106 5966 115108 6018
rect 113932 5684 113988 5694
rect 113932 5590 113988 5628
rect 115052 5236 115108 5966
rect 115612 6020 115668 6030
rect 115612 5926 115668 5964
rect 115724 5796 115780 6524
rect 115500 5740 115780 5796
rect 115500 5346 115556 5740
rect 115500 5294 115502 5346
rect 115554 5294 115556 5346
rect 115500 5282 115556 5294
rect 115052 5170 115108 5180
rect 113596 4900 113652 4910
rect 113596 4338 113652 4844
rect 114940 4900 114996 4910
rect 115836 4900 115892 8652
rect 119196 8260 119252 8270
rect 119196 8166 119252 8204
rect 120540 8260 120596 20132
rect 122108 15988 122164 33068
rect 122108 15922 122164 15932
rect 122444 26068 122500 26078
rect 120540 8166 120596 8204
rect 120988 10052 121044 10062
rect 118300 8148 118356 8158
rect 118300 8054 118356 8092
rect 119420 8148 119476 8158
rect 119420 8054 119476 8092
rect 119868 8146 119924 8158
rect 119868 8094 119870 8146
rect 119922 8094 119924 8146
rect 118860 8036 118916 8046
rect 118860 8034 119252 8036
rect 118860 7982 118862 8034
rect 118914 7982 119252 8034
rect 118860 7980 119252 7982
rect 118860 7970 118916 7980
rect 118076 7588 118132 7598
rect 117740 7586 118132 7588
rect 117740 7534 118078 7586
rect 118130 7534 118132 7586
rect 117740 7532 118132 7534
rect 115948 7362 116004 7374
rect 115948 7310 115950 7362
rect 116002 7310 116004 7362
rect 115948 5348 116004 7310
rect 116732 7362 116788 7374
rect 116732 7310 116734 7362
rect 116786 7310 116788 7362
rect 116508 6916 116564 6926
rect 116284 6580 116340 6590
rect 116284 6466 116340 6524
rect 116284 6414 116286 6466
rect 116338 6414 116340 6466
rect 116284 6356 116340 6414
rect 116284 6290 116340 6300
rect 116508 5906 116564 6860
rect 116732 6692 116788 7310
rect 117516 7364 117572 7374
rect 117516 7270 117572 7308
rect 116732 6468 116788 6636
rect 117628 6690 117684 6702
rect 117628 6638 117630 6690
rect 117682 6638 117684 6690
rect 117180 6468 117236 6478
rect 117628 6468 117684 6638
rect 116732 6466 117684 6468
rect 116732 6414 117182 6466
rect 117234 6414 117684 6466
rect 116732 6412 117684 6414
rect 117068 6132 117124 6142
rect 116508 5854 116510 5906
rect 116562 5854 116564 5906
rect 116508 5842 116564 5854
rect 116844 6130 117124 6132
rect 116844 6078 117070 6130
rect 117122 6078 117124 6130
rect 116844 6076 117124 6078
rect 116172 5796 116228 5806
rect 116172 5702 116228 5740
rect 116844 5460 116900 6076
rect 117068 6066 117124 6076
rect 116284 5404 116900 5460
rect 115948 5282 116004 5292
rect 116172 5348 116228 5358
rect 116172 5234 116228 5292
rect 116284 5346 116340 5404
rect 116284 5294 116286 5346
rect 116338 5294 116340 5346
rect 116284 5282 116340 5294
rect 116172 5182 116174 5234
rect 116226 5182 116228 5234
rect 116172 5170 116228 5182
rect 116732 5236 116788 5246
rect 114940 4898 115444 4900
rect 114940 4846 114942 4898
rect 114994 4846 115444 4898
rect 114940 4844 115444 4846
rect 114940 4834 114996 4844
rect 113596 4286 113598 4338
rect 113650 4286 113652 4338
rect 113596 4274 113652 4286
rect 115388 3780 115444 4844
rect 115836 4834 115892 4844
rect 116172 4562 116228 4574
rect 116172 4510 116174 4562
rect 116226 4510 116228 4562
rect 115948 4228 116004 4238
rect 115500 3780 115556 3790
rect 115388 3778 115556 3780
rect 115388 3726 115502 3778
rect 115554 3726 115556 3778
rect 115388 3724 115556 3726
rect 115500 3714 115556 3724
rect 113260 3614 113262 3666
rect 113314 3614 113316 3666
rect 113260 3602 113316 3614
rect 114604 3668 114660 3678
rect 112588 3502 112590 3554
rect 112642 3502 112644 3554
rect 112588 3490 112644 3502
rect 112364 3390 112366 3442
rect 112418 3390 112420 3442
rect 112364 3378 112420 3390
rect 113260 3444 113316 3454
rect 111916 924 112196 980
rect 111916 800 111972 924
rect 113260 800 113316 3388
rect 114604 3444 114660 3612
rect 114604 3312 114660 3388
rect 115612 3444 115668 3454
rect 115612 3350 115668 3388
rect 115948 800 116004 4172
rect 116172 3778 116228 4510
rect 116732 4562 116788 5180
rect 117180 5124 117236 6412
rect 117180 5030 117236 5068
rect 117628 5124 117684 5134
rect 117740 5124 117796 7532
rect 118076 7522 118132 7532
rect 118412 7476 118468 7486
rect 119084 7476 119140 7486
rect 118412 7474 119140 7476
rect 118412 7422 118414 7474
rect 118466 7422 119086 7474
rect 119138 7422 119140 7474
rect 118412 7420 119140 7422
rect 118412 7410 118468 7420
rect 119084 7410 119140 7420
rect 118300 6692 118356 6702
rect 118300 6690 119028 6692
rect 118300 6638 118302 6690
rect 118354 6638 119028 6690
rect 118300 6636 119028 6638
rect 118300 6626 118356 6636
rect 117628 5122 117796 5124
rect 117628 5070 117630 5122
rect 117682 5070 117796 5122
rect 117628 5068 117796 5070
rect 117628 5058 117684 5068
rect 116732 4510 116734 4562
rect 116786 4510 116788 4562
rect 116732 4498 116788 4510
rect 117180 4900 117236 4910
rect 116172 3726 116174 3778
rect 116226 3726 116228 3778
rect 116172 3714 116228 3726
rect 117180 3666 117236 4844
rect 118972 4562 119028 6636
rect 119196 6132 119252 7980
rect 119644 7586 119700 7598
rect 119644 7534 119646 7586
rect 119698 7534 119700 7586
rect 119420 7476 119476 7486
rect 119420 7382 119476 7420
rect 119644 7364 119700 7534
rect 119644 7298 119700 7308
rect 119868 6468 119924 8094
rect 120204 7586 120260 7598
rect 120204 7534 120206 7586
rect 120258 7534 120260 7586
rect 120204 6692 120260 7534
rect 120204 6636 120708 6692
rect 119868 6402 119924 6412
rect 120540 6466 120596 6478
rect 120540 6414 120542 6466
rect 120594 6414 120596 6466
rect 119196 6076 119364 6132
rect 118972 4510 118974 4562
rect 119026 4510 119028 4562
rect 118972 4498 119028 4510
rect 119308 4450 119364 6076
rect 119644 5908 119700 5918
rect 119644 5814 119700 5852
rect 119980 5906 120036 5918
rect 119980 5854 119982 5906
rect 120034 5854 120036 5906
rect 119980 5796 120036 5854
rect 119308 4398 119310 4450
rect 119362 4398 119364 4450
rect 119308 4386 119364 4398
rect 119868 5348 119924 5358
rect 119868 4450 119924 5292
rect 119980 4564 120036 5740
rect 119980 4498 120036 4508
rect 120092 4898 120148 4910
rect 120092 4846 120094 4898
rect 120146 4846 120148 4898
rect 119868 4398 119870 4450
rect 119922 4398 119924 4450
rect 119868 4386 119924 4398
rect 118188 4338 118244 4350
rect 118188 4286 118190 4338
rect 118242 4286 118244 4338
rect 117292 4228 117348 4238
rect 117292 4134 117348 4172
rect 118188 4116 118244 4286
rect 119980 4340 120036 4350
rect 120092 4340 120148 4846
rect 119980 4338 120148 4340
rect 119980 4286 119982 4338
rect 120034 4286 120148 4338
rect 119980 4284 120148 4286
rect 119980 4274 120036 4284
rect 118188 4050 118244 4060
rect 120428 4116 120484 4126
rect 119532 3780 119588 3790
rect 119756 3780 119812 3790
rect 119532 3778 119812 3780
rect 119532 3726 119534 3778
rect 119586 3726 119758 3778
rect 119810 3726 119812 3778
rect 119532 3724 119812 3726
rect 119532 3714 119588 3724
rect 119756 3714 119812 3724
rect 117180 3614 117182 3666
rect 117234 3614 117236 3666
rect 117180 3602 117236 3614
rect 119980 3668 120036 3678
rect 119980 3574 120036 3612
rect 120428 3666 120484 4060
rect 120540 3778 120596 6414
rect 120652 5124 120708 6636
rect 120988 6020 121044 9996
rect 121100 8036 121156 8046
rect 121436 8036 121492 8046
rect 121100 8034 121380 8036
rect 121100 7982 121102 8034
rect 121154 7982 121380 8034
rect 121100 7980 121380 7982
rect 121100 7970 121156 7980
rect 121324 7586 121380 7980
rect 121324 7534 121326 7586
rect 121378 7534 121380 7586
rect 121212 7474 121268 7486
rect 121212 7422 121214 7474
rect 121266 7422 121268 7474
rect 121212 7364 121268 7422
rect 121212 7298 121268 7308
rect 121324 6916 121380 7534
rect 121436 7476 121492 7980
rect 122444 8036 122500 26012
rect 123452 8428 123508 34638
rect 123788 34020 123844 34030
rect 123788 33926 123844 33964
rect 124796 34018 124852 35532
rect 125020 34356 125076 35756
rect 125132 35026 125188 37100
rect 125356 36370 125412 38556
rect 125580 36596 125636 39200
rect 125580 36540 126084 36596
rect 125356 36318 125358 36370
rect 125410 36318 125412 36370
rect 125356 36306 125412 36318
rect 125692 36370 125748 36382
rect 125692 36318 125694 36370
rect 125746 36318 125748 36370
rect 125692 36260 125748 36318
rect 125692 36194 125748 36204
rect 125804 35924 125860 35934
rect 125132 34974 125134 35026
rect 125186 34974 125188 35026
rect 125132 34962 125188 34974
rect 125580 35700 125636 35710
rect 125244 34356 125300 34366
rect 125020 34354 125300 34356
rect 125020 34302 125246 34354
rect 125298 34302 125300 34354
rect 125020 34300 125300 34302
rect 125244 34290 125300 34300
rect 124796 33966 124798 34018
rect 124850 33966 124852 34018
rect 123900 33234 123956 33246
rect 123900 33182 123902 33234
rect 123954 33182 123956 33234
rect 123564 33122 123620 33134
rect 123564 33070 123566 33122
rect 123618 33070 123620 33122
rect 123564 31892 123620 33070
rect 123900 33124 123956 33182
rect 123900 33058 123956 33068
rect 123564 31826 123620 31836
rect 124796 26292 124852 33966
rect 124908 33124 124964 33134
rect 124908 33030 124964 33068
rect 125580 32788 125636 35644
rect 125804 34916 125860 35868
rect 126028 35812 126084 36540
rect 126140 36372 126196 36382
rect 126140 36278 126196 36316
rect 126140 35812 126196 35822
rect 126028 35810 126196 35812
rect 126028 35758 126142 35810
rect 126194 35758 126196 35810
rect 126028 35756 126196 35758
rect 126028 34916 126084 34926
rect 125804 34914 126084 34916
rect 125804 34862 126030 34914
rect 126082 34862 126084 34914
rect 125804 34860 126084 34862
rect 125692 34356 125748 34366
rect 125804 34356 125860 34860
rect 126028 34850 126084 34860
rect 125692 34354 125860 34356
rect 125692 34302 125694 34354
rect 125746 34302 125860 34354
rect 125692 34300 125860 34302
rect 126140 34356 126196 35756
rect 126476 35140 126532 39200
rect 127372 37380 127428 39200
rect 127372 37324 127652 37380
rect 127596 36372 127652 37324
rect 127708 36372 127764 36382
rect 127596 36316 127708 36372
rect 127708 36240 127764 36316
rect 127932 36260 127988 36270
rect 126476 35074 126532 35084
rect 127484 35586 127540 35598
rect 127484 35534 127486 35586
rect 127538 35534 127540 35586
rect 126812 34916 126868 34926
rect 126588 34914 126868 34916
rect 126588 34862 126814 34914
rect 126866 34862 126868 34914
rect 126588 34860 126868 34862
rect 126252 34356 126308 34366
rect 126140 34354 126308 34356
rect 126140 34302 126254 34354
rect 126306 34302 126308 34354
rect 126140 34300 126308 34302
rect 125692 34290 125748 34300
rect 126252 34290 126308 34300
rect 125580 32722 125636 32732
rect 126028 34020 126084 34030
rect 124796 26226 124852 26236
rect 122444 7970 122500 7980
rect 123340 8372 123508 8428
rect 125132 26180 125188 26190
rect 123340 7698 123396 8372
rect 123340 7646 123342 7698
rect 123394 7646 123396 7698
rect 121436 7410 121492 7420
rect 121996 7476 122052 7486
rect 121996 7382 122052 7420
rect 123340 7476 123396 7646
rect 123340 7410 123396 7420
rect 122892 7364 122948 7374
rect 122892 7270 122948 7308
rect 122332 7252 122388 7262
rect 121324 6850 121380 6860
rect 122108 7250 122388 7252
rect 122108 7198 122334 7250
rect 122386 7198 122388 7250
rect 122108 7196 122388 7198
rect 122108 6690 122164 7196
rect 122332 7186 122388 7196
rect 122108 6638 122110 6690
rect 122162 6638 122164 6690
rect 122108 6626 122164 6638
rect 121324 6468 121380 6478
rect 121324 6374 121380 6412
rect 121772 6466 121828 6478
rect 121772 6414 121774 6466
rect 121826 6414 121828 6466
rect 120988 5964 121268 6020
rect 120988 5796 121044 5806
rect 120876 5794 121044 5796
rect 120876 5742 120990 5794
rect 121042 5742 121044 5794
rect 120876 5740 121044 5742
rect 120876 5124 120932 5740
rect 120988 5730 121044 5740
rect 120988 5348 121044 5358
rect 120988 5234 121044 5292
rect 120988 5182 120990 5234
rect 121042 5182 121044 5234
rect 120988 5170 121044 5182
rect 121100 5236 121156 5246
rect 120652 5122 120932 5124
rect 120652 5070 120654 5122
rect 120706 5070 120932 5122
rect 120652 5068 120932 5070
rect 120652 3892 120708 5068
rect 121100 4338 121156 5180
rect 121100 4286 121102 4338
rect 121154 4286 121156 4338
rect 121100 4274 121156 4286
rect 120652 3826 120708 3836
rect 120540 3726 120542 3778
rect 120594 3726 120596 3778
rect 120540 3714 120596 3726
rect 120428 3614 120430 3666
rect 120482 3614 120484 3666
rect 120428 3602 120484 3614
rect 121212 3666 121268 5964
rect 121772 5908 121828 6414
rect 121772 5842 121828 5852
rect 125020 6468 125076 6478
rect 125020 5122 125076 6412
rect 125020 5070 125022 5122
rect 125074 5070 125076 5122
rect 125020 5058 125076 5070
rect 124236 4564 124292 4574
rect 124236 4470 124292 4508
rect 124684 4564 124740 4574
rect 124684 4338 124740 4508
rect 124684 4286 124686 4338
rect 124738 4286 124740 4338
rect 124684 4274 124740 4286
rect 121212 3614 121214 3666
rect 121266 3614 121268 3666
rect 121212 3602 121268 3614
rect 121772 4226 121828 4238
rect 121772 4174 121774 4226
rect 121826 4174 121828 4226
rect 117292 3556 117348 3566
rect 116284 3444 116340 3454
rect 116284 3350 116340 3388
rect 117292 800 117348 3500
rect 118524 3556 118580 3566
rect 118524 3442 118580 3500
rect 118524 3390 118526 3442
rect 118578 3390 118580 3442
rect 118524 3378 118580 3390
rect 119420 3444 119476 3454
rect 119420 3350 119476 3388
rect 120092 3444 120148 3454
rect 120092 2100 120148 3388
rect 121772 3444 121828 4174
rect 125132 3666 125188 26124
rect 126028 25732 126084 33964
rect 126588 34018 126644 34860
rect 126812 34850 126868 34860
rect 127484 34132 127540 35534
rect 127932 35586 127988 36204
rect 127932 35534 127934 35586
rect 127986 35534 127988 35586
rect 127932 35476 127988 35534
rect 127932 35410 127988 35420
rect 127708 35140 127764 35150
rect 127708 35026 127764 35084
rect 127708 34974 127710 35026
rect 127762 34974 127764 35026
rect 127708 34962 127764 34974
rect 127484 34066 127540 34076
rect 127596 34692 127652 34702
rect 126588 33966 126590 34018
rect 126642 33966 126644 34018
rect 126588 33236 126644 33966
rect 126588 33170 126644 33180
rect 127596 30212 127652 34636
rect 128268 33460 128324 39200
rect 129052 36594 129108 36606
rect 129052 36542 129054 36594
rect 129106 36542 129108 36594
rect 128940 36484 128996 36494
rect 128828 34916 128884 34926
rect 128828 34822 128884 34860
rect 128940 34020 128996 36428
rect 129052 35812 129108 36542
rect 129164 35812 129220 39200
rect 130060 37044 130116 39200
rect 129948 36988 130116 37044
rect 129836 36484 129892 36494
rect 129836 36390 129892 36428
rect 129612 36258 129668 36270
rect 129612 36206 129614 36258
rect 129666 36206 129668 36258
rect 129500 35924 129556 35934
rect 129500 35812 129556 35868
rect 129164 35810 129556 35812
rect 129164 35758 129502 35810
rect 129554 35758 129556 35810
rect 129164 35756 129556 35758
rect 129052 35746 129108 35756
rect 129500 35746 129556 35756
rect 128828 34018 128996 34020
rect 128828 33966 128942 34018
rect 128994 33966 128996 34018
rect 128828 33964 128996 33966
rect 128604 33460 128660 33470
rect 128268 33458 128660 33460
rect 128268 33406 128606 33458
rect 128658 33406 128660 33458
rect 128268 33404 128660 33406
rect 128604 33394 128660 33404
rect 127596 30146 127652 30156
rect 126028 25666 126084 25676
rect 126812 27748 126868 27758
rect 126364 11172 126420 11182
rect 126364 7698 126420 11116
rect 126812 9940 126868 27692
rect 128828 12628 128884 33964
rect 128940 33954 128996 33964
rect 129164 35476 129220 35486
rect 129164 20188 129220 35420
rect 129388 34916 129444 34926
rect 129276 34692 129332 34702
rect 129276 34598 129332 34636
rect 129388 34354 129444 34860
rect 129388 34302 129390 34354
rect 129442 34302 129444 34354
rect 129388 34290 129444 34302
rect 129612 33346 129668 36206
rect 129948 35140 130004 36988
rect 130082 36876 130346 36886
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130082 36810 130346 36820
rect 130396 36372 130452 36382
rect 130396 36278 130452 36316
rect 130956 36372 131012 39200
rect 131292 36372 131348 36382
rect 130956 36370 131348 36372
rect 130956 36318 131294 36370
rect 131346 36318 131348 36370
rect 130956 36316 131348 36318
rect 130732 35812 130788 35822
rect 130620 35586 130676 35598
rect 130620 35534 130622 35586
rect 130674 35534 130676 35586
rect 130082 35308 130346 35318
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130082 35242 130346 35252
rect 129948 35084 130228 35140
rect 130060 34916 130116 34926
rect 130060 34822 130116 34860
rect 129948 34802 130004 34814
rect 129948 34750 129950 34802
rect 130002 34750 130004 34802
rect 129948 34692 130004 34750
rect 129948 34626 130004 34636
rect 129948 34020 130004 34030
rect 129948 33926 130004 33964
rect 130172 33908 130228 35084
rect 130508 34916 130564 34926
rect 130508 34130 130564 34860
rect 130620 34804 130676 35534
rect 130732 35138 130788 35756
rect 130732 35086 130734 35138
rect 130786 35086 130788 35138
rect 130732 35074 130788 35086
rect 130620 34748 130788 34804
rect 130508 34078 130510 34130
rect 130562 34078 130564 34130
rect 130508 34066 130564 34078
rect 130620 34242 130676 34254
rect 130620 34190 130622 34242
rect 130674 34190 130676 34242
rect 130620 34020 130676 34190
rect 130620 33954 130676 33964
rect 130732 33908 130788 34748
rect 130172 33852 130564 33908
rect 130082 33740 130346 33750
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130082 33674 130346 33684
rect 130508 33458 130564 33852
rect 130732 33842 130788 33852
rect 130508 33406 130510 33458
rect 130562 33406 130564 33458
rect 130508 33394 130564 33406
rect 129612 33294 129614 33346
rect 129666 33294 129668 33346
rect 129612 33282 129668 33294
rect 130956 32786 131012 36316
rect 131292 36306 131348 36316
rect 131628 36260 131684 36270
rect 131404 35810 131460 35822
rect 131404 35758 131406 35810
rect 131458 35758 131460 35810
rect 130956 32734 130958 32786
rect 131010 32734 131012 32786
rect 130956 32722 131012 32734
rect 131068 34690 131124 34702
rect 131068 34638 131070 34690
rect 131122 34638 131124 34690
rect 131068 32788 131124 34638
rect 131292 34132 131348 34142
rect 131292 34038 131348 34076
rect 131404 33346 131460 35758
rect 131628 35700 131684 36204
rect 131628 35606 131684 35644
rect 131852 35140 131908 39200
rect 132748 36820 132804 39200
rect 132748 36754 132804 36764
rect 132636 36596 132692 36606
rect 132636 36594 132804 36596
rect 132636 36542 132638 36594
rect 132690 36542 132804 36594
rect 132636 36540 132804 36542
rect 132636 36530 132692 36540
rect 132188 35924 132244 35934
rect 132188 35830 132244 35868
rect 131852 35074 131908 35084
rect 132636 35700 132692 35710
rect 131740 34802 131796 34814
rect 131740 34750 131742 34802
rect 131794 34750 131796 34802
rect 131404 33294 131406 33346
rect 131458 33294 131460 33346
rect 131404 33282 131460 33294
rect 131516 34468 131572 34478
rect 131068 32722 131124 32732
rect 131404 32788 131460 32798
rect 131516 32788 131572 34412
rect 131740 34468 131796 34750
rect 132076 34804 132132 34814
rect 132076 34710 132132 34748
rect 131740 34402 131796 34412
rect 132636 34354 132692 35644
rect 132748 35252 132804 36540
rect 133532 36370 133588 36382
rect 133532 36318 133534 36370
rect 133586 36318 133588 36370
rect 133196 36260 133252 36270
rect 133084 36258 133252 36260
rect 133084 36206 133198 36258
rect 133250 36206 133252 36258
rect 133084 36204 133252 36206
rect 132972 35588 133028 35598
rect 132748 35186 132804 35196
rect 132860 35586 133028 35588
rect 132860 35534 132974 35586
rect 133026 35534 133028 35586
rect 132860 35532 133028 35534
rect 132636 34302 132638 34354
rect 132690 34302 132692 34354
rect 132636 34290 132692 34302
rect 132300 34130 132356 34142
rect 132300 34078 132302 34130
rect 132354 34078 132356 34130
rect 131404 32786 131572 32788
rect 131404 32734 131406 32786
rect 131458 32734 131572 32786
rect 131404 32732 131572 32734
rect 131628 33906 131684 33918
rect 131628 33854 131630 33906
rect 131682 33854 131684 33906
rect 131404 32722 131460 32732
rect 130082 32172 130346 32182
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130082 32106 130346 32116
rect 131628 31108 131684 33854
rect 131964 33348 132020 33358
rect 131964 33254 132020 33292
rect 132300 33348 132356 34078
rect 132860 33460 132916 35532
rect 132972 35522 133028 35532
rect 132972 34914 133028 34926
rect 132972 34862 132974 34914
rect 133026 34862 133028 34914
rect 132972 34804 133028 34862
rect 132972 34738 133028 34748
rect 132860 33394 132916 33404
rect 132300 33282 132356 33292
rect 131628 31042 131684 31052
rect 130082 30604 130346 30614
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130082 30538 130346 30548
rect 130082 29036 130346 29046
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130082 28970 130346 28980
rect 133084 28420 133140 36204
rect 133196 36194 133252 36204
rect 133532 36036 133588 36318
rect 133532 34804 133588 35980
rect 133644 35812 133700 39200
rect 133868 36820 133924 36830
rect 133868 35812 133924 36764
rect 134540 36372 134596 39200
rect 135100 36594 135156 36606
rect 135100 36542 135102 36594
rect 135154 36542 135156 36594
rect 135100 36484 135156 36542
rect 135100 36418 135156 36428
rect 134540 36306 134596 36316
rect 135324 36372 135380 36382
rect 133980 36260 134036 36270
rect 133980 36166 134036 36204
rect 133980 35812 134036 35822
rect 133868 35810 134372 35812
rect 133868 35758 133982 35810
rect 134034 35758 134372 35810
rect 133868 35756 134372 35758
rect 133644 35746 133700 35756
rect 133980 35746 134036 35756
rect 133644 35140 133700 35150
rect 133644 35026 133700 35084
rect 133644 34974 133646 35026
rect 133698 34974 133700 35026
rect 133644 34962 133700 34974
rect 133532 34748 133700 34804
rect 133532 34132 133588 34142
rect 133084 28354 133140 28364
rect 133196 34130 133588 34132
rect 133196 34078 133534 34130
rect 133586 34078 133588 34130
rect 133196 34076 133588 34078
rect 133196 33458 133252 34076
rect 133532 34066 133588 34076
rect 133196 33406 133198 33458
rect 133250 33406 133252 33458
rect 130082 27468 130346 27478
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130082 27402 130346 27412
rect 133196 26180 133252 33406
rect 133196 26114 133252 26124
rect 130082 25900 130346 25910
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130082 25834 130346 25844
rect 130082 24332 130346 24342
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130082 24266 130346 24276
rect 130082 22764 130346 22774
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130082 22698 130346 22708
rect 133644 21812 133700 34748
rect 133868 34356 133924 34366
rect 133868 34262 133924 34300
rect 134316 34354 134372 35756
rect 134988 35700 135044 35710
rect 134988 35606 135044 35644
rect 134316 34302 134318 34354
rect 134370 34302 134372 34354
rect 134316 34290 134372 34302
rect 134764 35476 134820 35486
rect 134764 34802 134820 35420
rect 134764 34750 134766 34802
rect 134818 34750 134820 34802
rect 134764 34354 134820 34750
rect 134764 34302 134766 34354
rect 134818 34302 134820 34354
rect 134764 34290 134820 34302
rect 135100 34690 135156 34702
rect 135100 34638 135102 34690
rect 135154 34638 135156 34690
rect 135100 33348 135156 34638
rect 135324 34354 135380 36316
rect 135436 35140 135492 39200
rect 136108 36372 136164 36382
rect 136108 36278 136164 36316
rect 135660 35812 135716 35822
rect 135660 35586 135716 35756
rect 135660 35534 135662 35586
rect 135714 35534 135716 35586
rect 135660 35522 135716 35534
rect 136332 35364 136388 39200
rect 137116 36370 137172 36382
rect 137116 36318 137118 36370
rect 137170 36318 137172 36370
rect 137116 36260 137172 36318
rect 137116 36036 137172 36204
rect 137116 35970 137172 35980
rect 137004 35588 137060 35598
rect 137004 35494 137060 35532
rect 136332 35298 136388 35308
rect 136780 35364 136836 35374
rect 135436 35074 135492 35084
rect 136332 35140 136388 35150
rect 136332 35026 136388 35084
rect 136332 34974 136334 35026
rect 136386 34974 136388 35026
rect 136332 34962 136388 34974
rect 135324 34302 135326 34354
rect 135378 34302 135380 34354
rect 135324 34290 135380 34302
rect 135660 34914 135716 34926
rect 135660 34862 135662 34914
rect 135714 34862 135716 34914
rect 135660 34356 135716 34862
rect 136332 34804 136388 34814
rect 136332 34356 136388 34748
rect 135660 34290 135716 34300
rect 135996 34354 136388 34356
rect 135996 34302 136334 34354
rect 136386 34302 136388 34354
rect 135996 34300 136388 34302
rect 135100 33282 135156 33292
rect 135996 24164 136052 34300
rect 136332 34290 136388 34300
rect 136780 33458 136836 35308
rect 136780 33406 136782 33458
rect 136834 33406 136836 33458
rect 136780 33394 136836 33406
rect 137004 34244 137060 34254
rect 137004 26852 137060 34188
rect 137228 33460 137284 39200
rect 138124 36372 138180 39200
rect 139020 36932 139076 39200
rect 139916 36932 139972 39200
rect 139020 36876 139188 36932
rect 139916 36876 140308 36932
rect 138124 36306 138180 36316
rect 139020 36594 139076 36606
rect 139020 36542 139022 36594
rect 139074 36542 139076 36594
rect 137452 36258 137508 36270
rect 137452 36206 137454 36258
rect 137506 36206 137508 36258
rect 137340 34692 137396 34702
rect 137340 34598 137396 34636
rect 137340 34468 137396 34478
rect 137340 34018 137396 34412
rect 137452 34132 137508 36206
rect 138012 36260 138068 36270
rect 138012 36166 138068 36204
rect 139020 36148 139076 36542
rect 139020 36082 139076 36092
rect 138012 35810 138068 35822
rect 138012 35758 138014 35810
rect 138066 35758 138068 35810
rect 138012 35364 138068 35758
rect 138012 35298 138068 35308
rect 139020 35698 139076 35710
rect 139020 35646 139022 35698
rect 139074 35646 139076 35698
rect 138796 35252 138852 35262
rect 138796 35138 138852 35196
rect 138796 35086 138798 35138
rect 138850 35086 138852 35138
rect 138796 35074 138852 35086
rect 139020 34916 139076 35646
rect 139132 35140 139188 36876
rect 140028 36372 140084 36382
rect 139356 35810 139412 35822
rect 139356 35758 139358 35810
rect 139410 35758 139412 35810
rect 139356 35252 139412 35758
rect 139356 35186 139412 35196
rect 139132 35074 139188 35084
rect 140028 35028 140084 36316
rect 140252 35810 140308 36876
rect 140252 35758 140254 35810
rect 140306 35758 140308 35810
rect 140140 35028 140196 35038
rect 140028 35026 140196 35028
rect 140028 34974 140142 35026
rect 140194 34974 140196 35026
rect 140028 34972 140196 34974
rect 140140 34962 140196 34972
rect 139020 34860 139300 34916
rect 138012 34804 138068 34814
rect 138012 34710 138068 34748
rect 138572 34804 138628 34814
rect 138348 34244 138404 34254
rect 138348 34150 138404 34188
rect 137452 34066 137508 34076
rect 138572 34130 138628 34748
rect 139132 34692 139188 34702
rect 138572 34078 138574 34130
rect 138626 34078 138628 34130
rect 138572 34066 138628 34078
rect 138684 34690 139188 34692
rect 138684 34638 139134 34690
rect 139186 34638 139188 34690
rect 138684 34636 139188 34638
rect 137340 33966 137342 34018
rect 137394 33966 137396 34018
rect 137340 33908 137396 33966
rect 137340 33842 137396 33852
rect 137228 33394 137284 33404
rect 138124 33460 138180 33470
rect 138124 33366 138180 33404
rect 137452 33348 137508 33358
rect 137452 33254 137508 33292
rect 138684 31948 138740 34636
rect 139132 34626 139188 34636
rect 139020 34468 139076 34478
rect 139020 34130 139076 34412
rect 139020 34078 139022 34130
rect 139074 34078 139076 34130
rect 139020 34066 139076 34078
rect 139244 33460 139300 34860
rect 139692 34804 139748 34814
rect 139692 34710 139748 34748
rect 140028 34132 140084 34142
rect 140028 34038 140084 34076
rect 137004 26786 137060 26796
rect 138348 31892 138740 31948
rect 138796 33124 138852 33134
rect 135996 24098 136052 24108
rect 133644 21746 133700 21756
rect 134428 21812 134484 21822
rect 130082 21196 130346 21206
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130082 21130 130346 21140
rect 128828 12562 128884 12572
rect 129052 20132 129220 20188
rect 126812 9874 126868 9884
rect 128716 9940 128772 9950
rect 128716 9846 128772 9884
rect 128268 9154 128324 9166
rect 128268 9102 128270 9154
rect 128322 9102 128324 9154
rect 128044 9044 128100 9054
rect 128044 8950 128100 8988
rect 128268 8428 128324 9102
rect 128268 8372 128436 8428
rect 127372 8148 127428 8158
rect 127036 8146 127428 8148
rect 127036 8094 127374 8146
rect 127426 8094 127428 8146
rect 127036 8092 127428 8094
rect 126812 8036 126868 8046
rect 126812 8034 126980 8036
rect 126812 7982 126814 8034
rect 126866 7982 126980 8034
rect 126812 7980 126980 7982
rect 126812 7970 126868 7980
rect 126364 7646 126366 7698
rect 126418 7646 126420 7698
rect 126028 7588 126084 7598
rect 126028 7494 126084 7532
rect 126364 6916 126420 7646
rect 126588 6916 126644 6926
rect 126364 6914 126644 6916
rect 126364 6862 126590 6914
rect 126642 6862 126644 6914
rect 126364 6860 126644 6862
rect 126588 6850 126644 6860
rect 126924 6468 126980 7980
rect 127036 7698 127092 8092
rect 127372 8082 127428 8092
rect 127036 7646 127038 7698
rect 127090 7646 127092 7698
rect 127036 7634 127092 7646
rect 127708 8034 127764 8046
rect 127708 7982 127710 8034
rect 127762 7982 127764 8034
rect 127036 7476 127092 7486
rect 127036 6690 127092 7420
rect 127372 7250 127428 7262
rect 127372 7198 127374 7250
rect 127426 7198 127428 7250
rect 127372 6914 127428 7198
rect 127372 6862 127374 6914
rect 127426 6862 127428 6914
rect 127372 6850 127428 6862
rect 127708 6916 127764 7982
rect 128156 8034 128212 8046
rect 128156 7982 128158 8034
rect 128210 7982 128212 8034
rect 128156 7812 128212 7982
rect 128156 7746 128212 7756
rect 128044 7700 128100 7710
rect 128044 7586 128100 7644
rect 128044 7534 128046 7586
rect 128098 7534 128100 7586
rect 128044 7522 128100 7534
rect 128156 7476 128212 7486
rect 128156 7382 128212 7420
rect 127708 6860 128324 6916
rect 127036 6638 127038 6690
rect 127090 6638 127092 6690
rect 127036 6626 127092 6638
rect 128044 6690 128100 6702
rect 128044 6638 128046 6690
rect 128098 6638 128100 6690
rect 126476 6356 126532 6366
rect 126476 6130 126532 6300
rect 126476 6078 126478 6130
rect 126530 6078 126532 6130
rect 126476 6066 126532 6078
rect 125692 5234 125748 5246
rect 125692 5182 125694 5234
rect 125746 5182 125748 5234
rect 125356 4340 125412 4350
rect 125356 4246 125412 4284
rect 125132 3614 125134 3666
rect 125186 3614 125188 3666
rect 125132 3602 125188 3614
rect 123228 3556 123284 3566
rect 123228 3462 123284 3500
rect 121772 3378 121828 3388
rect 122108 3444 122164 3454
rect 119980 2044 120148 2100
rect 119980 800 120036 2044
rect 121324 924 121604 980
rect 121324 800 121380 924
rect 69244 700 69636 756
rect 70224 0 70336 800
rect 71568 0 71680 800
rect 72912 0 73024 800
rect 74256 0 74368 800
rect 75600 0 75712 800
rect 76944 0 77056 800
rect 78288 0 78400 800
rect 79632 0 79744 800
rect 80976 0 81088 800
rect 82320 0 82432 800
rect 83664 0 83776 800
rect 85008 0 85120 800
rect 86352 0 86464 800
rect 87696 0 87808 800
rect 89040 0 89152 800
rect 90384 0 90496 800
rect 91728 0 91840 800
rect 93072 0 93184 800
rect 94416 0 94528 800
rect 95760 0 95872 800
rect 97104 0 97216 800
rect 98448 0 98560 800
rect 99792 0 99904 800
rect 101136 0 101248 800
rect 102480 0 102592 800
rect 103824 0 103936 800
rect 105168 0 105280 800
rect 106512 0 106624 800
rect 107856 0 107968 800
rect 109200 0 109312 800
rect 110544 0 110656 800
rect 111888 0 112000 800
rect 113232 0 113344 800
rect 114576 0 114688 800
rect 115920 0 116032 800
rect 117264 0 117376 800
rect 118608 0 118720 800
rect 119952 0 120064 800
rect 121296 0 121408 800
rect 121548 756 121604 924
rect 122108 756 122164 3388
rect 123676 3444 123732 3454
rect 123676 3350 123732 3388
rect 124012 3444 124068 3454
rect 124012 800 124068 3388
rect 125692 3444 125748 5182
rect 126924 5234 126980 6412
rect 127372 6468 127428 6478
rect 127372 6374 127428 6412
rect 128044 6468 128100 6638
rect 127148 6356 127204 6366
rect 127148 5906 127204 6300
rect 127148 5854 127150 5906
rect 127202 5854 127204 5906
rect 127148 5842 127204 5854
rect 126924 5182 126926 5234
rect 126978 5182 126980 5234
rect 126924 5124 126980 5182
rect 126924 5058 126980 5068
rect 127372 5124 127428 5134
rect 127820 5124 127876 5134
rect 127372 5122 127876 5124
rect 127372 5070 127374 5122
rect 127426 5070 127822 5122
rect 127874 5070 127876 5122
rect 127372 5068 127876 5070
rect 127372 4564 127428 5068
rect 127820 5058 127876 5068
rect 127372 4498 127428 4508
rect 127820 4562 127876 4574
rect 127820 4510 127822 4562
rect 127874 4510 127876 4562
rect 127820 3780 127876 4510
rect 127820 3714 127876 3724
rect 128044 3666 128100 6412
rect 128044 3614 128046 3666
rect 128098 3614 128100 3666
rect 128044 3602 128100 3614
rect 128156 5794 128212 5806
rect 128156 5742 128158 5794
rect 128210 5742 128212 5794
rect 126028 3444 126084 3454
rect 125692 3378 125748 3388
rect 125804 3388 126028 3444
rect 125804 1764 125860 3388
rect 126028 3378 126084 3388
rect 126364 3444 126420 3454
rect 126364 3350 126420 3388
rect 127148 3444 127204 3454
rect 127148 3350 127204 3388
rect 128156 2884 128212 5742
rect 128268 5124 128324 6860
rect 128380 6690 128436 8372
rect 128940 8036 128996 8046
rect 128940 7942 128996 7980
rect 128940 7252 128996 7262
rect 128940 7158 128996 7196
rect 128380 6638 128382 6690
rect 128434 6638 128436 6690
rect 128380 6626 128436 6638
rect 128492 5348 128548 5358
rect 128380 5124 128436 5134
rect 128268 5122 128436 5124
rect 128268 5070 128382 5122
rect 128434 5070 128436 5122
rect 128268 5068 128436 5070
rect 128380 5058 128436 5068
rect 128380 4564 128436 4574
rect 128492 4564 128548 5292
rect 128380 4562 128548 4564
rect 128380 4510 128382 4562
rect 128434 4510 128548 4562
rect 128380 4508 128548 4510
rect 128604 4900 128660 4910
rect 128380 4498 128436 4508
rect 128604 4340 128660 4844
rect 128492 3668 128548 3678
rect 128604 3668 128660 4284
rect 128492 3666 128660 3668
rect 128492 3614 128494 3666
rect 128546 3614 128660 3666
rect 128492 3612 128660 3614
rect 129052 3666 129108 20132
rect 130082 19628 130346 19638
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130082 19562 130346 19572
rect 130082 18060 130346 18070
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130082 17994 130346 18004
rect 130082 16492 130346 16502
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130082 16426 130346 16436
rect 130082 14924 130346 14934
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130082 14858 130346 14868
rect 130082 13356 130346 13366
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130082 13290 130346 13300
rect 130082 11788 130346 11798
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130082 11722 130346 11732
rect 130082 10220 130346 10230
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130082 10154 130346 10164
rect 129500 9940 129556 9950
rect 129276 9602 129332 9614
rect 129276 9550 129278 9602
rect 129330 9550 129332 9602
rect 129164 9044 129220 9054
rect 129164 8950 129220 8988
rect 129276 8428 129332 9550
rect 129500 9042 129556 9884
rect 130172 9156 130228 9166
rect 130172 9062 130228 9100
rect 131292 9156 131348 9166
rect 129500 8990 129502 9042
rect 129554 8990 129556 9042
rect 129500 8978 129556 8990
rect 130284 9044 130340 9054
rect 130844 9044 130900 9054
rect 130284 9042 130900 9044
rect 130284 8990 130286 9042
rect 130338 8990 130846 9042
rect 130898 8990 130900 9042
rect 130284 8988 130900 8990
rect 130284 8978 130340 8988
rect 130082 8652 130346 8662
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130082 8586 130346 8596
rect 129164 8372 129332 8428
rect 129164 6468 129220 8372
rect 129724 7588 129780 7598
rect 129724 7494 129780 7532
rect 130844 7476 130900 8988
rect 131292 8428 131348 9100
rect 131292 8372 131572 8428
rect 131292 8258 131348 8270
rect 131292 8206 131294 8258
rect 131346 8206 131348 8258
rect 131292 7924 131348 8206
rect 131292 7858 131348 7868
rect 130844 7410 130900 7420
rect 129164 5906 129220 6412
rect 129164 5854 129166 5906
rect 129218 5854 129220 5906
rect 129164 4338 129220 5854
rect 129612 7364 129668 7374
rect 129612 5906 129668 7308
rect 130082 7084 130346 7094
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130082 7018 130346 7028
rect 130956 6580 131012 6590
rect 130956 6466 131012 6524
rect 130956 6414 130958 6466
rect 131010 6414 131012 6466
rect 130956 6402 131012 6414
rect 131516 6466 131572 8372
rect 131852 8258 131908 8270
rect 131852 8206 131854 8258
rect 131906 8206 131908 8258
rect 131516 6414 131518 6466
rect 131570 6414 131572 6466
rect 131516 6356 131572 6414
rect 131516 6290 131572 6300
rect 131628 7700 131684 7710
rect 131628 6804 131684 7644
rect 129612 5854 129614 5906
rect 129666 5854 129668 5906
rect 129612 5842 129668 5854
rect 130082 5516 130346 5526
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130082 5450 130346 5460
rect 131516 5348 131572 5358
rect 131628 5348 131684 6748
rect 131852 6468 131908 8206
rect 132300 8036 132356 8046
rect 132300 7942 132356 7980
rect 132860 8034 132916 8046
rect 132860 7982 132862 8034
rect 132914 7982 132916 8034
rect 132860 7924 132916 7982
rect 132860 7858 132916 7868
rect 133644 7588 133700 7598
rect 132076 7474 132132 7486
rect 132076 7422 132078 7474
rect 132130 7422 132132 7474
rect 132076 7140 132132 7422
rect 132076 7074 132132 7084
rect 132636 7474 132692 7486
rect 132636 7422 132638 7474
rect 132690 7422 132692 7474
rect 131964 6580 132020 6590
rect 131964 6486 132020 6524
rect 132076 6580 132132 6590
rect 132076 6578 132244 6580
rect 132076 6526 132078 6578
rect 132130 6526 132244 6578
rect 132076 6524 132244 6526
rect 132076 6514 132132 6524
rect 131852 6402 131908 6412
rect 132076 6132 132132 6142
rect 132076 6038 132132 6076
rect 132188 6020 132244 6524
rect 132636 6468 132692 7422
rect 133084 7362 133140 7374
rect 133084 7310 133086 7362
rect 133138 7310 133140 7362
rect 133084 7140 133140 7310
rect 133532 7364 133588 7374
rect 133532 7270 133588 7308
rect 133084 7074 133140 7084
rect 133644 6690 133700 7532
rect 133644 6638 133646 6690
rect 133698 6638 133700 6690
rect 133644 6626 133700 6638
rect 133084 6578 133140 6590
rect 133084 6526 133086 6578
rect 133138 6526 133140 6578
rect 132636 6402 132692 6412
rect 132972 6466 133028 6478
rect 132972 6414 132974 6466
rect 133026 6414 133028 6466
rect 131516 5346 131684 5348
rect 131516 5294 131518 5346
rect 131570 5294 131684 5346
rect 131516 5292 131684 5294
rect 131852 5684 131908 5694
rect 131516 5282 131572 5292
rect 130956 5124 131012 5134
rect 130956 4898 131012 5068
rect 130956 4846 130958 4898
rect 131010 4846 131012 4898
rect 130956 4834 131012 4846
rect 131852 4562 131908 5628
rect 132076 5236 132132 5246
rect 132188 5236 132244 5964
rect 132860 6244 132916 6254
rect 132076 5234 132244 5236
rect 132076 5182 132078 5234
rect 132130 5182 132244 5234
rect 132076 5180 132244 5182
rect 132636 5682 132692 5694
rect 132636 5630 132638 5682
rect 132690 5630 132692 5682
rect 132076 5170 132132 5180
rect 131964 5124 132020 5134
rect 131964 5030 132020 5068
rect 131852 4510 131854 4562
rect 131906 4510 131908 4562
rect 131852 4498 131908 4510
rect 132188 4564 132244 4574
rect 129164 4286 129166 4338
rect 129218 4286 129220 4338
rect 129164 4274 129220 4286
rect 129612 4340 129668 4350
rect 129612 4246 129668 4284
rect 132076 4228 132132 4238
rect 130082 3948 130346 3958
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130082 3882 130346 3892
rect 131516 3780 131572 3790
rect 131516 3686 131572 3724
rect 129052 3614 129054 3666
rect 129106 3614 129108 3666
rect 128492 3602 128548 3612
rect 129052 3602 129108 3614
rect 131628 3668 131684 3678
rect 131628 3574 131684 3612
rect 125356 1708 125860 1764
rect 128044 2828 128212 2884
rect 129388 3556 129444 3566
rect 125356 800 125412 1708
rect 128044 800 128100 2828
rect 129388 800 129444 3500
rect 130284 3556 130340 3566
rect 130284 3442 130340 3500
rect 130284 3390 130286 3442
rect 130338 3390 130340 3442
rect 130284 3378 130340 3390
rect 132076 800 132132 4172
rect 132188 3668 132244 4508
rect 132636 4452 132692 5630
rect 132860 5460 132916 6188
rect 132972 6132 133028 6414
rect 132972 6066 133028 6076
rect 133084 6020 133140 6526
rect 133084 5926 133140 5964
rect 133756 6578 133812 6590
rect 133756 6526 133758 6578
rect 133810 6526 133812 6578
rect 132860 5346 132916 5404
rect 132860 5294 132862 5346
rect 132914 5294 132916 5346
rect 132860 5282 132916 5294
rect 133308 5906 133364 5918
rect 133308 5854 133310 5906
rect 133362 5854 133364 5906
rect 132636 4386 132692 4396
rect 133308 5012 133364 5854
rect 133196 4228 133252 4238
rect 133196 4134 133252 4172
rect 132636 4116 132692 4126
rect 132636 4022 132692 4060
rect 133308 4004 133364 4956
rect 133308 3938 133364 3948
rect 133420 4898 133476 4910
rect 133420 4846 133422 4898
rect 133474 4846 133476 4898
rect 132300 3780 132356 3790
rect 132300 3686 132356 3724
rect 133420 3780 133476 4846
rect 133756 4564 133812 6526
rect 134204 6468 134260 6478
rect 134092 6020 134148 6030
rect 134092 5926 134148 5964
rect 133980 5684 134036 5694
rect 133980 5590 134036 5628
rect 134204 5124 134260 6412
rect 134204 5058 134260 5068
rect 134316 5796 134372 5806
rect 133756 4498 133812 4508
rect 134316 4338 134372 5740
rect 134316 4286 134318 4338
rect 134370 4286 134372 4338
rect 134316 4116 134372 4286
rect 134316 4050 134372 4060
rect 133420 3714 133476 3724
rect 132188 3536 132244 3612
rect 134316 3668 134372 3678
rect 134428 3668 134484 21756
rect 134764 8036 134820 8046
rect 134540 5794 134596 5806
rect 134540 5742 134542 5794
rect 134594 5742 134596 5794
rect 134540 5012 134596 5742
rect 134540 4946 134596 4956
rect 134316 3666 134484 3668
rect 134316 3614 134318 3666
rect 134370 3614 134484 3666
rect 134316 3612 134484 3614
rect 134316 3602 134372 3612
rect 133308 3444 133364 3454
rect 134764 3444 134820 7980
rect 137900 6020 137956 6030
rect 134988 5796 135044 5806
rect 135436 5796 135492 5806
rect 134988 5702 135044 5740
rect 135212 5794 135492 5796
rect 135212 5742 135438 5794
rect 135490 5742 135492 5794
rect 135212 5740 135492 5742
rect 135212 5012 135268 5740
rect 135436 5730 135492 5740
rect 137452 5794 137508 5806
rect 137452 5742 137454 5794
rect 137506 5742 137508 5794
rect 137340 5684 137396 5694
rect 136220 5236 136276 5246
rect 134876 4564 134932 4574
rect 134932 4508 135156 4564
rect 134876 4470 134932 4508
rect 135100 3668 135156 4508
rect 135212 4450 135268 4956
rect 135884 5122 135940 5134
rect 135884 5070 135886 5122
rect 135938 5070 135940 5122
rect 135884 4562 135940 5070
rect 135884 4510 135886 4562
rect 135938 4510 135940 4562
rect 135884 4498 135940 4510
rect 135212 4398 135214 4450
rect 135266 4398 135268 4450
rect 135212 4386 135268 4398
rect 136220 4450 136276 5180
rect 136332 5124 136388 5134
rect 136332 5030 136388 5068
rect 137340 5010 137396 5628
rect 137340 4958 137342 5010
rect 137394 4958 137396 5010
rect 137340 4946 137396 4958
rect 137004 4900 137060 4910
rect 137004 4806 137060 4844
rect 136220 4398 136222 4450
rect 136274 4398 136276 4450
rect 136220 4386 136276 4398
rect 137340 4452 137396 4462
rect 136892 4340 136948 4350
rect 136892 4246 136948 4284
rect 135212 3668 135268 3678
rect 135100 3666 135268 3668
rect 135100 3614 135214 3666
rect 135266 3614 135268 3666
rect 135100 3612 135268 3614
rect 135212 3602 135268 3612
rect 137340 3668 137396 4396
rect 135660 3556 135716 3566
rect 135660 3462 135716 3500
rect 137340 3554 137396 3612
rect 137340 3502 137342 3554
rect 137394 3502 137396 3554
rect 137340 3490 137396 3502
rect 137452 4452 137508 5742
rect 137900 5348 137956 5964
rect 137900 5282 137956 5292
rect 138348 5346 138404 31892
rect 138684 6020 138740 6030
rect 138684 5926 138740 5964
rect 138348 5294 138350 5346
rect 138402 5294 138404 5346
rect 138012 5236 138068 5246
rect 138012 5142 138068 5180
rect 138348 5236 138404 5294
rect 138348 5170 138404 5180
rect 137788 4452 137844 4462
rect 137452 4450 137844 4452
rect 137452 4398 137790 4450
rect 137842 4398 137844 4450
rect 137452 4396 137844 4398
rect 135100 3444 135156 3454
rect 136444 3444 136500 3454
rect 133364 3388 133476 3444
rect 134764 3442 135156 3444
rect 134764 3390 135102 3442
rect 135154 3390 135156 3442
rect 134764 3388 135156 3390
rect 133308 3350 133364 3388
rect 133420 800 133476 3388
rect 135100 3378 135156 3388
rect 136108 3442 136500 3444
rect 136108 3390 136446 3442
rect 136498 3390 136500 3442
rect 136108 3388 136500 3390
rect 136108 800 136164 3388
rect 136444 3378 136500 3388
rect 137452 800 137508 4396
rect 137788 4386 137844 4396
rect 138796 4228 138852 33068
rect 139244 33124 139300 33404
rect 139244 33058 139300 33068
rect 139356 33906 139412 33918
rect 139356 33854 139358 33906
rect 139410 33854 139412 33906
rect 139356 6132 139412 33854
rect 139580 33460 139636 33470
rect 139580 33366 139636 33404
rect 140140 33460 140196 33470
rect 140252 33460 140308 35758
rect 140700 35140 140756 35150
rect 140700 34018 140756 35084
rect 140812 35028 140868 39200
rect 141708 39060 141764 39200
rect 142044 39060 142100 39228
rect 141708 39004 142100 39060
rect 141036 38276 141092 38286
rect 140924 36260 140980 36270
rect 140924 36166 140980 36204
rect 141036 35812 141092 38220
rect 141820 37268 141876 37278
rect 141820 36484 141876 37212
rect 142380 36484 142436 39228
rect 142576 39200 142688 40000
rect 143472 39200 143584 40000
rect 144368 39200 144480 40000
rect 145264 39200 145376 40000
rect 142604 36596 142660 39200
rect 142604 36530 142660 36540
rect 143276 36484 143332 36494
rect 142380 36428 142548 36484
rect 141820 36352 141876 36428
rect 142156 36372 142212 36382
rect 142492 36372 142548 36428
rect 143052 36372 143108 36382
rect 142492 36370 143108 36372
rect 142492 36318 143054 36370
rect 143106 36318 143108 36370
rect 142492 36316 143108 36318
rect 142156 36278 142212 36316
rect 141036 35746 141092 35756
rect 142604 35700 142660 35710
rect 141596 35698 142660 35700
rect 141596 35646 142606 35698
rect 142658 35646 142660 35698
rect 141596 35644 142660 35646
rect 141596 35586 141652 35644
rect 142604 35634 142660 35644
rect 141596 35534 141598 35586
rect 141650 35534 141652 35586
rect 141596 35522 141652 35534
rect 142268 35474 142324 35486
rect 142268 35422 142270 35474
rect 142322 35422 142324 35474
rect 140812 34962 140868 34972
rect 141148 35252 141204 35262
rect 141148 34914 141204 35196
rect 141708 35028 141764 35038
rect 141708 34934 141764 34972
rect 141148 34862 141150 34914
rect 141202 34862 141204 34914
rect 141148 34850 141204 34862
rect 140700 33966 140702 34018
rect 140754 33966 140756 34018
rect 140700 33954 140756 33966
rect 141820 34132 141876 34142
rect 141820 34018 141876 34076
rect 141820 33966 141822 34018
rect 141874 33966 141876 34018
rect 140140 33458 140308 33460
rect 140140 33406 140142 33458
rect 140194 33406 140308 33458
rect 140140 33404 140308 33406
rect 140140 33394 140196 33404
rect 141820 32452 141876 33966
rect 141820 32386 141876 32396
rect 141484 7586 141540 7598
rect 141484 7534 141486 7586
rect 141538 7534 141540 7586
rect 139132 6018 139188 6030
rect 139132 5966 139134 6018
rect 139186 5966 139188 6018
rect 138908 5460 138964 5470
rect 138908 5010 138964 5404
rect 138908 4958 138910 5010
rect 138962 4958 138964 5010
rect 138908 4946 138964 4958
rect 139132 5122 139188 5966
rect 139356 5906 139412 6076
rect 139356 5854 139358 5906
rect 139410 5854 139412 5906
rect 139356 5842 139412 5854
rect 139916 6804 139972 6814
rect 139692 5684 139748 5694
rect 139692 5590 139748 5628
rect 139692 5460 139748 5470
rect 139692 5234 139748 5404
rect 139692 5182 139694 5234
rect 139746 5182 139748 5234
rect 139692 5170 139748 5182
rect 139132 5070 139134 5122
rect 139186 5070 139188 5122
rect 139132 5012 139188 5070
rect 139132 4946 139188 4956
rect 139020 4900 139076 4910
rect 138908 4228 138964 4238
rect 138796 4226 138964 4228
rect 138796 4174 138910 4226
rect 138962 4174 138964 4226
rect 138796 4172 138964 4174
rect 138908 4162 138964 4172
rect 139020 3668 139076 4844
rect 139020 3536 139076 3612
rect 139916 3892 139972 6748
rect 141260 6580 141316 6590
rect 141260 6466 141316 6524
rect 141260 6414 141262 6466
rect 141314 6414 141316 6466
rect 140252 6132 140308 6142
rect 140252 6038 140308 6076
rect 140812 5908 140868 5918
rect 140140 5236 140196 5246
rect 140140 5142 140196 5180
rect 140812 5234 140868 5852
rect 141260 5796 141316 6414
rect 141372 5908 141428 5918
rect 141372 5814 141428 5852
rect 141260 5730 141316 5740
rect 140812 5182 140814 5234
rect 140866 5182 140868 5234
rect 140812 5170 140868 5182
rect 141372 5684 141428 5694
rect 141372 5234 141428 5628
rect 141372 5182 141374 5234
rect 141426 5182 141428 5234
rect 141372 5170 141428 5182
rect 141484 4452 141540 7534
rect 141820 7474 141876 7486
rect 141820 7422 141822 7474
rect 141874 7422 141876 7474
rect 141820 6914 141876 7422
rect 141820 6862 141822 6914
rect 141874 6862 141876 6914
rect 141820 6850 141876 6862
rect 142156 6916 142212 6926
rect 142268 6916 142324 35422
rect 142380 34244 142436 34254
rect 142380 34018 142436 34188
rect 142380 33966 142382 34018
rect 142434 33966 142436 34018
rect 142380 28532 142436 33966
rect 142716 33458 142772 36316
rect 143052 36306 143108 36316
rect 142828 35812 142884 35822
rect 142828 35026 142884 35756
rect 142828 34974 142830 35026
rect 142882 34974 142884 35026
rect 142828 34962 142884 34974
rect 142940 35810 142996 35822
rect 142940 35758 142942 35810
rect 142994 35758 142996 35810
rect 142940 35252 142996 35758
rect 143164 35812 143220 35822
rect 143164 35718 143220 35756
rect 143276 35252 143332 36428
rect 142940 34132 142996 35196
rect 143164 35196 143332 35252
rect 143052 34244 143108 34254
rect 143052 34150 143108 34188
rect 142940 34038 142996 34076
rect 142716 33406 142718 33458
rect 142770 33406 142772 33458
rect 142716 33394 142772 33406
rect 143164 31948 143220 35196
rect 143276 35028 143332 35038
rect 143500 35028 143556 39200
rect 143276 35026 143556 35028
rect 143276 34974 143278 35026
rect 143330 34974 143556 35026
rect 143276 34972 143556 34974
rect 143276 34962 143332 34972
rect 143500 34804 143556 34972
rect 143724 37044 143780 37054
rect 143724 35026 143780 36988
rect 144172 36596 144228 36606
rect 143724 34974 143726 35026
rect 143778 34974 143780 35026
rect 143724 34962 143780 34974
rect 143836 36594 144228 36596
rect 143836 36542 144174 36594
rect 144226 36542 144228 36594
rect 143836 36540 144228 36542
rect 143500 34738 143556 34748
rect 143724 34132 143780 34142
rect 143836 34132 143892 36540
rect 144172 36530 144228 36540
rect 143948 35586 144004 35598
rect 143948 35534 143950 35586
rect 144002 35534 144004 35586
rect 143948 35252 144004 35534
rect 143948 35186 144004 35196
rect 143724 34130 143892 34132
rect 143724 34078 143726 34130
rect 143778 34078 143892 34130
rect 143724 34076 143892 34078
rect 143724 34066 143780 34076
rect 144396 34020 144452 39200
rect 145292 36708 145348 39200
rect 145292 36642 145348 36652
rect 146188 36708 146244 36718
rect 145740 36484 145796 36494
rect 145740 36390 145796 36428
rect 145292 36370 145348 36382
rect 145292 36318 145294 36370
rect 145346 36318 145348 36370
rect 144956 36260 145012 36270
rect 144956 36258 145124 36260
rect 144956 36206 144958 36258
rect 145010 36206 145124 36258
rect 144956 36204 145124 36206
rect 144956 36194 145012 36204
rect 144956 35586 145012 35598
rect 144956 35534 144958 35586
rect 145010 35534 145012 35586
rect 144732 34804 144788 34814
rect 144732 34710 144788 34748
rect 144396 33954 144452 33964
rect 144620 34692 144676 34702
rect 144060 33906 144116 33918
rect 144060 33854 144062 33906
rect 144114 33854 144116 33906
rect 143164 31892 143332 31948
rect 142380 28466 142436 28476
rect 142380 7586 142436 7598
rect 142380 7534 142382 7586
rect 142434 7534 142436 7586
rect 142380 7364 142436 7534
rect 142380 7298 142436 7308
rect 142492 7476 142548 7486
rect 142156 6914 142268 6916
rect 142156 6862 142158 6914
rect 142210 6862 142268 6914
rect 142156 6860 142268 6862
rect 142156 6850 142212 6860
rect 142268 6784 142324 6860
rect 142492 6578 142548 7420
rect 142492 6526 142494 6578
rect 142546 6526 142548 6578
rect 142492 6468 142548 6526
rect 142268 5908 142324 5918
rect 141932 5796 141988 5806
rect 141932 5702 141988 5740
rect 141708 5122 141764 5134
rect 141708 5070 141710 5122
rect 141762 5070 141764 5122
rect 141708 4900 141764 5070
rect 142268 5122 142324 5852
rect 142492 5908 142548 6412
rect 142604 7474 142660 7486
rect 142604 7422 142606 7474
rect 142658 7422 142660 7474
rect 142604 6132 142660 7422
rect 143164 7252 143220 7262
rect 142716 6580 142772 6590
rect 142716 6486 142772 6524
rect 142604 6066 142660 6076
rect 142716 6018 142772 6030
rect 142716 5966 142718 6018
rect 142770 5966 142772 6018
rect 142604 5908 142660 5918
rect 142492 5906 142660 5908
rect 142492 5854 142606 5906
rect 142658 5854 142660 5906
rect 142492 5852 142660 5854
rect 142492 5796 142548 5852
rect 142604 5842 142660 5852
rect 142492 5730 142548 5740
rect 142716 5460 142772 5966
rect 142268 5070 142270 5122
rect 142322 5070 142324 5122
rect 142268 5058 142324 5070
rect 142604 5404 142772 5460
rect 141708 4834 141764 4844
rect 142604 4900 142660 5404
rect 142716 5234 142772 5246
rect 142716 5182 142718 5234
rect 142770 5182 142772 5234
rect 142716 5012 142772 5182
rect 142716 4946 142772 4956
rect 142604 4834 142660 4844
rect 143164 4900 143220 7196
rect 143164 4834 143220 4844
rect 141484 4386 141540 4396
rect 141820 4450 141876 4462
rect 141820 4398 141822 4450
rect 141874 4398 141876 4450
rect 141260 4228 141316 4238
rect 141820 4228 141876 4398
rect 141260 4226 141876 4228
rect 141260 4174 141262 4226
rect 141314 4174 141876 4226
rect 141260 4172 141876 4174
rect 143164 4228 143220 4238
rect 143276 4228 143332 31892
rect 144060 8428 144116 33854
rect 143388 8372 144116 8428
rect 143388 6020 143444 8372
rect 143836 7924 143892 7934
rect 143612 7140 143668 7150
rect 143500 6468 143556 6478
rect 143500 6374 143556 6412
rect 143388 5906 143444 5964
rect 143388 5854 143390 5906
rect 143442 5854 143444 5906
rect 143388 5842 143444 5854
rect 143500 5122 143556 5134
rect 143500 5070 143502 5122
rect 143554 5070 143556 5122
rect 143500 4900 143556 5070
rect 143500 4834 143556 4844
rect 143612 4564 143668 7084
rect 143724 6132 143780 6142
rect 143724 6038 143780 6076
rect 143724 4564 143780 4574
rect 143612 4562 143780 4564
rect 143612 4510 143726 4562
rect 143778 4510 143780 4562
rect 143612 4508 143780 4510
rect 143724 4498 143780 4508
rect 143164 4226 143332 4228
rect 143164 4174 143166 4226
rect 143218 4174 143332 4226
rect 143164 4172 143332 4174
rect 141260 4162 141316 4172
rect 139916 3836 140420 3892
rect 139916 3666 139972 3836
rect 139916 3614 139918 3666
rect 139970 3614 139972 3666
rect 139916 3602 139972 3614
rect 140140 3668 140196 3678
rect 138012 3444 138068 3454
rect 138012 3350 138068 3388
rect 140140 800 140196 3612
rect 140364 3554 140420 3836
rect 141036 3668 141092 3678
rect 141036 3574 141092 3612
rect 140364 3502 140366 3554
rect 140418 3502 140420 3554
rect 140364 3490 140420 3502
rect 141484 800 141540 4172
rect 143164 4162 143220 4172
rect 143724 3332 143780 3342
rect 143836 3332 143892 7868
rect 143948 6916 144004 6926
rect 143948 6690 144004 6860
rect 143948 6638 143950 6690
rect 144002 6638 144004 6690
rect 143948 6626 144004 6638
rect 144508 5236 144564 5246
rect 144508 5142 144564 5180
rect 144172 4898 144228 4910
rect 144172 4846 144174 4898
rect 144226 4846 144228 4898
rect 144060 4452 144116 4462
rect 144172 4452 144228 4846
rect 144060 4450 144228 4452
rect 144060 4398 144062 4450
rect 144114 4398 144228 4450
rect 144060 4396 144228 4398
rect 144060 4386 144116 4396
rect 144172 3668 144228 3678
rect 144060 3556 144116 3566
rect 144060 3462 144116 3500
rect 143724 3330 143892 3332
rect 143724 3278 143726 3330
rect 143778 3278 143892 3330
rect 143724 3276 143892 3278
rect 143724 3266 143780 3276
rect 144172 800 144228 3612
rect 144620 3666 144676 34636
rect 144956 31948 145012 35534
rect 145068 34130 145124 36204
rect 145292 34692 145348 36318
rect 146188 35924 146244 36652
rect 147532 36596 147588 36606
rect 147532 36502 147588 36540
rect 146860 36482 146916 36494
rect 146860 36430 146862 36482
rect 146914 36430 146916 36482
rect 146860 36372 146916 36430
rect 146860 36306 146916 36316
rect 148492 36092 148756 36102
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148492 36026 148756 36036
rect 146188 35810 146244 35868
rect 146860 35924 146916 35934
rect 146860 35830 146916 35868
rect 146188 35758 146190 35810
rect 146242 35758 146244 35810
rect 146188 35746 146244 35758
rect 145292 34626 145348 34636
rect 145628 34692 145684 34702
rect 145628 34598 145684 34636
rect 148492 34524 148756 34534
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148492 34458 148756 34468
rect 145068 34078 145070 34130
rect 145122 34078 145124 34130
rect 145068 34066 145124 34078
rect 145628 34020 145684 34030
rect 145628 33926 145684 33964
rect 148492 32956 148756 32966
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148492 32890 148756 32900
rect 144844 31892 145012 31948
rect 147868 32788 147924 32798
rect 144844 31668 144900 31892
rect 144844 31602 144900 31612
rect 145964 7812 146020 7822
rect 145292 6132 145348 6142
rect 144844 6020 144900 6030
rect 144844 5926 144900 5964
rect 145180 5122 145236 5134
rect 145180 5070 145182 5122
rect 145234 5070 145236 5122
rect 145068 5010 145124 5022
rect 145068 4958 145070 5010
rect 145122 4958 145124 5010
rect 145068 4900 145124 4958
rect 145068 4834 145124 4844
rect 145180 5012 145236 5070
rect 145180 4452 145236 4956
rect 145180 4386 145236 4396
rect 145292 4340 145348 6076
rect 145852 5236 145908 5246
rect 145852 5142 145908 5180
rect 145964 4564 146020 7756
rect 145628 4452 145684 4490
rect 145628 4386 145684 4396
rect 145964 4450 146020 4508
rect 145964 4398 145966 4450
rect 146018 4398 146020 4450
rect 145964 4386 146020 4398
rect 146524 6356 146580 6366
rect 146524 5234 146580 6300
rect 146524 5182 146526 5234
rect 146578 5182 146580 5234
rect 145404 4340 145460 4350
rect 145292 4338 145460 4340
rect 145292 4286 145406 4338
rect 145458 4286 145460 4338
rect 145292 4284 145460 4286
rect 145404 4274 145460 4284
rect 145628 4228 145684 4238
rect 144620 3614 144622 3666
rect 144674 3614 144676 3666
rect 144620 3602 144676 3614
rect 145068 4114 145124 4126
rect 145068 4062 145070 4114
rect 145122 4062 145124 4114
rect 145068 3556 145124 4062
rect 145068 3490 145124 3500
rect 145628 3444 145684 4172
rect 146524 3556 146580 5182
rect 147868 5236 147924 32732
rect 148492 31388 148756 31398
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148492 31322 148756 31332
rect 147980 31108 148036 31118
rect 147980 6132 148036 31052
rect 148492 29820 148756 29830
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148492 29754 148756 29764
rect 148492 28252 148756 28262
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148492 28186 148756 28196
rect 148492 26684 148756 26694
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148492 26618 148756 26628
rect 148492 25116 148756 25126
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148492 25050 148756 25060
rect 148492 23548 148756 23558
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148492 23482 148756 23492
rect 148492 21980 148756 21990
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148492 21914 148756 21924
rect 148492 20412 148756 20422
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148492 20346 148756 20356
rect 148492 18844 148756 18854
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148492 18778 148756 18788
rect 148492 17276 148756 17286
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148492 17210 148756 17220
rect 148492 15708 148756 15718
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148492 15642 148756 15652
rect 148492 14140 148756 14150
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148492 14074 148756 14084
rect 148492 12572 148756 12582
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148492 12506 148756 12516
rect 148492 11004 148756 11014
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148492 10938 148756 10948
rect 148492 9436 148756 9446
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148492 9370 148756 9380
rect 148492 7868 148756 7878
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148492 7802 148756 7812
rect 148492 6300 148756 6310
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148492 6234 148756 6244
rect 147980 6066 148036 6076
rect 147868 5170 147924 5180
rect 148492 4732 148756 4742
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148492 4666 148756 4676
rect 146748 4564 146804 4574
rect 146748 4470 146804 4508
rect 147196 4228 147252 4238
rect 147196 4134 147252 4172
rect 147532 3668 147588 3678
rect 147532 3574 147588 3612
rect 146860 3556 146916 3566
rect 146524 3554 146916 3556
rect 146524 3502 146862 3554
rect 146914 3502 146916 3554
rect 146524 3500 146916 3502
rect 146860 3490 146916 3500
rect 145516 3442 145684 3444
rect 145516 3390 145630 3442
rect 145682 3390 145684 3442
rect 145516 3388 145684 3390
rect 145516 800 145572 3388
rect 145628 3378 145684 3388
rect 148492 3164 148756 3174
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148492 3098 148756 3108
rect 121548 700 122164 756
rect 122640 0 122752 800
rect 123984 0 124096 800
rect 125328 0 125440 800
rect 126672 0 126784 800
rect 128016 0 128128 800
rect 129360 0 129472 800
rect 130704 0 130816 800
rect 132048 0 132160 800
rect 133392 0 133504 800
rect 134736 0 134848 800
rect 136080 0 136192 800
rect 137424 0 137536 800
rect 138768 0 138880 800
rect 140112 0 140224 800
rect 141456 0 141568 800
rect 142800 0 142912 800
rect 144144 0 144256 800
rect 145488 0 145600 800
<< via2 >>
rect 6076 36258 6132 36260
rect 6076 36206 6078 36258
rect 6078 36206 6130 36258
rect 6130 36206 6132 36258
rect 6076 36204 6132 36206
rect 6636 36204 6692 36260
rect 6636 34636 6692 34692
rect 7868 35868 7924 35924
rect 8428 36876 8484 36932
rect 9100 36876 9156 36932
rect 7308 35084 7364 35140
rect 8428 35084 8484 35140
rect 9660 35922 9716 35924
rect 9660 35870 9662 35922
rect 9662 35870 9714 35922
rect 9714 35870 9716 35922
rect 9660 35868 9716 35870
rect 8876 34748 8932 34804
rect 9996 36258 10052 36260
rect 9996 36206 9998 36258
rect 9998 36206 10050 36258
rect 10050 36206 10052 36258
rect 9996 36204 10052 36206
rect 10780 36204 10836 36260
rect 9884 34972 9940 35028
rect 10332 35026 10388 35028
rect 10332 34974 10334 35026
rect 10334 34974 10386 35026
rect 10386 34974 10388 35026
rect 10332 34972 10388 34974
rect 11788 36316 11844 36372
rect 13916 36594 13972 36596
rect 13916 36542 13918 36594
rect 13918 36542 13970 36594
rect 13970 36542 13972 36594
rect 13916 36540 13972 36542
rect 12796 35756 12852 35812
rect 12908 36316 12964 36372
rect 11676 34972 11732 35028
rect 10780 34860 10836 34916
rect 8092 33852 8148 33908
rect 13356 35308 13412 35364
rect 15372 36540 15428 36596
rect 14252 35308 14308 35364
rect 16604 36988 16660 37044
rect 14924 34524 14980 34580
rect 8540 33852 8596 33908
rect 14588 33964 14644 34020
rect 15036 34300 15092 34356
rect 15596 34690 15652 34692
rect 15596 34638 15598 34690
rect 15598 34638 15650 34690
rect 15650 34638 15652 34690
rect 15596 34636 15652 34638
rect 15036 34018 15092 34020
rect 15036 33966 15038 34018
rect 15038 33966 15090 34018
rect 15090 33966 15092 34018
rect 15036 33964 15092 33966
rect 9884 32620 9940 32676
rect 11676 32620 11732 32676
rect 7196 31836 7252 31892
rect 16156 34636 16212 34692
rect 16492 34690 16548 34692
rect 16492 34638 16494 34690
rect 16494 34638 16546 34690
rect 16546 34638 16548 34690
rect 16492 34636 16548 34638
rect 16828 34412 16884 34468
rect 15932 34354 15988 34356
rect 15932 34302 15934 34354
rect 15934 34302 15986 34354
rect 15986 34302 15988 34354
rect 15932 34300 15988 34302
rect 19622 36874 19678 36876
rect 19622 36822 19624 36874
rect 19624 36822 19676 36874
rect 19676 36822 19678 36874
rect 19622 36820 19678 36822
rect 19726 36874 19782 36876
rect 19726 36822 19728 36874
rect 19728 36822 19780 36874
rect 19780 36822 19782 36874
rect 19726 36820 19782 36822
rect 19830 36874 19886 36876
rect 19830 36822 19832 36874
rect 19832 36822 19884 36874
rect 19884 36822 19886 36874
rect 19830 36820 19886 36822
rect 16940 34300 16996 34356
rect 17836 34748 17892 34804
rect 18620 36258 18676 36260
rect 18620 36206 18622 36258
rect 18622 36206 18674 36258
rect 18674 36206 18676 36258
rect 18620 36204 18676 36206
rect 18284 35980 18340 36036
rect 19068 35420 19124 35476
rect 18620 35084 18676 35140
rect 18396 34636 18452 34692
rect 18284 34354 18340 34356
rect 18284 34302 18286 34354
rect 18286 34302 18338 34354
rect 18338 34302 18340 34354
rect 18284 34300 18340 34302
rect 18172 33180 18228 33236
rect 18956 34802 19012 34804
rect 18956 34750 18958 34802
rect 18958 34750 19010 34802
rect 19010 34750 19012 34802
rect 18956 34748 19012 34750
rect 19740 35810 19796 35812
rect 19740 35758 19742 35810
rect 19742 35758 19794 35810
rect 19794 35758 19796 35810
rect 19740 35756 19796 35758
rect 19628 35420 19684 35476
rect 19622 35306 19678 35308
rect 19622 35254 19624 35306
rect 19624 35254 19676 35306
rect 19676 35254 19678 35306
rect 19622 35252 19678 35254
rect 19726 35306 19782 35308
rect 19726 35254 19728 35306
rect 19728 35254 19780 35306
rect 19780 35254 19782 35306
rect 19726 35252 19782 35254
rect 19830 35306 19886 35308
rect 19830 35254 19832 35306
rect 19832 35254 19884 35306
rect 19884 35254 19886 35306
rect 19830 35252 19886 35254
rect 19740 34636 19796 34692
rect 19852 34860 19908 34916
rect 19852 34412 19908 34468
rect 20636 36428 20692 36484
rect 20188 36204 20244 36260
rect 19964 34188 20020 34244
rect 19622 33738 19678 33740
rect 19622 33686 19624 33738
rect 19624 33686 19676 33738
rect 19676 33686 19678 33738
rect 19622 33684 19678 33686
rect 19726 33738 19782 33740
rect 19726 33686 19728 33738
rect 19728 33686 19780 33738
rect 19780 33686 19782 33738
rect 19726 33684 19782 33686
rect 19830 33738 19886 33740
rect 19830 33686 19832 33738
rect 19832 33686 19884 33738
rect 19884 33686 19886 33738
rect 19830 33684 19886 33686
rect 19740 33068 19796 33124
rect 19068 32956 19124 33012
rect 19622 32170 19678 32172
rect 19622 32118 19624 32170
rect 19624 32118 19676 32170
rect 19676 32118 19678 32170
rect 19622 32116 19678 32118
rect 19726 32170 19782 32172
rect 19726 32118 19728 32170
rect 19728 32118 19780 32170
rect 19780 32118 19782 32170
rect 19726 32116 19782 32118
rect 19830 32170 19886 32172
rect 19830 32118 19832 32170
rect 19832 32118 19884 32170
rect 19884 32118 19886 32170
rect 19830 32116 19886 32118
rect 19622 30602 19678 30604
rect 19622 30550 19624 30602
rect 19624 30550 19676 30602
rect 19676 30550 19678 30602
rect 19622 30548 19678 30550
rect 19726 30602 19782 30604
rect 19726 30550 19728 30602
rect 19728 30550 19780 30602
rect 19780 30550 19782 30602
rect 19726 30548 19782 30550
rect 19830 30602 19886 30604
rect 19830 30550 19832 30602
rect 19832 30550 19884 30602
rect 19884 30550 19886 30602
rect 19830 30548 19886 30550
rect 18396 29596 18452 29652
rect 19622 29034 19678 29036
rect 19622 28982 19624 29034
rect 19624 28982 19676 29034
rect 19676 28982 19678 29034
rect 19622 28980 19678 28982
rect 19726 29034 19782 29036
rect 19726 28982 19728 29034
rect 19728 28982 19780 29034
rect 19780 28982 19782 29034
rect 19726 28980 19782 28982
rect 19830 29034 19886 29036
rect 19830 28982 19832 29034
rect 19832 28982 19884 29034
rect 19884 28982 19886 29034
rect 19830 28980 19886 28982
rect 19622 27466 19678 27468
rect 19622 27414 19624 27466
rect 19624 27414 19676 27466
rect 19676 27414 19678 27466
rect 19622 27412 19678 27414
rect 19726 27466 19782 27468
rect 19726 27414 19728 27466
rect 19728 27414 19780 27466
rect 19780 27414 19782 27466
rect 19726 27412 19782 27414
rect 19830 27466 19886 27468
rect 19830 27414 19832 27466
rect 19832 27414 19884 27466
rect 19884 27414 19886 27466
rect 19830 27412 19886 27414
rect 18508 26012 18564 26068
rect 17948 17612 18004 17668
rect 15148 7532 15204 7588
rect 11676 6748 11732 6804
rect 14924 7420 14980 7476
rect 7420 6412 7476 6468
rect 10892 6578 10948 6580
rect 10892 6526 10894 6578
rect 10894 6526 10946 6578
rect 10946 6526 10948 6578
rect 10892 6524 10948 6526
rect 13580 6524 13636 6580
rect 6860 4396 6916 4452
rect 5852 3948 5908 4004
rect 6412 3948 6468 4004
rect 7420 4450 7476 4452
rect 7420 4398 7422 4450
rect 7422 4398 7474 4450
rect 7474 4398 7476 4450
rect 7420 4396 7476 4398
rect 6636 4172 6692 4228
rect 6412 3612 6468 3668
rect 6300 3554 6356 3556
rect 6300 3502 6302 3554
rect 6302 3502 6354 3554
rect 6354 3502 6356 3554
rect 6300 3500 6356 3502
rect 8316 4508 8372 4564
rect 6860 3442 6916 3444
rect 6860 3390 6862 3442
rect 6862 3390 6914 3442
rect 6914 3390 6916 3442
rect 6860 3388 6916 3390
rect 8764 4226 8820 4228
rect 8764 4174 8766 4226
rect 8766 4174 8818 4226
rect 8818 4174 8820 4226
rect 8764 4172 8820 4174
rect 10220 5122 10276 5124
rect 10220 5070 10222 5122
rect 10222 5070 10274 5122
rect 10274 5070 10276 5122
rect 10220 5068 10276 5070
rect 10108 4508 10164 4564
rect 11228 6466 11284 6468
rect 11228 6414 11230 6466
rect 11230 6414 11282 6466
rect 11282 6414 11284 6466
rect 11228 6412 11284 6414
rect 12908 6412 12964 6468
rect 11676 5122 11732 5124
rect 11676 5070 11678 5122
rect 11678 5070 11730 5122
rect 11730 5070 11732 5122
rect 11676 5068 11732 5070
rect 11788 5010 11844 5012
rect 11788 4958 11790 5010
rect 11790 4958 11842 5010
rect 11842 4958 11844 5010
rect 11788 4956 11844 4958
rect 11116 4898 11172 4900
rect 11116 4846 11118 4898
rect 11118 4846 11170 4898
rect 11170 4846 11172 4898
rect 11116 4844 11172 4846
rect 10332 4508 10388 4564
rect 9772 4396 9828 4452
rect 5740 2492 5796 2548
rect 8876 3164 8932 3220
rect 11004 4450 11060 4452
rect 11004 4398 11006 4450
rect 11006 4398 11058 4450
rect 11058 4398 11060 4450
rect 11004 4396 11060 4398
rect 10220 4172 10276 4228
rect 11340 3666 11396 3668
rect 11340 3614 11342 3666
rect 11342 3614 11394 3666
rect 11394 3614 11396 3666
rect 11340 3612 11396 3614
rect 11116 3500 11172 3556
rect 9884 3388 9940 3444
rect 10108 3442 10164 3444
rect 10108 3390 10110 3442
rect 10110 3390 10162 3442
rect 10162 3390 10164 3442
rect 10108 3388 10164 3390
rect 10332 3276 10388 3332
rect 12236 5010 12292 5012
rect 12236 4958 12238 5010
rect 12238 4958 12290 5010
rect 12290 4958 12292 5010
rect 12236 4956 12292 4958
rect 12012 4562 12068 4564
rect 12012 4510 12014 4562
rect 12014 4510 12066 4562
rect 12066 4510 12068 4562
rect 12012 4508 12068 4510
rect 12684 5234 12740 5236
rect 12684 5182 12686 5234
rect 12686 5182 12738 5234
rect 12738 5182 12740 5234
rect 12684 5180 12740 5182
rect 12460 4956 12516 5012
rect 13580 5180 13636 5236
rect 11900 3500 11956 3556
rect 12348 3500 12404 3556
rect 13916 3948 13972 4004
rect 14364 3948 14420 4004
rect 16604 7196 16660 7252
rect 16156 6412 16212 6468
rect 16044 6130 16100 6132
rect 16044 6078 16046 6130
rect 16046 6078 16098 6130
rect 16098 6078 16100 6130
rect 16044 6076 16100 6078
rect 16716 6076 16772 6132
rect 16828 6412 16884 6468
rect 15820 5906 15876 5908
rect 15820 5854 15822 5906
rect 15822 5854 15874 5906
rect 15874 5854 15876 5906
rect 15820 5852 15876 5854
rect 15820 4956 15876 5012
rect 16492 4956 16548 5012
rect 17836 6130 17892 6132
rect 17836 6078 17838 6130
rect 17838 6078 17890 6130
rect 17890 6078 17892 6130
rect 17836 6076 17892 6078
rect 19622 25898 19678 25900
rect 19622 25846 19624 25898
rect 19624 25846 19676 25898
rect 19676 25846 19678 25898
rect 19622 25844 19678 25846
rect 19726 25898 19782 25900
rect 19726 25846 19728 25898
rect 19728 25846 19780 25898
rect 19780 25846 19782 25898
rect 19726 25844 19782 25846
rect 19830 25898 19886 25900
rect 19830 25846 19832 25898
rect 19832 25846 19884 25898
rect 19884 25846 19886 25898
rect 19830 25844 19886 25846
rect 19622 24330 19678 24332
rect 19622 24278 19624 24330
rect 19624 24278 19676 24330
rect 19676 24278 19678 24330
rect 19622 24276 19678 24278
rect 19726 24330 19782 24332
rect 19726 24278 19728 24330
rect 19728 24278 19780 24330
rect 19780 24278 19782 24330
rect 19726 24276 19782 24278
rect 19830 24330 19886 24332
rect 19830 24278 19832 24330
rect 19832 24278 19884 24330
rect 19884 24278 19886 24330
rect 19830 24276 19886 24278
rect 19622 22762 19678 22764
rect 19622 22710 19624 22762
rect 19624 22710 19676 22762
rect 19676 22710 19678 22762
rect 19622 22708 19678 22710
rect 19726 22762 19782 22764
rect 19726 22710 19728 22762
rect 19728 22710 19780 22762
rect 19780 22710 19782 22762
rect 19726 22708 19782 22710
rect 19830 22762 19886 22764
rect 19830 22710 19832 22762
rect 19832 22710 19884 22762
rect 19884 22710 19886 22762
rect 19830 22708 19886 22710
rect 19622 21194 19678 21196
rect 19622 21142 19624 21194
rect 19624 21142 19676 21194
rect 19676 21142 19678 21194
rect 19622 21140 19678 21142
rect 19726 21194 19782 21196
rect 19726 21142 19728 21194
rect 19728 21142 19780 21194
rect 19780 21142 19782 21194
rect 19726 21140 19782 21142
rect 19830 21194 19886 21196
rect 19830 21142 19832 21194
rect 19832 21142 19884 21194
rect 19884 21142 19886 21194
rect 19830 21140 19886 21142
rect 21420 36370 21476 36372
rect 21420 36318 21422 36370
rect 21422 36318 21474 36370
rect 21474 36318 21476 36370
rect 21420 36316 21476 36318
rect 20412 35698 20468 35700
rect 20412 35646 20414 35698
rect 20414 35646 20466 35698
rect 20466 35646 20468 35698
rect 20412 35644 20468 35646
rect 21420 35922 21476 35924
rect 21420 35870 21422 35922
rect 21422 35870 21474 35922
rect 21474 35870 21476 35922
rect 21420 35868 21476 35870
rect 22204 36370 22260 36372
rect 22204 36318 22206 36370
rect 22206 36318 22258 36370
rect 22258 36318 22260 36370
rect 22204 36316 22260 36318
rect 21868 35980 21924 36036
rect 20636 35084 20692 35140
rect 20748 34690 20804 34692
rect 20748 34638 20750 34690
rect 20750 34638 20802 34690
rect 20802 34638 20804 34690
rect 20748 34636 20804 34638
rect 20748 34188 20804 34244
rect 20524 32956 20580 33012
rect 20076 26012 20132 26068
rect 19622 19626 19678 19628
rect 19622 19574 19624 19626
rect 19624 19574 19676 19626
rect 19676 19574 19678 19626
rect 19622 19572 19678 19574
rect 19726 19626 19782 19628
rect 19726 19574 19728 19626
rect 19728 19574 19780 19626
rect 19780 19574 19782 19626
rect 19726 19572 19782 19574
rect 19830 19626 19886 19628
rect 19830 19574 19832 19626
rect 19832 19574 19884 19626
rect 19884 19574 19886 19626
rect 19830 19572 19886 19574
rect 19622 18058 19678 18060
rect 19622 18006 19624 18058
rect 19624 18006 19676 18058
rect 19676 18006 19678 18058
rect 19622 18004 19678 18006
rect 19726 18058 19782 18060
rect 19726 18006 19728 18058
rect 19728 18006 19780 18058
rect 19780 18006 19782 18058
rect 19726 18004 19782 18006
rect 19830 18058 19886 18060
rect 19830 18006 19832 18058
rect 19832 18006 19884 18058
rect 19884 18006 19886 18058
rect 19830 18004 19886 18006
rect 19622 16490 19678 16492
rect 19622 16438 19624 16490
rect 19624 16438 19676 16490
rect 19676 16438 19678 16490
rect 19622 16436 19678 16438
rect 19726 16490 19782 16492
rect 19726 16438 19728 16490
rect 19728 16438 19780 16490
rect 19780 16438 19782 16490
rect 19726 16436 19782 16438
rect 19830 16490 19886 16492
rect 19830 16438 19832 16490
rect 19832 16438 19884 16490
rect 19884 16438 19886 16490
rect 19830 16436 19886 16438
rect 19622 14922 19678 14924
rect 19622 14870 19624 14922
rect 19624 14870 19676 14922
rect 19676 14870 19678 14922
rect 19622 14868 19678 14870
rect 19726 14922 19782 14924
rect 19726 14870 19728 14922
rect 19728 14870 19780 14922
rect 19780 14870 19782 14922
rect 19726 14868 19782 14870
rect 19830 14922 19886 14924
rect 19830 14870 19832 14922
rect 19832 14870 19884 14922
rect 19884 14870 19886 14922
rect 19830 14868 19886 14870
rect 19622 13354 19678 13356
rect 19622 13302 19624 13354
rect 19624 13302 19676 13354
rect 19676 13302 19678 13354
rect 19622 13300 19678 13302
rect 19726 13354 19782 13356
rect 19726 13302 19728 13354
rect 19728 13302 19780 13354
rect 19780 13302 19782 13354
rect 19726 13300 19782 13302
rect 19830 13354 19886 13356
rect 19830 13302 19832 13354
rect 19832 13302 19884 13354
rect 19884 13302 19886 13354
rect 19830 13300 19886 13302
rect 19622 11786 19678 11788
rect 19622 11734 19624 11786
rect 19624 11734 19676 11786
rect 19676 11734 19678 11786
rect 19622 11732 19678 11734
rect 19726 11786 19782 11788
rect 19726 11734 19728 11786
rect 19728 11734 19780 11786
rect 19780 11734 19782 11786
rect 19726 11732 19782 11734
rect 19830 11786 19886 11788
rect 19830 11734 19832 11786
rect 19832 11734 19884 11786
rect 19884 11734 19886 11786
rect 19830 11732 19886 11734
rect 19622 10218 19678 10220
rect 19622 10166 19624 10218
rect 19624 10166 19676 10218
rect 19676 10166 19678 10218
rect 19622 10164 19678 10166
rect 19726 10218 19782 10220
rect 19726 10166 19728 10218
rect 19728 10166 19780 10218
rect 19780 10166 19782 10218
rect 19726 10164 19782 10166
rect 19830 10218 19886 10220
rect 19830 10166 19832 10218
rect 19832 10166 19884 10218
rect 19884 10166 19886 10218
rect 19830 10164 19886 10166
rect 19622 8650 19678 8652
rect 19622 8598 19624 8650
rect 19624 8598 19676 8650
rect 19676 8598 19678 8650
rect 19622 8596 19678 8598
rect 19726 8650 19782 8652
rect 19726 8598 19728 8650
rect 19728 8598 19780 8650
rect 19780 8598 19782 8650
rect 19726 8596 19782 8598
rect 19830 8650 19886 8652
rect 19830 8598 19832 8650
rect 19832 8598 19884 8650
rect 19884 8598 19886 8650
rect 19830 8596 19886 8598
rect 18508 7644 18564 7700
rect 19964 7698 20020 7700
rect 19964 7646 19966 7698
rect 19966 7646 20018 7698
rect 20018 7646 20020 7698
rect 19964 7644 20020 7646
rect 19068 7586 19124 7588
rect 19068 7534 19070 7586
rect 19070 7534 19122 7586
rect 19122 7534 19124 7586
rect 19068 7532 19124 7534
rect 18172 7250 18228 7252
rect 18172 7198 18174 7250
rect 18174 7198 18226 7250
rect 18226 7198 18228 7250
rect 18172 7196 18228 7198
rect 18620 6748 18676 6804
rect 18396 5906 18452 5908
rect 18396 5854 18398 5906
rect 18398 5854 18450 5906
rect 18450 5854 18452 5906
rect 18396 5852 18452 5854
rect 17948 4844 18004 4900
rect 16604 3948 16660 4004
rect 16492 3724 16548 3780
rect 14476 3442 14532 3444
rect 14476 3390 14478 3442
rect 14478 3390 14530 3442
rect 14530 3390 14532 3442
rect 14476 3388 14532 3390
rect 15148 3388 15204 3444
rect 16268 3442 16324 3444
rect 16268 3390 16270 3442
rect 16270 3390 16322 3442
rect 16322 3390 16324 3442
rect 16268 3388 16324 3390
rect 16492 3388 16548 3444
rect 19622 7082 19678 7084
rect 19622 7030 19624 7082
rect 19624 7030 19676 7082
rect 19676 7030 19678 7082
rect 19622 7028 19678 7030
rect 19726 7082 19782 7084
rect 19726 7030 19728 7082
rect 19728 7030 19780 7082
rect 19780 7030 19782 7082
rect 19726 7028 19782 7030
rect 19830 7082 19886 7084
rect 19830 7030 19832 7082
rect 19832 7030 19884 7082
rect 19884 7030 19886 7082
rect 19830 7028 19886 7030
rect 19068 6748 19124 6804
rect 18956 6636 19012 6692
rect 18956 6076 19012 6132
rect 18732 5964 18788 6020
rect 19180 6076 19236 6132
rect 19622 5514 19678 5516
rect 19622 5462 19624 5514
rect 19624 5462 19676 5514
rect 19676 5462 19678 5514
rect 19622 5460 19678 5462
rect 19726 5514 19782 5516
rect 19726 5462 19728 5514
rect 19728 5462 19780 5514
rect 19780 5462 19782 5514
rect 19726 5460 19782 5462
rect 19830 5514 19886 5516
rect 19830 5462 19832 5514
rect 19832 5462 19884 5514
rect 19884 5462 19886 5514
rect 19830 5460 19886 5462
rect 17612 3442 17668 3444
rect 17612 3390 17614 3442
rect 17614 3390 17666 3442
rect 17666 3390 17668 3442
rect 17612 3388 17668 3390
rect 20300 6636 20356 6692
rect 20412 7196 20468 7252
rect 20748 7196 20804 7252
rect 20412 6524 20468 6580
rect 20748 6748 20804 6804
rect 20524 6130 20580 6132
rect 20524 6078 20526 6130
rect 20526 6078 20578 6130
rect 20578 6078 20580 6130
rect 20524 6076 20580 6078
rect 20636 5794 20692 5796
rect 20636 5742 20638 5794
rect 20638 5742 20690 5794
rect 20690 5742 20692 5794
rect 20636 5740 20692 5742
rect 20860 6690 20916 6692
rect 20860 6638 20862 6690
rect 20862 6638 20914 6690
rect 20914 6638 20916 6690
rect 20860 6636 20916 6638
rect 21868 35084 21924 35140
rect 21532 34412 21588 34468
rect 21868 34412 21924 34468
rect 22092 32956 22148 33012
rect 22204 29932 22260 29988
rect 22540 36316 22596 36372
rect 22540 35868 22596 35924
rect 22764 38892 22820 38948
rect 22876 36370 22932 36372
rect 22876 36318 22878 36370
rect 22878 36318 22930 36370
rect 22930 36318 22932 36370
rect 22876 36316 22932 36318
rect 22764 35644 22820 35700
rect 23100 35532 23156 35588
rect 24220 36652 24276 36708
rect 23884 35532 23940 35588
rect 24220 34636 24276 34692
rect 22876 34188 22932 34244
rect 23212 34242 23268 34244
rect 23212 34190 23214 34242
rect 23214 34190 23266 34242
rect 23266 34190 23268 34242
rect 23212 34188 23268 34190
rect 22316 10892 22372 10948
rect 23884 33964 23940 34020
rect 21308 5964 21364 6020
rect 21532 6466 21588 6468
rect 21532 6414 21534 6466
rect 21534 6414 21586 6466
rect 21586 6414 21588 6466
rect 21532 6412 21588 6414
rect 21196 5794 21252 5796
rect 21196 5742 21198 5794
rect 21198 5742 21250 5794
rect 21250 5742 21252 5794
rect 21196 5740 21252 5742
rect 21196 5180 21252 5236
rect 21980 6018 22036 6020
rect 21980 5966 21982 6018
rect 21982 5966 22034 6018
rect 22034 5966 22036 6018
rect 21980 5964 22036 5966
rect 21756 5234 21812 5236
rect 21756 5182 21758 5234
rect 21758 5182 21810 5234
rect 21810 5182 21812 5234
rect 21756 5180 21812 5182
rect 22204 5234 22260 5236
rect 22204 5182 22206 5234
rect 22206 5182 22258 5234
rect 22258 5182 22260 5234
rect 22204 5180 22260 5182
rect 21532 5068 21588 5124
rect 20300 4898 20356 4900
rect 20300 4846 20302 4898
rect 20302 4846 20354 4898
rect 20354 4846 20356 4898
rect 20300 4844 20356 4846
rect 21644 4898 21700 4900
rect 21644 4846 21646 4898
rect 21646 4846 21698 4898
rect 21698 4846 21700 4898
rect 21644 4844 21700 4846
rect 20524 4396 20580 4452
rect 19622 3946 19678 3948
rect 19622 3894 19624 3946
rect 19624 3894 19676 3946
rect 19676 3894 19678 3946
rect 19622 3892 19678 3894
rect 19726 3946 19782 3948
rect 19726 3894 19728 3946
rect 19728 3894 19780 3946
rect 19780 3894 19782 3946
rect 19726 3892 19782 3894
rect 19830 3946 19886 3948
rect 19830 3894 19832 3946
rect 19832 3894 19884 3946
rect 19884 3894 19886 3946
rect 19830 3892 19886 3894
rect 19404 3554 19460 3556
rect 19404 3502 19406 3554
rect 19406 3502 19458 3554
rect 19458 3502 19460 3554
rect 19404 3500 19460 3502
rect 21084 4450 21140 4452
rect 21084 4398 21086 4450
rect 21086 4398 21138 4450
rect 21138 4398 21140 4450
rect 21084 4396 21140 4398
rect 20524 3388 20580 3444
rect 24444 34412 24500 34468
rect 24892 35308 24948 35364
rect 24780 34412 24836 34468
rect 24892 34018 24948 34020
rect 24892 33966 24894 34018
rect 24894 33966 24946 34018
rect 24946 33966 24948 34018
rect 24892 33964 24948 33966
rect 25564 35308 25620 35364
rect 26908 36428 26964 36484
rect 27692 36594 27748 36596
rect 27692 36542 27694 36594
rect 27694 36542 27746 36594
rect 27746 36542 27748 36594
rect 27692 36540 27748 36542
rect 27580 36204 27636 36260
rect 27020 35868 27076 35924
rect 27804 35196 27860 35252
rect 28364 35196 28420 35252
rect 28140 35084 28196 35140
rect 25788 33964 25844 34020
rect 26012 33740 26068 33796
rect 24220 27580 24276 27636
rect 26012 33068 26068 33124
rect 25004 9996 25060 10052
rect 24556 5740 24612 5796
rect 23324 3666 23380 3668
rect 23324 3614 23326 3666
rect 23326 3614 23378 3666
rect 23378 3614 23380 3666
rect 23324 3612 23380 3614
rect 22204 3442 22260 3444
rect 22204 3390 22206 3442
rect 22206 3390 22258 3442
rect 22258 3390 22260 3442
rect 22204 3388 22260 3390
rect 23212 3388 23268 3444
rect 24108 3442 24164 3444
rect 24108 3390 24110 3442
rect 24110 3390 24162 3442
rect 24162 3390 24164 3442
rect 24108 3388 24164 3390
rect 25116 5122 25172 5124
rect 25116 5070 25118 5122
rect 25118 5070 25170 5122
rect 25170 5070 25172 5122
rect 25116 5068 25172 5070
rect 25788 5794 25844 5796
rect 25788 5742 25790 5794
rect 25790 5742 25842 5794
rect 25842 5742 25844 5794
rect 25788 5740 25844 5742
rect 28364 33964 28420 34020
rect 30044 38780 30100 38836
rect 29260 36370 29316 36372
rect 29260 36318 29262 36370
rect 29262 36318 29314 36370
rect 29314 36318 29316 36370
rect 29260 36316 29316 36318
rect 29596 36092 29652 36148
rect 28812 35084 28868 35140
rect 28476 26460 28532 26516
rect 28588 33964 28644 34020
rect 26124 26124 26180 26180
rect 27132 7308 27188 7364
rect 26348 6748 26404 6804
rect 27804 6524 27860 6580
rect 26908 5740 26964 5796
rect 26012 4844 26068 4900
rect 28028 5906 28084 5908
rect 28028 5854 28030 5906
rect 28030 5854 28082 5906
rect 28082 5854 28084 5906
rect 28028 5852 28084 5854
rect 27916 5740 27972 5796
rect 27916 5292 27972 5348
rect 28252 5180 28308 5236
rect 27468 4396 27524 4452
rect 25004 3612 25060 3668
rect 25228 3442 25284 3444
rect 25228 3390 25230 3442
rect 25230 3390 25282 3442
rect 25282 3390 25284 3442
rect 25228 3388 25284 3390
rect 27580 4226 27636 4228
rect 27580 4174 27582 4226
rect 27582 4174 27634 4226
rect 27634 4174 27636 4226
rect 27580 4172 27636 4174
rect 28252 4060 28308 4116
rect 28812 33292 28868 33348
rect 29372 34354 29428 34356
rect 29372 34302 29374 34354
rect 29374 34302 29426 34354
rect 29426 34302 29428 34354
rect 29372 34300 29428 34302
rect 29484 33852 29540 33908
rect 30940 36540 30996 36596
rect 30604 36316 30660 36372
rect 29820 33852 29876 33908
rect 30044 33404 30100 33460
rect 32284 36594 32340 36596
rect 32284 36542 32286 36594
rect 32286 36542 32338 36594
rect 32338 36542 32340 36594
rect 32284 36540 32340 36542
rect 30604 34300 30660 34356
rect 30828 33122 30884 33124
rect 30828 33070 30830 33122
rect 30830 33070 30882 33122
rect 30882 33070 30884 33122
rect 30828 33068 30884 33070
rect 31500 34748 31556 34804
rect 31276 32844 31332 32900
rect 31388 32284 31444 32340
rect 30156 24668 30212 24724
rect 29484 9996 29540 10052
rect 30492 12684 30548 12740
rect 29148 7362 29204 7364
rect 29148 7310 29150 7362
rect 29150 7310 29202 7362
rect 29202 7310 29204 7362
rect 29148 7308 29204 7310
rect 29820 9324 29876 9380
rect 28812 6578 28868 6580
rect 28812 6526 28814 6578
rect 28814 6526 28866 6578
rect 28866 6526 28868 6578
rect 28812 6524 28868 6526
rect 28700 5346 28756 5348
rect 28700 5294 28702 5346
rect 28702 5294 28754 5346
rect 28754 5294 28756 5346
rect 28700 5292 28756 5294
rect 29484 5122 29540 5124
rect 29484 5070 29486 5122
rect 29486 5070 29538 5122
rect 29538 5070 29540 5122
rect 29484 5068 29540 5070
rect 28924 4450 28980 4452
rect 28924 4398 28926 4450
rect 28926 4398 28978 4450
rect 28978 4398 28980 4450
rect 28924 4396 28980 4398
rect 26572 3442 26628 3444
rect 26572 3390 26574 3442
rect 26574 3390 26626 3442
rect 26626 3390 26628 3442
rect 26572 3388 26628 3390
rect 30044 6914 30100 6916
rect 30044 6862 30046 6914
rect 30046 6862 30098 6914
rect 30098 6862 30100 6914
rect 30044 6860 30100 6862
rect 30268 6578 30324 6580
rect 30268 6526 30270 6578
rect 30270 6526 30322 6578
rect 30322 6526 30324 6578
rect 30268 6524 30324 6526
rect 29820 4172 29876 4228
rect 27244 3442 27300 3444
rect 27244 3390 27246 3442
rect 27246 3390 27298 3442
rect 27298 3390 27300 3442
rect 27244 3388 27300 3390
rect 29260 4060 29316 4116
rect 29484 3724 29540 3780
rect 31500 7644 31556 7700
rect 33516 36482 33572 36484
rect 33516 36430 33518 36482
rect 33518 36430 33570 36482
rect 33570 36430 33572 36482
rect 33516 36428 33572 36430
rect 33964 36258 34020 36260
rect 33964 36206 33966 36258
rect 33966 36206 34018 36258
rect 34018 36206 34020 36258
rect 33964 36204 34020 36206
rect 32508 35532 32564 35588
rect 32844 34748 32900 34804
rect 33180 34636 33236 34692
rect 33292 34748 33348 34804
rect 32844 34300 32900 34356
rect 33292 33964 33348 34020
rect 32620 33516 32676 33572
rect 31836 33458 31892 33460
rect 31836 33406 31838 33458
rect 31838 33406 31890 33458
rect 31890 33406 31892 33458
rect 31836 33404 31892 33406
rect 31948 32956 32004 33012
rect 31836 32844 31892 32900
rect 35084 36428 35140 36484
rect 33964 34636 34020 34692
rect 33516 34354 33572 34356
rect 33516 34302 33518 34354
rect 33518 34302 33570 34354
rect 33570 34302 33572 34354
rect 33516 34300 33572 34302
rect 35756 36652 35812 36708
rect 35756 35756 35812 35812
rect 34524 33852 34580 33908
rect 32620 33068 32676 33124
rect 32284 32844 32340 32900
rect 31948 31052 32004 31108
rect 31836 24892 31892 24948
rect 31612 6860 31668 6916
rect 32956 10780 33012 10836
rect 30940 5292 30996 5348
rect 31836 5906 31892 5908
rect 31836 5854 31838 5906
rect 31838 5854 31890 5906
rect 31890 5854 31892 5906
rect 31836 5852 31892 5854
rect 31948 5346 32004 5348
rect 31948 5294 31950 5346
rect 31950 5294 32002 5346
rect 32002 5294 32004 5346
rect 31948 5292 32004 5294
rect 31388 4844 31444 4900
rect 31276 4396 31332 4452
rect 30716 4226 30772 4228
rect 30716 4174 30718 4226
rect 30718 4174 30770 4226
rect 30770 4174 30772 4226
rect 30716 4172 30772 4174
rect 30044 3724 30100 3780
rect 31164 3666 31220 3668
rect 31164 3614 31166 3666
rect 31166 3614 31218 3666
rect 31218 3614 31220 3666
rect 31164 3612 31220 3614
rect 30044 3500 30100 3556
rect 32732 4450 32788 4452
rect 32732 4398 32734 4450
rect 32734 4398 32786 4450
rect 32786 4398 32788 4450
rect 32732 4396 32788 4398
rect 32060 4172 32116 4228
rect 36316 37884 36372 37940
rect 36652 36316 36708 36372
rect 35196 33068 35252 33124
rect 35644 34524 35700 34580
rect 36204 34524 36260 34580
rect 34860 31948 34916 32004
rect 35420 16044 35476 16100
rect 34524 9212 34580 9268
rect 34972 10892 35028 10948
rect 35084 8316 35140 8372
rect 32956 3612 33012 3668
rect 33404 7644 33460 7700
rect 36092 33404 36148 33460
rect 37436 36482 37492 36484
rect 37436 36430 37438 36482
rect 37438 36430 37490 36482
rect 37490 36430 37492 36482
rect 37436 36428 37492 36430
rect 36652 34748 36708 34804
rect 36764 33404 36820 33460
rect 36988 34972 37044 35028
rect 37660 34802 37716 34804
rect 37660 34750 37662 34802
rect 37662 34750 37714 34802
rect 37714 34750 37716 34802
rect 37660 34748 37716 34750
rect 37100 34412 37156 34468
rect 36988 34188 37044 34244
rect 39004 37548 39060 37604
rect 38892 36428 38948 36484
rect 38032 36090 38088 36092
rect 38032 36038 38034 36090
rect 38034 36038 38086 36090
rect 38086 36038 38088 36090
rect 38032 36036 38088 36038
rect 38136 36090 38192 36092
rect 38136 36038 38138 36090
rect 38138 36038 38190 36090
rect 38190 36038 38192 36090
rect 38136 36036 38192 36038
rect 38240 36090 38296 36092
rect 38240 36038 38242 36090
rect 38242 36038 38294 36090
rect 38294 36038 38296 36090
rect 38240 36036 38296 36038
rect 39116 35980 39172 36036
rect 37884 34972 37940 35028
rect 38444 35026 38500 35028
rect 38444 34974 38446 35026
rect 38446 34974 38498 35026
rect 38498 34974 38500 35026
rect 38444 34972 38500 34974
rect 38032 34522 38088 34524
rect 38032 34470 38034 34522
rect 38034 34470 38086 34522
rect 38086 34470 38088 34522
rect 38032 34468 38088 34470
rect 38136 34522 38192 34524
rect 38136 34470 38138 34522
rect 38138 34470 38190 34522
rect 38190 34470 38192 34522
rect 38136 34468 38192 34470
rect 38240 34522 38296 34524
rect 38240 34470 38242 34522
rect 38242 34470 38294 34522
rect 38294 34470 38296 34522
rect 38240 34468 38296 34470
rect 38444 33516 38500 33572
rect 38108 33180 38164 33236
rect 38032 32954 38088 32956
rect 38032 32902 38034 32954
rect 38034 32902 38086 32954
rect 38086 32902 38088 32954
rect 38032 32900 38088 32902
rect 38136 32954 38192 32956
rect 38136 32902 38138 32954
rect 38138 32902 38190 32954
rect 38190 32902 38192 32954
rect 38136 32900 38192 32902
rect 38240 32954 38296 32956
rect 38240 32902 38242 32954
rect 38242 32902 38294 32954
rect 38294 32902 38296 32954
rect 38240 32900 38296 32902
rect 38444 32844 38500 32900
rect 37884 32620 37940 32676
rect 38668 33234 38724 33236
rect 38668 33182 38670 33234
rect 38670 33182 38722 33234
rect 38722 33182 38724 33234
rect 38668 33180 38724 33182
rect 38444 32674 38500 32676
rect 38444 32622 38446 32674
rect 38446 32622 38498 32674
rect 38498 32622 38500 32674
rect 38444 32620 38500 32622
rect 38032 31386 38088 31388
rect 38032 31334 38034 31386
rect 38034 31334 38086 31386
rect 38086 31334 38088 31386
rect 38032 31332 38088 31334
rect 38136 31386 38192 31388
rect 38136 31334 38138 31386
rect 38138 31334 38190 31386
rect 38190 31334 38192 31386
rect 38136 31332 38192 31334
rect 38240 31386 38296 31388
rect 38240 31334 38242 31386
rect 38242 31334 38294 31386
rect 38294 31334 38296 31386
rect 38240 31332 38296 31334
rect 38032 29818 38088 29820
rect 38032 29766 38034 29818
rect 38034 29766 38086 29818
rect 38086 29766 38088 29818
rect 38032 29764 38088 29766
rect 38136 29818 38192 29820
rect 38136 29766 38138 29818
rect 38138 29766 38190 29818
rect 38190 29766 38192 29818
rect 38136 29764 38192 29766
rect 38240 29818 38296 29820
rect 38240 29766 38242 29818
rect 38242 29766 38294 29818
rect 38294 29766 38296 29818
rect 38240 29764 38296 29766
rect 38032 28250 38088 28252
rect 38032 28198 38034 28250
rect 38034 28198 38086 28250
rect 38086 28198 38088 28250
rect 38032 28196 38088 28198
rect 38136 28250 38192 28252
rect 38136 28198 38138 28250
rect 38138 28198 38190 28250
rect 38190 28198 38192 28250
rect 38136 28196 38192 28198
rect 38240 28250 38296 28252
rect 38240 28198 38242 28250
rect 38242 28198 38294 28250
rect 38294 28198 38296 28250
rect 38240 28196 38296 28198
rect 37660 27692 37716 27748
rect 36540 27244 36596 27300
rect 38032 26682 38088 26684
rect 38032 26630 38034 26682
rect 38034 26630 38086 26682
rect 38086 26630 38088 26682
rect 38032 26628 38088 26630
rect 38136 26682 38192 26684
rect 38136 26630 38138 26682
rect 38138 26630 38190 26682
rect 38190 26630 38192 26682
rect 38136 26628 38192 26630
rect 38240 26682 38296 26684
rect 38240 26630 38242 26682
rect 38242 26630 38294 26682
rect 38294 26630 38296 26682
rect 38240 26628 38296 26630
rect 38032 25114 38088 25116
rect 38032 25062 38034 25114
rect 38034 25062 38086 25114
rect 38086 25062 38088 25114
rect 38032 25060 38088 25062
rect 38136 25114 38192 25116
rect 38136 25062 38138 25114
rect 38138 25062 38190 25114
rect 38190 25062 38192 25114
rect 38136 25060 38192 25062
rect 38240 25114 38296 25116
rect 38240 25062 38242 25114
rect 38242 25062 38294 25114
rect 38294 25062 38296 25114
rect 38240 25060 38296 25062
rect 38032 23546 38088 23548
rect 38032 23494 38034 23546
rect 38034 23494 38086 23546
rect 38086 23494 38088 23546
rect 38032 23492 38088 23494
rect 38136 23546 38192 23548
rect 38136 23494 38138 23546
rect 38138 23494 38190 23546
rect 38190 23494 38192 23546
rect 38136 23492 38192 23494
rect 38240 23546 38296 23548
rect 38240 23494 38242 23546
rect 38242 23494 38294 23546
rect 38294 23494 38296 23546
rect 38240 23492 38296 23494
rect 38032 21978 38088 21980
rect 38032 21926 38034 21978
rect 38034 21926 38086 21978
rect 38086 21926 38088 21978
rect 38032 21924 38088 21926
rect 38136 21978 38192 21980
rect 38136 21926 38138 21978
rect 38138 21926 38190 21978
rect 38190 21926 38192 21978
rect 38136 21924 38192 21926
rect 38240 21978 38296 21980
rect 38240 21926 38242 21978
rect 38242 21926 38294 21978
rect 38294 21926 38296 21978
rect 38240 21924 38296 21926
rect 38032 20410 38088 20412
rect 38032 20358 38034 20410
rect 38034 20358 38086 20410
rect 38086 20358 38088 20410
rect 38032 20356 38088 20358
rect 38136 20410 38192 20412
rect 38136 20358 38138 20410
rect 38138 20358 38190 20410
rect 38190 20358 38192 20410
rect 38136 20356 38192 20358
rect 38240 20410 38296 20412
rect 38240 20358 38242 20410
rect 38242 20358 38294 20410
rect 38294 20358 38296 20410
rect 38240 20356 38296 20358
rect 38032 18842 38088 18844
rect 38032 18790 38034 18842
rect 38034 18790 38086 18842
rect 38086 18790 38088 18842
rect 38032 18788 38088 18790
rect 38136 18842 38192 18844
rect 38136 18790 38138 18842
rect 38138 18790 38190 18842
rect 38190 18790 38192 18842
rect 38136 18788 38192 18790
rect 38240 18842 38296 18844
rect 38240 18790 38242 18842
rect 38242 18790 38294 18842
rect 38294 18790 38296 18842
rect 38240 18788 38296 18790
rect 38032 17274 38088 17276
rect 38032 17222 38034 17274
rect 38034 17222 38086 17274
rect 38086 17222 38088 17274
rect 38032 17220 38088 17222
rect 38136 17274 38192 17276
rect 38136 17222 38138 17274
rect 38138 17222 38190 17274
rect 38190 17222 38192 17274
rect 38136 17220 38192 17222
rect 38240 17274 38296 17276
rect 38240 17222 38242 17274
rect 38242 17222 38294 17274
rect 38294 17222 38296 17274
rect 38240 17220 38296 17222
rect 38032 15706 38088 15708
rect 38032 15654 38034 15706
rect 38034 15654 38086 15706
rect 38086 15654 38088 15706
rect 38032 15652 38088 15654
rect 38136 15706 38192 15708
rect 38136 15654 38138 15706
rect 38138 15654 38190 15706
rect 38190 15654 38192 15706
rect 38136 15652 38192 15654
rect 38240 15706 38296 15708
rect 38240 15654 38242 15706
rect 38242 15654 38294 15706
rect 38294 15654 38296 15706
rect 38240 15652 38296 15654
rect 39340 35810 39396 35812
rect 39340 35758 39342 35810
rect 39342 35758 39394 35810
rect 39394 35758 39396 35810
rect 39340 35756 39396 35758
rect 39004 32844 39060 32900
rect 39004 32562 39060 32564
rect 39004 32510 39006 32562
rect 39006 32510 39058 32562
rect 39058 32510 39060 32562
rect 39004 32508 39060 32510
rect 39228 32844 39284 32900
rect 39452 34972 39508 35028
rect 40348 36428 40404 36484
rect 41132 36258 41188 36260
rect 41132 36206 41134 36258
rect 41134 36206 41186 36258
rect 41186 36206 41188 36258
rect 41132 36204 41188 36206
rect 40012 35474 40068 35476
rect 40012 35422 40014 35474
rect 40014 35422 40066 35474
rect 40066 35422 40068 35474
rect 40012 35420 40068 35422
rect 39788 34860 39844 34916
rect 39564 32284 39620 32340
rect 39900 34188 39956 34244
rect 39116 27804 39172 27860
rect 38444 15036 38500 15092
rect 38032 14138 38088 14140
rect 38032 14086 38034 14138
rect 38034 14086 38086 14138
rect 38086 14086 38088 14138
rect 38032 14084 38088 14086
rect 38136 14138 38192 14140
rect 38136 14086 38138 14138
rect 38138 14086 38190 14138
rect 38190 14086 38192 14138
rect 38136 14084 38192 14086
rect 38240 14138 38296 14140
rect 38240 14086 38242 14138
rect 38242 14086 38294 14138
rect 38294 14086 38296 14138
rect 38240 14084 38296 14086
rect 38032 12570 38088 12572
rect 38032 12518 38034 12570
rect 38034 12518 38086 12570
rect 38086 12518 38088 12570
rect 38032 12516 38088 12518
rect 38136 12570 38192 12572
rect 38136 12518 38138 12570
rect 38138 12518 38190 12570
rect 38190 12518 38192 12570
rect 38136 12516 38192 12518
rect 38240 12570 38296 12572
rect 38240 12518 38242 12570
rect 38242 12518 38294 12570
rect 38294 12518 38296 12570
rect 38240 12516 38296 12518
rect 38032 11002 38088 11004
rect 38032 10950 38034 11002
rect 38034 10950 38086 11002
rect 38086 10950 38088 11002
rect 38032 10948 38088 10950
rect 38136 11002 38192 11004
rect 38136 10950 38138 11002
rect 38138 10950 38190 11002
rect 38190 10950 38192 11002
rect 38136 10948 38192 10950
rect 38240 11002 38296 11004
rect 38240 10950 38242 11002
rect 38242 10950 38294 11002
rect 38294 10950 38296 11002
rect 38240 10948 38296 10950
rect 35644 9324 35700 9380
rect 38032 9434 38088 9436
rect 38032 9382 38034 9434
rect 38034 9382 38086 9434
rect 38086 9382 38088 9434
rect 38032 9380 38088 9382
rect 38136 9434 38192 9436
rect 38136 9382 38138 9434
rect 38138 9382 38190 9434
rect 38190 9382 38192 9434
rect 38136 9380 38192 9382
rect 38240 9434 38296 9436
rect 38240 9382 38242 9434
rect 38242 9382 38294 9434
rect 38294 9382 38296 9434
rect 38240 9380 38296 9382
rect 38032 7866 38088 7868
rect 38032 7814 38034 7866
rect 38034 7814 38086 7866
rect 38086 7814 38088 7866
rect 38032 7812 38088 7814
rect 38136 7866 38192 7868
rect 38136 7814 38138 7866
rect 38138 7814 38190 7866
rect 38190 7814 38192 7866
rect 38136 7812 38192 7814
rect 38240 7866 38296 7868
rect 38240 7814 38242 7866
rect 38242 7814 38294 7866
rect 38294 7814 38296 7866
rect 38240 7812 38296 7814
rect 37884 7308 37940 7364
rect 37436 6524 37492 6580
rect 36764 5964 36820 6020
rect 37436 5964 37492 6020
rect 35532 5068 35588 5124
rect 33516 4450 33572 4452
rect 33516 4398 33518 4450
rect 33518 4398 33570 4450
rect 33570 4398 33572 4450
rect 33516 4396 33572 4398
rect 33404 3612 33460 3668
rect 34860 3666 34916 3668
rect 34860 3614 34862 3666
rect 34862 3614 34914 3666
rect 34914 3614 34916 3666
rect 34860 3612 34916 3614
rect 35532 3612 35588 3668
rect 36764 5628 36820 5684
rect 40124 31836 40180 31892
rect 39900 12684 39956 12740
rect 39228 7362 39284 7364
rect 39228 7310 39230 7362
rect 39230 7310 39282 7362
rect 39282 7310 39284 7362
rect 39228 7308 39284 7310
rect 39116 6802 39172 6804
rect 39116 6750 39118 6802
rect 39118 6750 39170 6802
rect 39170 6750 39172 6802
rect 39116 6748 39172 6750
rect 38332 6578 38388 6580
rect 38332 6526 38334 6578
rect 38334 6526 38386 6578
rect 38386 6526 38388 6578
rect 38332 6524 38388 6526
rect 38892 6412 38948 6468
rect 38032 6298 38088 6300
rect 38032 6246 38034 6298
rect 38034 6246 38086 6298
rect 38086 6246 38088 6298
rect 38032 6244 38088 6246
rect 38136 6298 38192 6300
rect 38136 6246 38138 6298
rect 38138 6246 38190 6298
rect 38190 6246 38192 6298
rect 38136 6244 38192 6246
rect 38240 6298 38296 6300
rect 38240 6246 38242 6298
rect 38242 6246 38294 6298
rect 38294 6246 38296 6298
rect 38240 6244 38296 6246
rect 37548 5682 37604 5684
rect 37548 5630 37550 5682
rect 37550 5630 37602 5682
rect 37602 5630 37604 5682
rect 37548 5628 37604 5630
rect 38220 5628 38276 5684
rect 38032 4730 38088 4732
rect 38032 4678 38034 4730
rect 38034 4678 38086 4730
rect 38086 4678 38088 4730
rect 38032 4676 38088 4678
rect 38136 4730 38192 4732
rect 38136 4678 38138 4730
rect 38138 4678 38190 4730
rect 38190 4678 38192 4730
rect 38136 4676 38192 4678
rect 38240 4730 38296 4732
rect 38240 4678 38242 4730
rect 38242 4678 38294 4730
rect 38294 4678 38296 4730
rect 38240 4676 38296 4678
rect 41580 35308 41636 35364
rect 40460 34242 40516 34244
rect 40460 34190 40462 34242
rect 40462 34190 40514 34242
rect 40514 34190 40516 34242
rect 40460 34188 40516 34190
rect 40796 34076 40852 34132
rect 41580 33740 41636 33796
rect 41020 33628 41076 33684
rect 40460 32732 40516 32788
rect 40796 32562 40852 32564
rect 40796 32510 40798 32562
rect 40798 32510 40850 32562
rect 40850 32510 40852 32562
rect 40796 32508 40852 32510
rect 40908 29260 40964 29316
rect 41244 32732 41300 32788
rect 40124 6802 40180 6804
rect 40124 6750 40126 6802
rect 40126 6750 40178 6802
rect 40178 6750 40180 6802
rect 40124 6748 40180 6750
rect 40572 10892 40628 10948
rect 41804 33628 41860 33684
rect 43036 37996 43092 38052
rect 41916 33516 41972 33572
rect 42028 35420 42084 35476
rect 42140 33740 42196 33796
rect 42028 24780 42084 24836
rect 42140 33516 42196 33572
rect 42364 33516 42420 33572
rect 42364 33068 42420 33124
rect 42140 32956 42196 33012
rect 43932 38668 43988 38724
rect 42812 35084 42868 35140
rect 43148 35084 43204 35140
rect 44604 37212 44660 37268
rect 45276 36988 45332 37044
rect 45276 36370 45332 36372
rect 45276 36318 45278 36370
rect 45278 36318 45330 36370
rect 45330 36318 45332 36370
rect 45276 36316 45332 36318
rect 44716 36092 44772 36148
rect 44716 34636 44772 34692
rect 45724 35980 45780 36036
rect 45836 36204 45892 36260
rect 45612 34914 45668 34916
rect 45612 34862 45614 34914
rect 45614 34862 45666 34914
rect 45666 34862 45668 34914
rect 45612 34860 45668 34862
rect 44604 34076 44660 34132
rect 43596 33740 43652 33796
rect 43148 33628 43204 33684
rect 44604 31164 44660 31220
rect 45052 31836 45108 31892
rect 42476 27132 42532 27188
rect 42812 27692 42868 27748
rect 42140 13356 42196 13412
rect 41244 10780 41300 10836
rect 40572 8316 40628 8372
rect 39788 6412 39844 6468
rect 40460 6466 40516 6468
rect 40460 6414 40462 6466
rect 40462 6414 40514 6466
rect 40514 6414 40516 6466
rect 40460 6412 40516 6414
rect 39676 6018 39732 6020
rect 39676 5966 39678 6018
rect 39678 5966 39730 6018
rect 39730 5966 39732 6018
rect 39676 5964 39732 5966
rect 40460 5964 40516 6020
rect 40236 5794 40292 5796
rect 40236 5742 40238 5794
rect 40238 5742 40290 5794
rect 40290 5742 40292 5794
rect 40236 5740 40292 5742
rect 40348 5682 40404 5684
rect 40348 5630 40350 5682
rect 40350 5630 40402 5682
rect 40402 5630 40404 5682
rect 40348 5628 40404 5630
rect 38444 4508 38500 4564
rect 38556 5068 38612 5124
rect 39116 4562 39172 4564
rect 39116 4510 39118 4562
rect 39118 4510 39170 4562
rect 39170 4510 39172 4562
rect 39116 4508 39172 4510
rect 39564 4508 39620 4564
rect 40236 4284 40292 4340
rect 39340 4172 39396 4228
rect 36204 3442 36260 3444
rect 36204 3390 36206 3442
rect 36206 3390 36258 3442
rect 36258 3390 36260 3442
rect 36204 3388 36260 3390
rect 36876 3388 36932 3444
rect 37772 3442 37828 3444
rect 37772 3390 37774 3442
rect 37774 3390 37826 3442
rect 37826 3390 37828 3442
rect 37772 3388 37828 3390
rect 38332 3442 38388 3444
rect 38332 3390 38334 3442
rect 38334 3390 38386 3442
rect 38386 3390 38388 3442
rect 38332 3388 38388 3390
rect 38032 3162 38088 3164
rect 38032 3110 38034 3162
rect 38034 3110 38086 3162
rect 38086 3110 38088 3162
rect 38032 3108 38088 3110
rect 38136 3162 38192 3164
rect 38136 3110 38138 3162
rect 38138 3110 38190 3162
rect 38190 3110 38192 3162
rect 38136 3108 38192 3110
rect 38240 3162 38296 3164
rect 38240 3110 38242 3162
rect 38242 3110 38294 3162
rect 38294 3110 38296 3162
rect 38240 3108 38296 3110
rect 39676 3724 39732 3780
rect 40348 4226 40404 4228
rect 40348 4174 40350 4226
rect 40350 4174 40402 4226
rect 40402 4174 40404 4226
rect 40348 4172 40404 4174
rect 41020 5852 41076 5908
rect 40908 5794 40964 5796
rect 40908 5742 40910 5794
rect 40910 5742 40962 5794
rect 40962 5742 40964 5794
rect 40908 5740 40964 5742
rect 40908 5180 40964 5236
rect 41468 5906 41524 5908
rect 41468 5854 41470 5906
rect 41470 5854 41522 5906
rect 41522 5854 41524 5906
rect 41468 5852 41524 5854
rect 41692 5234 41748 5236
rect 41692 5182 41694 5234
rect 41694 5182 41746 5234
rect 41746 5182 41748 5234
rect 41692 5180 41748 5182
rect 41580 5122 41636 5124
rect 41580 5070 41582 5122
rect 41582 5070 41634 5122
rect 41634 5070 41636 5122
rect 41580 5068 41636 5070
rect 42252 5122 42308 5124
rect 42252 5070 42254 5122
rect 42254 5070 42306 5122
rect 42306 5070 42308 5122
rect 42252 5068 42308 5070
rect 40572 3724 40628 3780
rect 40236 3666 40292 3668
rect 40236 3614 40238 3666
rect 40238 3614 40290 3666
rect 40290 3614 40292 3666
rect 40236 3612 40292 3614
rect 40684 3388 40740 3444
rect 41244 3442 41300 3444
rect 41244 3390 41246 3442
rect 41246 3390 41298 3442
rect 41298 3390 41300 3442
rect 41244 3388 41300 3390
rect 45052 23324 45108 23380
rect 43932 15036 43988 15092
rect 41692 3388 41748 3444
rect 44604 5404 44660 5460
rect 44716 4956 44772 5012
rect 45388 33068 45444 33124
rect 45388 31724 45444 31780
rect 46844 36370 46900 36372
rect 46844 36318 46846 36370
rect 46846 36318 46898 36370
rect 46898 36318 46900 36370
rect 46844 36316 46900 36318
rect 46060 34300 46116 34356
rect 46284 36092 46340 36148
rect 46396 35308 46452 35364
rect 46396 34412 46452 34468
rect 45836 22988 45892 23044
rect 47404 36540 47460 36596
rect 47068 34636 47124 34692
rect 45724 20076 45780 20132
rect 45276 16044 45332 16100
rect 46956 32060 47012 32116
rect 47180 28028 47236 28084
rect 47292 34860 47348 34916
rect 48076 36594 48132 36596
rect 48076 36542 48078 36594
rect 48078 36542 48130 36594
rect 48130 36542 48132 36594
rect 48076 36540 48132 36542
rect 47628 36316 47684 36372
rect 47516 34972 47572 35028
rect 47404 34636 47460 34692
rect 48412 35922 48468 35924
rect 48412 35870 48414 35922
rect 48414 35870 48466 35922
rect 48466 35870 48468 35922
rect 48412 35868 48468 35870
rect 48300 34972 48356 35028
rect 47852 34914 47908 34916
rect 47852 34862 47854 34914
rect 47854 34862 47906 34914
rect 47906 34862 47908 34914
rect 47852 34860 47908 34862
rect 47292 26348 47348 26404
rect 46508 14364 46564 14420
rect 46732 13356 46788 13412
rect 45276 4956 45332 5012
rect 45612 5010 45668 5012
rect 45612 4958 45614 5010
rect 45614 4958 45666 5010
rect 45666 4958 45668 5010
rect 45612 4956 45668 4958
rect 45052 4172 45108 4228
rect 45276 4338 45332 4340
rect 45276 4286 45278 4338
rect 45278 4286 45330 4338
rect 45330 4286 45332 4338
rect 45276 4284 45332 4286
rect 47068 9212 47124 9268
rect 46956 6018 47012 6020
rect 46956 5966 46958 6018
rect 46958 5966 47010 6018
rect 47010 5966 47012 6018
rect 46956 5964 47012 5966
rect 48188 34300 48244 34356
rect 49532 36652 49588 36708
rect 49196 36482 49252 36484
rect 49196 36430 49198 36482
rect 49198 36430 49250 36482
rect 49250 36430 49252 36482
rect 49196 36428 49252 36430
rect 48748 35698 48804 35700
rect 48748 35646 48750 35698
rect 48750 35646 48802 35698
rect 48802 35646 48804 35698
rect 48748 35644 48804 35646
rect 48748 34354 48804 34356
rect 48748 34302 48750 34354
rect 48750 34302 48802 34354
rect 48802 34302 48804 34354
rect 48748 34300 48804 34302
rect 48524 34188 48580 34244
rect 49644 36204 49700 36260
rect 49980 36258 50036 36260
rect 49980 36206 49982 36258
rect 49982 36206 50034 36258
rect 50034 36206 50036 36258
rect 49980 36204 50036 36206
rect 49532 34860 49588 34916
rect 48972 34636 49028 34692
rect 49644 34242 49700 34244
rect 49644 34190 49646 34242
rect 49646 34190 49698 34242
rect 49698 34190 49700 34242
rect 49644 34188 49700 34190
rect 47964 33516 48020 33572
rect 48860 33292 48916 33348
rect 48524 32562 48580 32564
rect 48524 32510 48526 32562
rect 48526 32510 48578 32562
rect 48578 32510 48580 32562
rect 48524 32508 48580 32510
rect 49756 33852 49812 33908
rect 49196 33234 49252 33236
rect 49196 33182 49198 33234
rect 49198 33182 49250 33234
rect 49250 33182 49252 33234
rect 49196 33180 49252 33182
rect 49420 33180 49476 33236
rect 49868 33122 49924 33124
rect 49868 33070 49870 33122
rect 49870 33070 49922 33122
rect 49922 33070 49924 33122
rect 49868 33068 49924 33070
rect 50204 35420 50260 35476
rect 49196 23436 49252 23492
rect 48972 16828 49028 16884
rect 47852 7420 47908 7476
rect 48748 7474 48804 7476
rect 48748 7422 48750 7474
rect 48750 7422 48802 7474
rect 48802 7422 48804 7474
rect 48748 7420 48804 7422
rect 50988 36428 51044 36484
rect 51548 36204 51604 36260
rect 51100 35980 51156 36036
rect 50316 34972 50372 35028
rect 50428 35532 50484 35588
rect 50876 35026 50932 35028
rect 50876 34974 50878 35026
rect 50878 34974 50930 35026
rect 50930 34974 50932 35026
rect 50876 34972 50932 34974
rect 50428 34860 50484 34916
rect 50764 34188 50820 34244
rect 50764 33852 50820 33908
rect 51436 33740 51492 33796
rect 51324 33516 51380 33572
rect 51212 33404 51268 33460
rect 51660 35474 51716 35476
rect 51660 35422 51662 35474
rect 51662 35422 51714 35474
rect 51714 35422 51716 35474
rect 51660 35420 51716 35422
rect 51772 33740 51828 33796
rect 51548 32844 51604 32900
rect 51996 34748 52052 34804
rect 51996 32844 52052 32900
rect 51884 31724 51940 31780
rect 51660 27916 51716 27972
rect 52220 35810 52276 35812
rect 52220 35758 52222 35810
rect 52222 35758 52274 35810
rect 52274 35758 52276 35810
rect 52220 35756 52276 35758
rect 52892 36316 52948 36372
rect 52780 35868 52836 35924
rect 52668 35756 52724 35812
rect 52108 24556 52164 24612
rect 52444 33740 52500 33796
rect 53116 36482 53172 36484
rect 53116 36430 53118 36482
rect 53118 36430 53170 36482
rect 53170 36430 53172 36482
rect 53116 36428 53172 36430
rect 52892 34524 52948 34580
rect 52556 33516 52612 33572
rect 53564 35084 53620 35140
rect 54796 36428 54852 36484
rect 56252 38108 56308 38164
rect 54572 35644 54628 35700
rect 53564 33404 53620 33460
rect 52556 31724 52612 31780
rect 52444 22876 52500 22932
rect 52892 23436 52948 23492
rect 51324 17612 51380 17668
rect 51436 16828 51492 16884
rect 50316 8428 50372 8484
rect 50316 7586 50372 7588
rect 50316 7534 50318 7586
rect 50318 7534 50370 7586
rect 50370 7534 50372 7586
rect 50316 7532 50372 7534
rect 50092 7420 50148 7476
rect 49756 7196 49812 7252
rect 50540 7196 50596 7252
rect 51100 7196 51156 7252
rect 48300 6636 48356 6692
rect 49532 6690 49588 6692
rect 49532 6638 49534 6690
rect 49534 6638 49586 6690
rect 49586 6638 49588 6690
rect 49532 6636 49588 6638
rect 48076 6412 48132 6468
rect 47516 5964 47572 6020
rect 46732 3612 46788 3668
rect 45276 3388 45332 3444
rect 48748 5906 48804 5908
rect 48748 5854 48750 5906
rect 48750 5854 48802 5906
rect 48802 5854 48804 5906
rect 48748 5852 48804 5854
rect 49084 5852 49140 5908
rect 48412 5404 48468 5460
rect 48860 5404 48916 5460
rect 48076 5122 48132 5124
rect 48076 5070 48078 5122
rect 48078 5070 48130 5122
rect 48130 5070 48132 5122
rect 48076 5068 48132 5070
rect 48636 5122 48692 5124
rect 48636 5070 48638 5122
rect 48638 5070 48690 5122
rect 48690 5070 48692 5122
rect 48636 5068 48692 5070
rect 49420 5852 49476 5908
rect 50540 6578 50596 6580
rect 50540 6526 50542 6578
rect 50542 6526 50594 6578
rect 50594 6526 50596 6578
rect 50540 6524 50596 6526
rect 49756 6076 49812 6132
rect 50316 6412 50372 6468
rect 51100 6130 51156 6132
rect 51100 6078 51102 6130
rect 51102 6078 51154 6130
rect 51154 6078 51156 6130
rect 51100 6076 51156 6078
rect 49868 5068 49924 5124
rect 47516 3666 47572 3668
rect 47516 3614 47518 3666
rect 47518 3614 47570 3666
rect 47570 3614 47572 3666
rect 47516 3612 47572 3614
rect 48860 3442 48916 3444
rect 48860 3390 48862 3442
rect 48862 3390 48914 3442
rect 48914 3390 48916 3442
rect 48860 3388 48916 3390
rect 50764 4226 50820 4228
rect 50764 4174 50766 4226
rect 50766 4174 50818 4226
rect 50818 4174 50820 4226
rect 50764 4172 50820 4174
rect 51548 7474 51604 7476
rect 51548 7422 51550 7474
rect 51550 7422 51602 7474
rect 51602 7422 51604 7474
rect 51548 7420 51604 7422
rect 52108 6578 52164 6580
rect 52108 6526 52110 6578
rect 52110 6526 52162 6578
rect 52162 6526 52164 6578
rect 52108 6524 52164 6526
rect 51548 6466 51604 6468
rect 51548 6414 51550 6466
rect 51550 6414 51602 6466
rect 51602 6414 51604 6466
rect 51548 6412 51604 6414
rect 52892 5906 52948 5908
rect 52892 5854 52894 5906
rect 52894 5854 52946 5906
rect 52946 5854 52948 5906
rect 52892 5852 52948 5854
rect 52556 5740 52612 5796
rect 52556 5180 52612 5236
rect 54124 34242 54180 34244
rect 54124 34190 54126 34242
rect 54126 34190 54178 34242
rect 54178 34190 54180 34242
rect 54124 34188 54180 34190
rect 53900 33458 53956 33460
rect 53900 33406 53902 33458
rect 53902 33406 53954 33458
rect 53954 33406 53956 33458
rect 53900 33404 53956 33406
rect 53676 12796 53732 12852
rect 54236 32060 54292 32116
rect 53340 5906 53396 5908
rect 53340 5854 53342 5906
rect 53342 5854 53394 5906
rect 53394 5854 53396 5906
rect 53340 5852 53396 5854
rect 53564 5292 53620 5348
rect 54124 5292 54180 5348
rect 53452 5122 53508 5124
rect 53452 5070 53454 5122
rect 53454 5070 53506 5122
rect 53506 5070 53508 5122
rect 53452 5068 53508 5070
rect 54124 5068 54180 5124
rect 53004 4956 53060 5012
rect 55356 34914 55412 34916
rect 55356 34862 55358 34914
rect 55358 34862 55410 34914
rect 55410 34862 55412 34914
rect 55356 34860 55412 34862
rect 54572 34188 54628 34244
rect 54348 22540 54404 22596
rect 56442 36874 56498 36876
rect 56442 36822 56444 36874
rect 56444 36822 56496 36874
rect 56496 36822 56498 36874
rect 56442 36820 56498 36822
rect 56546 36874 56602 36876
rect 56546 36822 56548 36874
rect 56548 36822 56600 36874
rect 56600 36822 56602 36874
rect 56546 36820 56602 36822
rect 56650 36874 56706 36876
rect 56650 36822 56652 36874
rect 56652 36822 56704 36874
rect 56704 36822 56706 36874
rect 56650 36820 56706 36822
rect 56812 35756 56868 35812
rect 56442 35306 56498 35308
rect 56442 35254 56444 35306
rect 56444 35254 56496 35306
rect 56496 35254 56498 35306
rect 56442 35252 56498 35254
rect 56546 35306 56602 35308
rect 56546 35254 56548 35306
rect 56548 35254 56600 35306
rect 56600 35254 56602 35306
rect 56546 35252 56602 35254
rect 56650 35306 56706 35308
rect 56650 35254 56652 35306
rect 56652 35254 56704 35306
rect 56704 35254 56706 35306
rect 56650 35252 56706 35254
rect 56700 34802 56756 34804
rect 56700 34750 56702 34802
rect 56702 34750 56754 34802
rect 56754 34750 56756 34802
rect 56700 34748 56756 34750
rect 56252 34690 56308 34692
rect 56252 34638 56254 34690
rect 56254 34638 56306 34690
rect 56306 34638 56308 34690
rect 56252 34636 56308 34638
rect 57036 35196 57092 35252
rect 57036 34636 57092 34692
rect 56442 33738 56498 33740
rect 56442 33686 56444 33738
rect 56444 33686 56496 33738
rect 56496 33686 56498 33738
rect 56442 33684 56498 33686
rect 56546 33738 56602 33740
rect 56546 33686 56548 33738
rect 56548 33686 56600 33738
rect 56600 33686 56602 33738
rect 56546 33684 56602 33686
rect 56650 33738 56706 33740
rect 56650 33686 56652 33738
rect 56652 33686 56704 33738
rect 56704 33686 56706 33738
rect 56650 33684 56706 33686
rect 56442 32170 56498 32172
rect 56442 32118 56444 32170
rect 56444 32118 56496 32170
rect 56496 32118 56498 32170
rect 56442 32116 56498 32118
rect 56546 32170 56602 32172
rect 56546 32118 56548 32170
rect 56548 32118 56600 32170
rect 56600 32118 56602 32170
rect 56546 32116 56602 32118
rect 56650 32170 56706 32172
rect 56650 32118 56652 32170
rect 56652 32118 56704 32170
rect 56704 32118 56706 32170
rect 56650 32116 56706 32118
rect 56442 30602 56498 30604
rect 56442 30550 56444 30602
rect 56444 30550 56496 30602
rect 56496 30550 56498 30602
rect 56442 30548 56498 30550
rect 56546 30602 56602 30604
rect 56546 30550 56548 30602
rect 56548 30550 56600 30602
rect 56600 30550 56602 30602
rect 56546 30548 56602 30550
rect 56650 30602 56706 30604
rect 56650 30550 56652 30602
rect 56652 30550 56704 30602
rect 56704 30550 56706 30602
rect 56650 30548 56706 30550
rect 56442 29034 56498 29036
rect 56442 28982 56444 29034
rect 56444 28982 56496 29034
rect 56496 28982 56498 29034
rect 56442 28980 56498 28982
rect 56546 29034 56602 29036
rect 56546 28982 56548 29034
rect 56548 28982 56600 29034
rect 56600 28982 56602 29034
rect 56546 28980 56602 28982
rect 56650 29034 56706 29036
rect 56650 28982 56652 29034
rect 56652 28982 56704 29034
rect 56704 28982 56706 29034
rect 56650 28980 56706 28982
rect 56442 27466 56498 27468
rect 56442 27414 56444 27466
rect 56444 27414 56496 27466
rect 56496 27414 56498 27466
rect 56442 27412 56498 27414
rect 56546 27466 56602 27468
rect 56546 27414 56548 27466
rect 56548 27414 56600 27466
rect 56600 27414 56602 27466
rect 56546 27412 56602 27414
rect 56650 27466 56706 27468
rect 56650 27414 56652 27466
rect 56652 27414 56704 27466
rect 56704 27414 56706 27466
rect 56650 27412 56706 27414
rect 56442 25898 56498 25900
rect 56442 25846 56444 25898
rect 56444 25846 56496 25898
rect 56496 25846 56498 25898
rect 56442 25844 56498 25846
rect 56546 25898 56602 25900
rect 56546 25846 56548 25898
rect 56548 25846 56600 25898
rect 56600 25846 56602 25898
rect 56546 25844 56602 25846
rect 56650 25898 56706 25900
rect 56650 25846 56652 25898
rect 56652 25846 56704 25898
rect 56704 25846 56706 25898
rect 56650 25844 56706 25846
rect 55692 25676 55748 25732
rect 56442 24330 56498 24332
rect 56442 24278 56444 24330
rect 56444 24278 56496 24330
rect 56496 24278 56498 24330
rect 56442 24276 56498 24278
rect 56546 24330 56602 24332
rect 56546 24278 56548 24330
rect 56548 24278 56600 24330
rect 56600 24278 56602 24330
rect 56546 24276 56602 24278
rect 56650 24330 56706 24332
rect 56650 24278 56652 24330
rect 56652 24278 56704 24330
rect 56704 24278 56706 24330
rect 56650 24276 56706 24278
rect 56442 22762 56498 22764
rect 56442 22710 56444 22762
rect 56444 22710 56496 22762
rect 56496 22710 56498 22762
rect 56442 22708 56498 22710
rect 56546 22762 56602 22764
rect 56546 22710 56548 22762
rect 56548 22710 56600 22762
rect 56600 22710 56602 22762
rect 56546 22708 56602 22710
rect 56650 22762 56706 22764
rect 56650 22710 56652 22762
rect 56652 22710 56704 22762
rect 56704 22710 56706 22762
rect 56650 22708 56706 22710
rect 54908 21308 54964 21364
rect 56442 21194 56498 21196
rect 56442 21142 56444 21194
rect 56444 21142 56496 21194
rect 56496 21142 56498 21194
rect 56442 21140 56498 21142
rect 56546 21194 56602 21196
rect 56546 21142 56548 21194
rect 56548 21142 56600 21194
rect 56600 21142 56602 21194
rect 56546 21140 56602 21142
rect 56650 21194 56706 21196
rect 56650 21142 56652 21194
rect 56652 21142 56704 21194
rect 56704 21142 56706 21194
rect 56650 21140 56706 21142
rect 56442 19626 56498 19628
rect 56442 19574 56444 19626
rect 56444 19574 56496 19626
rect 56496 19574 56498 19626
rect 56442 19572 56498 19574
rect 56546 19626 56602 19628
rect 56546 19574 56548 19626
rect 56548 19574 56600 19626
rect 56600 19574 56602 19626
rect 56546 19572 56602 19574
rect 56650 19626 56706 19628
rect 56650 19574 56652 19626
rect 56652 19574 56704 19626
rect 56704 19574 56706 19626
rect 56650 19572 56706 19574
rect 56442 18058 56498 18060
rect 56442 18006 56444 18058
rect 56444 18006 56496 18058
rect 56496 18006 56498 18058
rect 56442 18004 56498 18006
rect 56546 18058 56602 18060
rect 56546 18006 56548 18058
rect 56548 18006 56600 18058
rect 56600 18006 56602 18058
rect 56546 18004 56602 18006
rect 56650 18058 56706 18060
rect 56650 18006 56652 18058
rect 56652 18006 56704 18058
rect 56704 18006 56706 18058
rect 56650 18004 56706 18006
rect 57596 35810 57652 35812
rect 57596 35758 57598 35810
rect 57598 35758 57650 35810
rect 57650 35758 57652 35810
rect 57596 35756 57652 35758
rect 57484 34354 57540 34356
rect 57484 34302 57486 34354
rect 57486 34302 57538 34354
rect 57538 34302 57540 34354
rect 57484 34300 57540 34302
rect 57148 32732 57204 32788
rect 57036 17612 57092 17668
rect 56442 16490 56498 16492
rect 56442 16438 56444 16490
rect 56444 16438 56496 16490
rect 56496 16438 56498 16490
rect 56442 16436 56498 16438
rect 56546 16490 56602 16492
rect 56546 16438 56548 16490
rect 56548 16438 56600 16490
rect 56600 16438 56602 16490
rect 56546 16436 56602 16438
rect 56650 16490 56706 16492
rect 56650 16438 56652 16490
rect 56652 16438 56704 16490
rect 56704 16438 56706 16490
rect 56650 16436 56706 16438
rect 56442 14922 56498 14924
rect 56442 14870 56444 14922
rect 56444 14870 56496 14922
rect 56496 14870 56498 14922
rect 56442 14868 56498 14870
rect 56546 14922 56602 14924
rect 56546 14870 56548 14922
rect 56548 14870 56600 14922
rect 56600 14870 56602 14922
rect 56546 14868 56602 14870
rect 56650 14922 56706 14924
rect 56650 14870 56652 14922
rect 56652 14870 56704 14922
rect 56704 14870 56706 14922
rect 56650 14868 56706 14870
rect 58268 33964 58324 34020
rect 59500 36092 59556 36148
rect 58604 33964 58660 34020
rect 58492 33740 58548 33796
rect 58716 33516 58772 33572
rect 57932 26236 57988 26292
rect 58828 32508 58884 32564
rect 58604 23100 58660 23156
rect 58940 31612 58996 31668
rect 59500 34748 59556 34804
rect 59500 33852 59556 33908
rect 59612 33740 59668 33796
rect 59164 33516 59220 33572
rect 59052 30156 59108 30212
rect 60844 36370 60900 36372
rect 60844 36318 60846 36370
rect 60846 36318 60898 36370
rect 60898 36318 60900 36370
rect 60844 36316 60900 36318
rect 59836 34748 59892 34804
rect 59724 26796 59780 26852
rect 61292 34860 61348 34916
rect 57820 14252 57876 14308
rect 58044 14364 58100 14420
rect 56442 13354 56498 13356
rect 56442 13302 56444 13354
rect 56444 13302 56496 13354
rect 56496 13302 56498 13354
rect 56442 13300 56498 13302
rect 56546 13354 56602 13356
rect 56546 13302 56548 13354
rect 56548 13302 56600 13354
rect 56600 13302 56602 13354
rect 56546 13300 56602 13302
rect 56650 13354 56706 13356
rect 56650 13302 56652 13354
rect 56652 13302 56704 13354
rect 56704 13302 56706 13354
rect 56650 13300 56706 13302
rect 56442 11786 56498 11788
rect 56442 11734 56444 11786
rect 56444 11734 56496 11786
rect 56496 11734 56498 11786
rect 56442 11732 56498 11734
rect 56546 11786 56602 11788
rect 56546 11734 56548 11786
rect 56548 11734 56600 11786
rect 56600 11734 56602 11786
rect 56546 11732 56602 11734
rect 56650 11786 56706 11788
rect 56650 11734 56652 11786
rect 56652 11734 56704 11786
rect 56704 11734 56706 11786
rect 56650 11732 56706 11734
rect 56442 10218 56498 10220
rect 56442 10166 56444 10218
rect 56444 10166 56496 10218
rect 56496 10166 56498 10218
rect 56442 10164 56498 10166
rect 56546 10218 56602 10220
rect 56546 10166 56548 10218
rect 56548 10166 56600 10218
rect 56600 10166 56602 10218
rect 56546 10164 56602 10166
rect 56650 10218 56706 10220
rect 56650 10166 56652 10218
rect 56652 10166 56704 10218
rect 56704 10166 56706 10218
rect 56650 10164 56706 10166
rect 56442 8650 56498 8652
rect 56442 8598 56444 8650
rect 56444 8598 56496 8650
rect 56496 8598 56498 8650
rect 56442 8596 56498 8598
rect 56546 8650 56602 8652
rect 56546 8598 56548 8650
rect 56548 8598 56600 8650
rect 56600 8598 56602 8650
rect 56546 8596 56602 8598
rect 56650 8650 56706 8652
rect 56650 8598 56652 8650
rect 56652 8598 56704 8650
rect 56704 8598 56706 8650
rect 56650 8596 56706 8598
rect 56442 7082 56498 7084
rect 56442 7030 56444 7082
rect 56444 7030 56496 7082
rect 56496 7030 56498 7082
rect 56442 7028 56498 7030
rect 56546 7082 56602 7084
rect 56546 7030 56548 7082
rect 56548 7030 56600 7082
rect 56600 7030 56602 7082
rect 56546 7028 56602 7030
rect 56650 7082 56706 7084
rect 56650 7030 56652 7082
rect 56652 7030 56704 7082
rect 56704 7030 56706 7082
rect 56650 7028 56706 7030
rect 54460 5234 54516 5236
rect 54460 5182 54462 5234
rect 54462 5182 54514 5234
rect 54514 5182 54516 5234
rect 54460 5180 54516 5182
rect 55692 4956 55748 5012
rect 55020 4562 55076 4564
rect 55020 4510 55022 4562
rect 55022 4510 55074 4562
rect 55074 4510 55076 4562
rect 55020 4508 55076 4510
rect 56442 5514 56498 5516
rect 56442 5462 56444 5514
rect 56444 5462 56496 5514
rect 56496 5462 56498 5514
rect 56442 5460 56498 5462
rect 56546 5514 56602 5516
rect 56546 5462 56548 5514
rect 56548 5462 56600 5514
rect 56600 5462 56602 5514
rect 56546 5460 56602 5462
rect 56650 5514 56706 5516
rect 56650 5462 56652 5514
rect 56652 5462 56704 5514
rect 56704 5462 56706 5514
rect 56650 5460 56706 5462
rect 56812 4898 56868 4900
rect 56812 4846 56814 4898
rect 56814 4846 56866 4898
rect 56866 4846 56868 4898
rect 56812 4844 56868 4846
rect 57260 4898 57316 4900
rect 57260 4846 57262 4898
rect 57262 4846 57314 4898
rect 57314 4846 57316 4898
rect 57260 4844 57316 4846
rect 56476 4508 56532 4564
rect 56812 4396 56868 4452
rect 56442 3946 56498 3948
rect 56442 3894 56444 3946
rect 56444 3894 56496 3946
rect 56496 3894 56498 3946
rect 56442 3892 56498 3894
rect 56546 3946 56602 3948
rect 56546 3894 56548 3946
rect 56548 3894 56600 3946
rect 56600 3894 56602 3946
rect 56546 3892 56602 3894
rect 56650 3946 56706 3948
rect 56650 3894 56652 3946
rect 56652 3894 56704 3946
rect 56704 3894 56706 3946
rect 56650 3892 56706 3894
rect 55916 3276 55972 3332
rect 56700 3276 56756 3332
rect 57820 5068 57876 5124
rect 57596 4450 57652 4452
rect 57596 4398 57598 4450
rect 57598 4398 57650 4450
rect 57650 4398 57652 4450
rect 57596 4396 57652 4398
rect 57036 3948 57092 4004
rect 58156 4844 58212 4900
rect 60396 31052 60452 31108
rect 60732 30940 60788 30996
rect 62524 37660 62580 37716
rect 61516 32620 61572 32676
rect 60844 30828 60900 30884
rect 60396 30268 60452 30324
rect 62300 35196 62356 35252
rect 62412 35420 62468 35476
rect 61964 33852 62020 33908
rect 62412 34412 62468 34468
rect 62636 35586 62692 35588
rect 62636 35534 62638 35586
rect 62638 35534 62690 35586
rect 62690 35534 62692 35586
rect 62636 35532 62692 35534
rect 63644 37772 63700 37828
rect 64092 37436 64148 37492
rect 63084 35532 63140 35588
rect 61852 32172 61908 32228
rect 61740 30268 61796 30324
rect 62300 32786 62356 32788
rect 62300 32734 62302 32786
rect 62302 32734 62354 32786
rect 62354 32734 62356 32786
rect 62300 32732 62356 32734
rect 63420 33122 63476 33124
rect 63420 33070 63422 33122
rect 63422 33070 63474 33122
rect 63474 33070 63476 33122
rect 63420 33068 63476 33070
rect 63196 32786 63252 32788
rect 63196 32734 63198 32786
rect 63198 32734 63250 32786
rect 63250 32734 63252 32786
rect 63196 32732 63252 32734
rect 65436 37436 65492 37492
rect 63644 33852 63700 33908
rect 63980 33852 64036 33908
rect 63868 33122 63924 33124
rect 63868 33070 63870 33122
rect 63870 33070 63922 33122
rect 63922 33070 63924 33122
rect 63868 33068 63924 33070
rect 63308 31836 63364 31892
rect 62972 31724 63028 31780
rect 62188 24332 62244 24388
rect 62636 25116 62692 25172
rect 61628 24108 61684 24164
rect 60396 23212 60452 23268
rect 61740 22988 61796 23044
rect 59836 10892 59892 10948
rect 60844 6412 60900 6468
rect 59948 6300 60004 6356
rect 60396 6300 60452 6356
rect 58828 3948 58884 4004
rect 58044 3612 58100 3668
rect 60844 6130 60900 6132
rect 60844 6078 60846 6130
rect 60846 6078 60898 6130
rect 60898 6078 60900 6130
rect 60844 6076 60900 6078
rect 59836 3948 59892 4004
rect 59388 3500 59444 3556
rect 59612 3666 59668 3668
rect 59612 3614 59614 3666
rect 59614 3614 59666 3666
rect 59666 3614 59668 3666
rect 59612 3612 59668 3614
rect 60620 5180 60676 5236
rect 61740 5068 61796 5124
rect 60844 3554 60900 3556
rect 60844 3502 60846 3554
rect 60846 3502 60898 3554
rect 60898 3502 60900 3554
rect 60844 3500 60900 3502
rect 61964 3836 62020 3892
rect 62300 5180 62356 5236
rect 64428 33516 64484 33572
rect 64876 35420 64932 35476
rect 64764 33516 64820 33572
rect 65100 33852 65156 33908
rect 64540 32732 64596 32788
rect 64428 31948 64484 32004
rect 64876 31890 64932 31892
rect 64876 31838 64878 31890
rect 64878 31838 64930 31890
rect 64930 31838 64932 31890
rect 64876 31836 64932 31838
rect 65548 36316 65604 36372
rect 65660 37884 65716 37940
rect 65884 36370 65940 36372
rect 65884 36318 65886 36370
rect 65886 36318 65938 36370
rect 65938 36318 65940 36370
rect 65884 36316 65940 36318
rect 65548 35420 65604 35476
rect 66332 35474 66388 35476
rect 66332 35422 66334 35474
rect 66334 35422 66386 35474
rect 66386 35422 66388 35474
rect 66332 35420 66388 35422
rect 65660 34018 65716 34020
rect 65660 33966 65662 34018
rect 65662 33966 65714 34018
rect 65714 33966 65716 34018
rect 65660 33964 65716 33966
rect 66220 35308 66276 35364
rect 65884 33068 65940 33124
rect 65996 33292 66052 33348
rect 64988 29484 65044 29540
rect 64316 27692 64372 27748
rect 67228 38332 67284 38388
rect 66556 36876 66612 36932
rect 68012 37548 68068 37604
rect 66556 34300 66612 34356
rect 67004 35420 67060 35476
rect 66780 34690 66836 34692
rect 66780 34638 66782 34690
rect 66782 34638 66834 34690
rect 66834 34638 66836 34690
rect 66780 34636 66836 34638
rect 66668 33292 66724 33348
rect 66668 33122 66724 33124
rect 66668 33070 66670 33122
rect 66670 33070 66722 33122
rect 66722 33070 66724 33122
rect 66668 33068 66724 33070
rect 67116 34748 67172 34804
rect 67340 34802 67396 34804
rect 67340 34750 67342 34802
rect 67342 34750 67394 34802
rect 67394 34750 67396 34802
rect 67340 34748 67396 34750
rect 67900 34636 67956 34692
rect 68124 35138 68180 35140
rect 68124 35086 68126 35138
rect 68126 35086 68178 35138
rect 68178 35086 68180 35138
rect 68124 35084 68180 35086
rect 69020 37548 69076 37604
rect 68460 36594 68516 36596
rect 68460 36542 68462 36594
rect 68462 36542 68514 36594
rect 68514 36542 68516 36594
rect 68460 36540 68516 36542
rect 68908 36370 68964 36372
rect 68908 36318 68910 36370
rect 68910 36318 68962 36370
rect 68962 36318 68964 36370
rect 68908 36316 68964 36318
rect 68908 35532 68964 35588
rect 69916 38444 69972 38500
rect 69132 36540 69188 36596
rect 69804 37884 69860 37940
rect 69692 36204 69748 36260
rect 69692 35922 69748 35924
rect 69692 35870 69694 35922
rect 69694 35870 69746 35922
rect 69746 35870 69748 35922
rect 69692 35868 69748 35870
rect 69356 35084 69412 35140
rect 68236 34300 68292 34356
rect 67340 34130 67396 34132
rect 67340 34078 67342 34130
rect 67342 34078 67394 34130
rect 67394 34078 67396 34130
rect 67340 34076 67396 34078
rect 68236 34076 68292 34132
rect 67340 32956 67396 33012
rect 67228 32732 67284 32788
rect 66668 31948 66724 32004
rect 62860 8764 62916 8820
rect 62524 5068 62580 5124
rect 62188 4956 62244 5012
rect 63868 7474 63924 7476
rect 63868 7422 63870 7474
rect 63870 7422 63922 7474
rect 63922 7422 63924 7474
rect 63868 7420 63924 7422
rect 63196 4956 63252 5012
rect 62188 3388 62244 3444
rect 64652 9154 64708 9156
rect 64652 9102 64654 9154
rect 64654 9102 64706 9154
rect 64706 9102 64708 9154
rect 64652 9100 64708 9102
rect 64876 9100 64932 9156
rect 64092 6524 64148 6580
rect 64652 6636 64708 6692
rect 65548 8818 65604 8820
rect 65548 8766 65550 8818
rect 65550 8766 65602 8818
rect 65602 8766 65604 8818
rect 65548 8764 65604 8766
rect 65996 9212 66052 9268
rect 67228 9266 67284 9268
rect 67228 9214 67230 9266
rect 67230 9214 67282 9266
rect 67282 9214 67284 9266
rect 67228 9212 67284 9214
rect 65772 8316 65828 8372
rect 65548 7474 65604 7476
rect 65548 7422 65550 7474
rect 65550 7422 65602 7474
rect 65602 7422 65604 7474
rect 65548 7420 65604 7422
rect 66444 9154 66500 9156
rect 66444 9102 66446 9154
rect 66446 9102 66498 9154
rect 66498 9102 66500 9154
rect 66444 9100 66500 9102
rect 68572 34636 68628 34692
rect 69468 34690 69524 34692
rect 69468 34638 69470 34690
rect 69470 34638 69522 34690
rect 69522 34638 69524 34690
rect 69468 34636 69524 34638
rect 69468 33964 69524 34020
rect 71148 38556 71204 38612
rect 70812 38220 70868 38276
rect 69916 35084 69972 35140
rect 69916 34300 69972 34356
rect 70252 33404 70308 33460
rect 71148 34076 71204 34132
rect 73164 37212 73220 37268
rect 71708 36594 71764 36596
rect 71708 36542 71710 36594
rect 71710 36542 71762 36594
rect 71762 36542 71764 36594
rect 71708 36540 71764 36542
rect 72380 36370 72436 36372
rect 72380 36318 72382 36370
rect 72382 36318 72434 36370
rect 72434 36318 72436 36370
rect 72380 36316 72436 36318
rect 72492 36258 72548 36260
rect 72492 36206 72494 36258
rect 72494 36206 72546 36258
rect 72546 36206 72548 36258
rect 72492 36204 72548 36206
rect 73500 37324 73556 37380
rect 72716 35644 72772 35700
rect 70812 31948 70868 32004
rect 69468 30044 69524 30100
rect 71932 31836 71988 31892
rect 73612 34972 73668 35028
rect 73724 37324 73780 37380
rect 73276 34748 73332 34804
rect 74508 36540 74564 36596
rect 75292 38668 75348 38724
rect 74852 36090 74908 36092
rect 74852 36038 74854 36090
rect 74854 36038 74906 36090
rect 74906 36038 74908 36090
rect 74852 36036 74908 36038
rect 74956 36090 75012 36092
rect 74956 36038 74958 36090
rect 74958 36038 75010 36090
rect 75010 36038 75012 36090
rect 74956 36036 75012 36038
rect 75060 36090 75116 36092
rect 75060 36038 75062 36090
rect 75062 36038 75114 36090
rect 75114 36038 75116 36090
rect 75060 36036 75116 36038
rect 74732 35756 74788 35812
rect 74508 35026 74564 35028
rect 74508 34974 74510 35026
rect 74510 34974 74562 35026
rect 74562 34974 74564 35026
rect 74508 34972 74564 34974
rect 73500 34130 73556 34132
rect 73500 34078 73502 34130
rect 73502 34078 73554 34130
rect 73554 34078 73556 34130
rect 73500 34076 73556 34078
rect 74172 34860 74228 34916
rect 75292 35756 75348 35812
rect 74844 35586 74900 35588
rect 74844 35534 74846 35586
rect 74846 35534 74898 35586
rect 74898 35534 74900 35586
rect 74844 35532 74900 35534
rect 74852 34522 74908 34524
rect 74852 34470 74854 34522
rect 74854 34470 74906 34522
rect 74906 34470 74908 34522
rect 74852 34468 74908 34470
rect 74956 34522 75012 34524
rect 74956 34470 74958 34522
rect 74958 34470 75010 34522
rect 75010 34470 75012 34522
rect 74956 34468 75012 34470
rect 75060 34522 75116 34524
rect 75060 34470 75062 34522
rect 75062 34470 75114 34522
rect 75114 34470 75116 34522
rect 75060 34468 75116 34470
rect 75628 36988 75684 37044
rect 75628 35810 75684 35812
rect 75628 35758 75630 35810
rect 75630 35758 75682 35810
rect 75682 35758 75684 35810
rect 75628 35756 75684 35758
rect 75740 34412 75796 34468
rect 74172 34076 74228 34132
rect 75068 33852 75124 33908
rect 75740 33852 75796 33908
rect 76300 35756 76356 35812
rect 76412 37996 76468 38052
rect 77196 36764 77252 36820
rect 77308 37996 77364 38052
rect 78764 38668 78820 38724
rect 78652 37996 78708 38052
rect 76300 35474 76356 35476
rect 76300 35422 76302 35474
rect 76302 35422 76354 35474
rect 76354 35422 76356 35474
rect 76300 35420 76356 35422
rect 76076 34636 76132 34692
rect 72380 28476 72436 28532
rect 71484 28364 71540 28420
rect 71708 22876 71764 22932
rect 67676 8370 67732 8372
rect 67676 8318 67678 8370
rect 67678 8318 67730 8370
rect 67730 8318 67732 8370
rect 67676 8316 67732 8318
rect 65884 7196 65940 7252
rect 65324 6466 65380 6468
rect 65324 6414 65326 6466
rect 65326 6414 65378 6466
rect 65378 6414 65380 6466
rect 65324 6412 65380 6414
rect 65548 6130 65604 6132
rect 65548 6078 65550 6130
rect 65550 6078 65602 6130
rect 65602 6078 65604 6130
rect 65548 6076 65604 6078
rect 64876 5740 64932 5796
rect 66444 7196 66500 7252
rect 66332 6578 66388 6580
rect 66332 6526 66334 6578
rect 66334 6526 66386 6578
rect 66386 6526 66388 6578
rect 66332 6524 66388 6526
rect 66668 5964 66724 6020
rect 66108 5906 66164 5908
rect 66108 5854 66110 5906
rect 66110 5854 66162 5906
rect 66162 5854 66164 5906
rect 66108 5852 66164 5854
rect 66668 5628 66724 5684
rect 67228 7196 67284 7252
rect 67340 6748 67396 6804
rect 67564 6578 67620 6580
rect 67564 6526 67566 6578
rect 67566 6526 67618 6578
rect 67618 6526 67620 6578
rect 67564 6524 67620 6526
rect 67564 6300 67620 6356
rect 67340 5964 67396 6020
rect 66780 5516 66836 5572
rect 67116 5740 67172 5796
rect 68124 6914 68180 6916
rect 68124 6862 68126 6914
rect 68126 6862 68178 6914
rect 68178 6862 68180 6914
rect 68124 6860 68180 6862
rect 68236 6636 68292 6692
rect 67788 5628 67844 5684
rect 67900 5852 67956 5908
rect 67004 5180 67060 5236
rect 65884 4508 65940 4564
rect 66668 4284 66724 4340
rect 67564 5068 67620 5124
rect 64652 3666 64708 3668
rect 64652 3614 64654 3666
rect 64654 3614 64706 3666
rect 64706 3614 64708 3666
rect 64652 3612 64708 3614
rect 64876 3500 64932 3556
rect 65212 3500 65268 3556
rect 68460 5516 68516 5572
rect 67676 3836 67732 3892
rect 68684 6076 68740 6132
rect 71708 12684 71764 12740
rect 76188 34524 76244 34580
rect 76300 34354 76356 34356
rect 76300 34302 76302 34354
rect 76302 34302 76354 34354
rect 76354 34302 76356 34354
rect 76300 34300 76356 34302
rect 74852 32954 74908 32956
rect 74852 32902 74854 32954
rect 74854 32902 74906 32954
rect 74906 32902 74908 32954
rect 74852 32900 74908 32902
rect 74956 32954 75012 32956
rect 74956 32902 74958 32954
rect 74958 32902 75010 32954
rect 75010 32902 75012 32954
rect 74956 32900 75012 32902
rect 75060 32954 75116 32956
rect 75060 32902 75062 32954
rect 75062 32902 75114 32954
rect 75114 32902 75116 32954
rect 75060 32900 75116 32902
rect 74852 31386 74908 31388
rect 74852 31334 74854 31386
rect 74854 31334 74906 31386
rect 74906 31334 74908 31386
rect 74852 31332 74908 31334
rect 74956 31386 75012 31388
rect 74956 31334 74958 31386
rect 74958 31334 75010 31386
rect 75010 31334 75012 31386
rect 74956 31332 75012 31334
rect 75060 31386 75116 31388
rect 75060 31334 75062 31386
rect 75062 31334 75114 31386
rect 75114 31334 75116 31386
rect 75060 31332 75116 31334
rect 74852 29818 74908 29820
rect 74852 29766 74854 29818
rect 74854 29766 74906 29818
rect 74906 29766 74908 29818
rect 74852 29764 74908 29766
rect 74956 29818 75012 29820
rect 74956 29766 74958 29818
rect 74958 29766 75010 29818
rect 75010 29766 75012 29818
rect 74956 29764 75012 29766
rect 75060 29818 75116 29820
rect 75060 29766 75062 29818
rect 75062 29766 75114 29818
rect 75114 29766 75116 29818
rect 75060 29764 75116 29766
rect 74852 28250 74908 28252
rect 74852 28198 74854 28250
rect 74854 28198 74906 28250
rect 74906 28198 74908 28250
rect 74852 28196 74908 28198
rect 74956 28250 75012 28252
rect 74956 28198 74958 28250
rect 74958 28198 75010 28250
rect 75010 28198 75012 28250
rect 74956 28196 75012 28198
rect 75060 28250 75116 28252
rect 75060 28198 75062 28250
rect 75062 28198 75114 28250
rect 75114 28198 75116 28250
rect 75060 28196 75116 28198
rect 75516 26908 75572 26964
rect 74852 26682 74908 26684
rect 74852 26630 74854 26682
rect 74854 26630 74906 26682
rect 74906 26630 74908 26682
rect 74852 26628 74908 26630
rect 74956 26682 75012 26684
rect 74956 26630 74958 26682
rect 74958 26630 75010 26682
rect 75010 26630 75012 26682
rect 74956 26628 75012 26630
rect 75060 26682 75116 26684
rect 75060 26630 75062 26682
rect 75062 26630 75114 26682
rect 75114 26630 75116 26682
rect 75060 26628 75116 26630
rect 74852 25114 74908 25116
rect 74852 25062 74854 25114
rect 74854 25062 74906 25114
rect 74906 25062 74908 25114
rect 74852 25060 74908 25062
rect 74956 25114 75012 25116
rect 74956 25062 74958 25114
rect 74958 25062 75010 25114
rect 75010 25062 75012 25114
rect 74956 25060 75012 25062
rect 75060 25114 75116 25116
rect 75060 25062 75062 25114
rect 75062 25062 75114 25114
rect 75114 25062 75116 25114
rect 75060 25060 75116 25062
rect 74852 23546 74908 23548
rect 74852 23494 74854 23546
rect 74854 23494 74906 23546
rect 74906 23494 74908 23546
rect 74852 23492 74908 23494
rect 74956 23546 75012 23548
rect 74956 23494 74958 23546
rect 74958 23494 75010 23546
rect 75010 23494 75012 23546
rect 74956 23492 75012 23494
rect 75060 23546 75116 23548
rect 75060 23494 75062 23546
rect 75062 23494 75114 23546
rect 75114 23494 75116 23546
rect 75060 23492 75116 23494
rect 74852 21978 74908 21980
rect 74852 21926 74854 21978
rect 74854 21926 74906 21978
rect 74906 21926 74908 21978
rect 74852 21924 74908 21926
rect 74956 21978 75012 21980
rect 74956 21926 74958 21978
rect 74958 21926 75010 21978
rect 75010 21926 75012 21978
rect 74956 21924 75012 21926
rect 75060 21978 75116 21980
rect 75060 21926 75062 21978
rect 75062 21926 75114 21978
rect 75114 21926 75116 21978
rect 75060 21924 75116 21926
rect 74852 20410 74908 20412
rect 74852 20358 74854 20410
rect 74854 20358 74906 20410
rect 74906 20358 74908 20410
rect 74852 20356 74908 20358
rect 74956 20410 75012 20412
rect 74956 20358 74958 20410
rect 74958 20358 75010 20410
rect 75010 20358 75012 20410
rect 74956 20356 75012 20358
rect 75060 20410 75116 20412
rect 75060 20358 75062 20410
rect 75062 20358 75114 20410
rect 75114 20358 75116 20410
rect 75060 20356 75116 20358
rect 74852 18842 74908 18844
rect 74852 18790 74854 18842
rect 74854 18790 74906 18842
rect 74906 18790 74908 18842
rect 74852 18788 74908 18790
rect 74956 18842 75012 18844
rect 74956 18790 74958 18842
rect 74958 18790 75010 18842
rect 75010 18790 75012 18842
rect 74956 18788 75012 18790
rect 75060 18842 75116 18844
rect 75060 18790 75062 18842
rect 75062 18790 75114 18842
rect 75114 18790 75116 18842
rect 75060 18788 75116 18790
rect 74852 17274 74908 17276
rect 74852 17222 74854 17274
rect 74854 17222 74906 17274
rect 74906 17222 74908 17274
rect 74852 17220 74908 17222
rect 74956 17274 75012 17276
rect 74956 17222 74958 17274
rect 74958 17222 75010 17274
rect 75010 17222 75012 17274
rect 74956 17220 75012 17222
rect 75060 17274 75116 17276
rect 75060 17222 75062 17274
rect 75062 17222 75114 17274
rect 75114 17222 75116 17274
rect 75060 17220 75116 17222
rect 74852 15706 74908 15708
rect 74852 15654 74854 15706
rect 74854 15654 74906 15706
rect 74906 15654 74908 15706
rect 74852 15652 74908 15654
rect 74956 15706 75012 15708
rect 74956 15654 74958 15706
rect 74958 15654 75010 15706
rect 75010 15654 75012 15706
rect 74956 15652 75012 15654
rect 75060 15706 75116 15708
rect 75060 15654 75062 15706
rect 75062 15654 75114 15706
rect 75114 15654 75116 15706
rect 75060 15652 75116 15654
rect 74852 14138 74908 14140
rect 74852 14086 74854 14138
rect 74854 14086 74906 14138
rect 74906 14086 74908 14138
rect 74852 14084 74908 14086
rect 74956 14138 75012 14140
rect 74956 14086 74958 14138
rect 74958 14086 75010 14138
rect 75010 14086 75012 14138
rect 74956 14084 75012 14086
rect 75060 14138 75116 14140
rect 75060 14086 75062 14138
rect 75062 14086 75114 14138
rect 75114 14086 75116 14138
rect 75060 14084 75116 14086
rect 74852 12570 74908 12572
rect 74852 12518 74854 12570
rect 74854 12518 74906 12570
rect 74906 12518 74908 12570
rect 74852 12516 74908 12518
rect 74956 12570 75012 12572
rect 74956 12518 74958 12570
rect 74958 12518 75010 12570
rect 75010 12518 75012 12570
rect 74956 12516 75012 12518
rect 75060 12570 75116 12572
rect 75060 12518 75062 12570
rect 75062 12518 75114 12570
rect 75114 12518 75116 12570
rect 75060 12516 75116 12518
rect 73724 11676 73780 11732
rect 74852 11002 74908 11004
rect 74852 10950 74854 11002
rect 74854 10950 74906 11002
rect 74906 10950 74908 11002
rect 74852 10948 74908 10950
rect 74956 11002 75012 11004
rect 74956 10950 74958 11002
rect 74958 10950 75010 11002
rect 75010 10950 75012 11002
rect 74956 10948 75012 10950
rect 75060 11002 75116 11004
rect 75060 10950 75062 11002
rect 75062 10950 75114 11002
rect 75114 10950 75116 11002
rect 75060 10948 75116 10950
rect 74852 9434 74908 9436
rect 74852 9382 74854 9434
rect 74854 9382 74906 9434
rect 74906 9382 74908 9434
rect 74852 9380 74908 9382
rect 74956 9434 75012 9436
rect 74956 9382 74958 9434
rect 74958 9382 75010 9434
rect 75010 9382 75012 9434
rect 74956 9380 75012 9382
rect 75060 9434 75116 9436
rect 75060 9382 75062 9434
rect 75062 9382 75114 9434
rect 75114 9382 75116 9434
rect 75060 9380 75116 9382
rect 69468 6860 69524 6916
rect 69132 6524 69188 6580
rect 69356 6466 69412 6468
rect 69356 6414 69358 6466
rect 69358 6414 69410 6466
rect 69410 6414 69412 6466
rect 69356 6412 69412 6414
rect 69132 5852 69188 5908
rect 68684 5740 68740 5796
rect 69468 5122 69524 5124
rect 69468 5070 69470 5122
rect 69470 5070 69522 5122
rect 69522 5070 69524 5122
rect 69468 5068 69524 5070
rect 69356 4844 69412 4900
rect 68572 4284 68628 4340
rect 69244 4338 69300 4340
rect 69244 4286 69246 4338
rect 69246 4286 69298 4338
rect 69298 4286 69300 4338
rect 69244 4284 69300 4286
rect 68572 3666 68628 3668
rect 68572 3614 68574 3666
rect 68574 3614 68626 3666
rect 68626 3614 68628 3666
rect 68572 3612 68628 3614
rect 69356 3612 69412 3668
rect 70140 5964 70196 6020
rect 70476 5628 70532 5684
rect 71148 6018 71204 6020
rect 71148 5966 71150 6018
rect 71150 5966 71202 6018
rect 71202 5966 71204 6018
rect 71148 5964 71204 5966
rect 70700 5906 70756 5908
rect 70700 5854 70702 5906
rect 70702 5854 70754 5906
rect 70754 5854 70756 5906
rect 70700 5852 70756 5854
rect 71484 5010 71540 5012
rect 71484 4958 71486 5010
rect 71486 4958 71538 5010
rect 71538 4958 71540 5010
rect 71484 4956 71540 4958
rect 71148 4898 71204 4900
rect 71148 4846 71150 4898
rect 71150 4846 71202 4898
rect 71202 4846 71204 4898
rect 71148 4844 71204 4846
rect 70588 2492 70644 2548
rect 74852 7866 74908 7868
rect 74852 7814 74854 7866
rect 74854 7814 74906 7866
rect 74906 7814 74908 7866
rect 74852 7812 74908 7814
rect 74956 7866 75012 7868
rect 74956 7814 74958 7866
rect 74958 7814 75010 7866
rect 75010 7814 75012 7866
rect 74956 7812 75012 7814
rect 75060 7866 75116 7868
rect 75060 7814 75062 7866
rect 75062 7814 75114 7866
rect 75114 7814 75116 7866
rect 75060 7812 75116 7814
rect 74620 7308 74676 7364
rect 74060 7196 74116 7252
rect 72604 6524 72660 6580
rect 72156 6130 72212 6132
rect 72156 6078 72158 6130
rect 72158 6078 72210 6130
rect 72210 6078 72212 6130
rect 72156 6076 72212 6078
rect 73276 6578 73332 6580
rect 73276 6526 73278 6578
rect 73278 6526 73330 6578
rect 73330 6526 73332 6578
rect 73276 6524 73332 6526
rect 72380 5292 72436 5348
rect 71932 5010 71988 5012
rect 71932 4958 71934 5010
rect 71934 4958 71986 5010
rect 71986 4958 71988 5010
rect 71932 4956 71988 4958
rect 72940 5964 72996 6020
rect 72940 5346 72996 5348
rect 72940 5294 72942 5346
rect 72942 5294 72994 5346
rect 72994 5294 72996 5346
rect 72940 5292 72996 5294
rect 72492 5068 72548 5124
rect 72492 4284 72548 4340
rect 72604 3554 72660 3556
rect 72604 3502 72606 3554
rect 72606 3502 72658 3554
rect 72658 3502 72660 3554
rect 72604 3500 72660 3502
rect 73724 4898 73780 4900
rect 73724 4846 73726 4898
rect 73726 4846 73778 4898
rect 73778 4846 73780 4898
rect 73724 4844 73780 4846
rect 77308 35698 77364 35700
rect 77308 35646 77310 35698
rect 77310 35646 77362 35698
rect 77362 35646 77364 35698
rect 77308 35644 77364 35646
rect 76860 34524 76916 34580
rect 76860 34300 76916 34356
rect 77756 33404 77812 33460
rect 78092 35756 78148 35812
rect 78204 34802 78260 34804
rect 78204 34750 78206 34802
rect 78206 34750 78258 34802
rect 78258 34750 78260 34802
rect 78204 34748 78260 34750
rect 77644 33068 77700 33124
rect 77196 31276 77252 31332
rect 76636 26908 76692 26964
rect 77980 24668 78036 24724
rect 75068 7362 75124 7364
rect 75068 7310 75070 7362
rect 75070 7310 75122 7362
rect 75122 7310 75124 7362
rect 75068 7308 75124 7310
rect 75180 7196 75236 7252
rect 74852 6298 74908 6300
rect 74852 6246 74854 6298
rect 74854 6246 74906 6298
rect 74906 6246 74908 6298
rect 74852 6244 74908 6246
rect 74956 6298 75012 6300
rect 74956 6246 74958 6298
rect 74958 6246 75010 6298
rect 75010 6246 75012 6298
rect 74956 6244 75012 6246
rect 75060 6298 75116 6300
rect 75060 6246 75062 6298
rect 75062 6246 75114 6298
rect 75114 6246 75116 6298
rect 75060 6244 75116 6246
rect 74732 6018 74788 6020
rect 74732 5966 74734 6018
rect 74734 5966 74786 6018
rect 74786 5966 74788 6018
rect 74732 5964 74788 5966
rect 75852 12796 75908 12852
rect 75740 6524 75796 6580
rect 75628 5068 75684 5124
rect 74852 4730 74908 4732
rect 74852 4678 74854 4730
rect 74854 4678 74906 4730
rect 74906 4678 74908 4730
rect 74852 4676 74908 4678
rect 74956 4730 75012 4732
rect 74956 4678 74958 4730
rect 74958 4678 75010 4730
rect 75010 4678 75012 4730
rect 74956 4676 75012 4678
rect 75060 4730 75116 4732
rect 75060 4678 75062 4730
rect 75062 4678 75114 4730
rect 75114 4678 75116 4730
rect 75060 4676 75116 4678
rect 76972 12796 77028 12852
rect 76972 11788 77028 11844
rect 78428 35532 78484 35588
rect 78540 34802 78596 34804
rect 78540 34750 78542 34802
rect 78542 34750 78594 34802
rect 78594 34750 78596 34802
rect 78540 34748 78596 34750
rect 78988 36764 79044 36820
rect 79100 36316 79156 36372
rect 78764 35420 78820 35476
rect 78988 34524 79044 34580
rect 79436 34802 79492 34804
rect 79436 34750 79438 34802
rect 79438 34750 79490 34802
rect 79490 34750 79492 34802
rect 79436 34748 79492 34750
rect 79100 29596 79156 29652
rect 79772 35586 79828 35588
rect 79772 35534 79774 35586
rect 79774 35534 79826 35586
rect 79826 35534 79828 35586
rect 79772 35532 79828 35534
rect 81564 37212 81620 37268
rect 81228 36370 81284 36372
rect 81228 36318 81230 36370
rect 81230 36318 81282 36370
rect 81282 36318 81284 36370
rect 81228 36316 81284 36318
rect 82796 38892 82852 38948
rect 82572 37100 82628 37156
rect 82236 36204 82292 36260
rect 80892 35084 80948 35140
rect 80444 34748 80500 34804
rect 80444 33852 80500 33908
rect 80556 33180 80612 33236
rect 81788 34300 81844 34356
rect 81340 33180 81396 33236
rect 83020 36370 83076 36372
rect 83020 36318 83022 36370
rect 83022 36318 83074 36370
rect 83074 36318 83076 36370
rect 83020 36316 83076 36318
rect 84028 38108 84084 38164
rect 83468 35756 83524 35812
rect 82572 35084 82628 35140
rect 82572 34748 82628 34804
rect 83804 34748 83860 34804
rect 82684 34300 82740 34356
rect 83804 34130 83860 34132
rect 83804 34078 83806 34130
rect 83806 34078 83858 34130
rect 83858 34078 83860 34130
rect 83804 34076 83860 34078
rect 84924 36258 84980 36260
rect 84924 36206 84926 36258
rect 84926 36206 84978 36258
rect 84978 36206 84980 36258
rect 84924 36204 84980 36206
rect 84476 36092 84532 36148
rect 84924 35810 84980 35812
rect 84924 35758 84926 35810
rect 84926 35758 84978 35810
rect 84978 35758 84980 35810
rect 84924 35756 84980 35758
rect 85820 38780 85876 38836
rect 86156 36428 86212 36484
rect 86828 36428 86884 36484
rect 85260 35756 85316 35812
rect 86716 35810 86772 35812
rect 86716 35758 86718 35810
rect 86718 35758 86770 35810
rect 86770 35758 86772 35810
rect 86716 35756 86772 35758
rect 84364 35084 84420 35140
rect 84140 34076 84196 34132
rect 84588 32956 84644 33012
rect 85932 35084 85988 35140
rect 87052 35084 87108 35140
rect 82236 32620 82292 32676
rect 82012 31164 82068 31220
rect 81452 29932 81508 29988
rect 85148 27916 85204 27972
rect 79772 27804 79828 27860
rect 79660 27580 79716 27636
rect 87948 35084 88004 35140
rect 87612 34354 87668 34356
rect 87612 34302 87614 34354
rect 87614 34302 87666 34354
rect 87666 34302 87668 34354
rect 87612 34300 87668 34302
rect 87612 33628 87668 33684
rect 88620 34748 88676 34804
rect 88396 34300 88452 34356
rect 88508 34636 88564 34692
rect 88172 34018 88228 34020
rect 88172 33966 88174 34018
rect 88174 33966 88226 34018
rect 88226 33966 88228 34018
rect 88172 33964 88228 33966
rect 88060 33404 88116 33460
rect 87724 30828 87780 30884
rect 87500 27244 87556 27300
rect 87052 26460 87108 26516
rect 85484 26124 85540 26180
rect 80668 24332 80724 24388
rect 79772 22988 79828 23044
rect 86492 22876 86548 22932
rect 84924 21308 84980 21364
rect 83132 20972 83188 21028
rect 79772 11788 79828 11844
rect 76076 6412 76132 6468
rect 76972 7474 77028 7476
rect 76972 7422 76974 7474
rect 76974 7422 77026 7474
rect 77026 7422 77028 7474
rect 76972 7420 77028 7422
rect 78316 7420 78372 7476
rect 78428 11676 78484 11732
rect 76748 7196 76804 7252
rect 77868 7196 77924 7252
rect 77644 6578 77700 6580
rect 77644 6526 77646 6578
rect 77646 6526 77698 6578
rect 77698 6526 77700 6578
rect 77644 6524 77700 6526
rect 77308 6466 77364 6468
rect 77308 6414 77310 6466
rect 77310 6414 77362 6466
rect 77362 6414 77364 6466
rect 77308 6412 77364 6414
rect 76300 5682 76356 5684
rect 76300 5630 76302 5682
rect 76302 5630 76354 5682
rect 76354 5630 76356 5682
rect 76300 5628 76356 5630
rect 76300 5068 76356 5124
rect 76636 5122 76692 5124
rect 76636 5070 76638 5122
rect 76638 5070 76690 5122
rect 76690 5070 76692 5122
rect 76636 5068 76692 5070
rect 77308 5180 77364 5236
rect 77084 3724 77140 3780
rect 80780 8316 80836 8372
rect 78540 6466 78596 6468
rect 78540 6414 78542 6466
rect 78542 6414 78594 6466
rect 78594 6414 78596 6466
rect 78540 6412 78596 6414
rect 79324 6412 79380 6468
rect 79212 3778 79268 3780
rect 79212 3726 79214 3778
rect 79214 3726 79266 3778
rect 79266 3726 79268 3778
rect 79212 3724 79268 3726
rect 79324 3666 79380 3668
rect 79324 3614 79326 3666
rect 79326 3614 79378 3666
rect 79378 3614 79380 3666
rect 79324 3612 79380 3614
rect 76972 3500 77028 3556
rect 73836 3388 73892 3444
rect 75628 3388 75684 3444
rect 74852 3162 74908 3164
rect 74852 3110 74854 3162
rect 74854 3110 74906 3162
rect 74906 3110 74908 3162
rect 74852 3108 74908 3110
rect 74956 3162 75012 3164
rect 74956 3110 74958 3162
rect 74958 3110 75010 3162
rect 75010 3110 75012 3162
rect 74956 3108 75012 3110
rect 75060 3162 75116 3164
rect 75060 3110 75062 3162
rect 75062 3110 75114 3162
rect 75114 3110 75116 3162
rect 75060 3108 75116 3110
rect 77308 3500 77364 3556
rect 80444 5068 80500 5124
rect 80220 4844 80276 4900
rect 80444 4620 80500 4676
rect 84924 15932 84980 15988
rect 83132 8316 83188 8372
rect 84700 14252 84756 14308
rect 81788 7532 81844 7588
rect 81116 6524 81172 6580
rect 81564 6578 81620 6580
rect 81564 6526 81566 6578
rect 81566 6526 81618 6578
rect 81618 6526 81620 6578
rect 81564 6524 81620 6526
rect 81228 4620 81284 4676
rect 81676 4620 81732 4676
rect 84476 5122 84532 5124
rect 84476 5070 84478 5122
rect 84478 5070 84530 5122
rect 84530 5070 84532 5122
rect 84476 5068 84532 5070
rect 82236 5010 82292 5012
rect 82236 4958 82238 5010
rect 82238 4958 82290 5010
rect 82290 4958 82292 5010
rect 82236 4956 82292 4958
rect 81788 3836 81844 3892
rect 80332 3666 80388 3668
rect 80332 3614 80334 3666
rect 80334 3614 80386 3666
rect 80386 3614 80388 3666
rect 80332 3612 80388 3614
rect 81004 3388 81060 3444
rect 82908 3442 82964 3444
rect 82908 3390 82910 3442
rect 82910 3390 82962 3442
rect 82962 3390 82964 3442
rect 82908 3388 82964 3390
rect 86492 14252 86548 14308
rect 88620 34242 88676 34244
rect 88620 34190 88622 34242
rect 88622 34190 88674 34242
rect 88674 34190 88676 34242
rect 88620 34188 88676 34190
rect 89068 36482 89124 36484
rect 89068 36430 89070 36482
rect 89070 36430 89122 36482
rect 89122 36430 89124 36482
rect 89068 36428 89124 36430
rect 89180 36316 89236 36372
rect 88956 35196 89012 35252
rect 88844 33516 88900 33572
rect 88956 34524 89012 34580
rect 89068 33458 89124 33460
rect 89068 33406 89070 33458
rect 89070 33406 89122 33458
rect 89122 33406 89124 33458
rect 89068 33404 89124 33406
rect 89516 36316 89572 36372
rect 89628 34690 89684 34692
rect 89628 34638 89630 34690
rect 89630 34638 89682 34690
rect 89682 34638 89684 34690
rect 89628 34636 89684 34638
rect 89852 36316 89908 36372
rect 90188 36204 90244 36260
rect 89964 35644 90020 35700
rect 90412 35644 90468 35700
rect 90300 35196 90356 35252
rect 88956 28028 89012 28084
rect 89516 24892 89572 24948
rect 89628 33964 89684 34020
rect 91420 36988 91476 37044
rect 90748 36370 90804 36372
rect 90748 36318 90750 36370
rect 90750 36318 90802 36370
rect 90802 36318 90804 36370
rect 90748 36316 90804 36318
rect 90524 34524 90580 34580
rect 90300 34300 90356 34356
rect 90412 34242 90468 34244
rect 90412 34190 90414 34242
rect 90414 34190 90466 34242
rect 90466 34190 90468 34242
rect 90412 34188 90468 34190
rect 90076 32620 90132 32676
rect 89740 27132 89796 27188
rect 90748 35196 90804 35252
rect 90860 34076 90916 34132
rect 91196 35644 91252 35700
rect 91084 34018 91140 34020
rect 91084 33966 91086 34018
rect 91086 33966 91138 34018
rect 91138 33966 91140 34018
rect 91084 33964 91140 33966
rect 90748 33516 90804 33572
rect 91308 35084 91364 35140
rect 91532 35084 91588 35140
rect 91308 34524 91364 34580
rect 89628 24444 89684 24500
rect 89404 23100 89460 23156
rect 88620 15932 88676 15988
rect 87612 7196 87668 7252
rect 85596 6412 85652 6468
rect 85484 5122 85540 5124
rect 85484 5070 85486 5122
rect 85486 5070 85538 5122
rect 85538 5070 85540 5122
rect 85484 5068 85540 5070
rect 87388 6130 87444 6132
rect 87388 6078 87390 6130
rect 87390 6078 87442 6130
rect 87442 6078 87444 6130
rect 87388 6076 87444 6078
rect 88172 6578 88228 6580
rect 88172 6526 88174 6578
rect 88174 6526 88226 6578
rect 88226 6526 88228 6578
rect 88172 6524 88228 6526
rect 88508 6130 88564 6132
rect 88508 6078 88510 6130
rect 88510 6078 88562 6130
rect 88562 6078 88564 6130
rect 88508 6076 88564 6078
rect 88396 5180 88452 5236
rect 86268 4956 86324 5012
rect 86828 4450 86884 4452
rect 86828 4398 86830 4450
rect 86830 4398 86882 4450
rect 86882 4398 86884 4450
rect 86828 4396 86884 4398
rect 88508 4396 88564 4452
rect 86268 4284 86324 4340
rect 84028 3442 84084 3444
rect 84028 3390 84030 3442
rect 84030 3390 84082 3442
rect 84082 3390 84084 3442
rect 84028 3388 84084 3390
rect 85036 3388 85092 3444
rect 86828 3442 86884 3444
rect 86828 3390 86830 3442
rect 86830 3390 86882 3442
rect 86882 3390 86884 3442
rect 86828 3388 86884 3390
rect 91644 32674 91700 32676
rect 91644 32622 91646 32674
rect 91646 32622 91698 32674
rect 91698 32622 91700 32674
rect 91644 32620 91700 32622
rect 92092 35586 92148 35588
rect 92092 35534 92094 35586
rect 92094 35534 92146 35586
rect 92146 35534 92148 35586
rect 92092 35532 92148 35534
rect 91868 33964 91924 34020
rect 92764 36988 92820 37044
rect 93324 36988 93380 37044
rect 93262 36874 93318 36876
rect 93262 36822 93264 36874
rect 93264 36822 93316 36874
rect 93316 36822 93318 36874
rect 93262 36820 93318 36822
rect 93366 36874 93422 36876
rect 93366 36822 93368 36874
rect 93368 36822 93420 36874
rect 93420 36822 93422 36874
rect 93366 36820 93422 36822
rect 93470 36874 93526 36876
rect 93470 36822 93472 36874
rect 93472 36822 93524 36874
rect 93524 36822 93526 36874
rect 93470 36820 93526 36822
rect 93660 36764 93716 36820
rect 92428 35868 92484 35924
rect 93660 36204 93716 36260
rect 92428 34524 92484 34580
rect 92316 34188 92372 34244
rect 91980 32562 92036 32564
rect 91980 32510 91982 32562
rect 91982 32510 92034 32562
rect 92034 32510 92036 32562
rect 91980 32508 92036 32510
rect 91756 32396 91812 32452
rect 92428 34076 92484 34132
rect 92204 29260 92260 29316
rect 92764 35196 92820 35252
rect 92652 27692 92708 27748
rect 92988 35868 93044 35924
rect 92988 34860 93044 34916
rect 92876 24780 92932 24836
rect 93262 35306 93318 35308
rect 93262 35254 93264 35306
rect 93264 35254 93316 35306
rect 93316 35254 93318 35306
rect 93262 35252 93318 35254
rect 93366 35306 93422 35308
rect 93366 35254 93368 35306
rect 93368 35254 93420 35306
rect 93420 35254 93422 35306
rect 93366 35252 93422 35254
rect 93470 35306 93526 35308
rect 93470 35254 93472 35306
rect 93472 35254 93524 35306
rect 93524 35254 93526 35306
rect 93470 35252 93526 35254
rect 93324 35084 93380 35140
rect 93262 33738 93318 33740
rect 93262 33686 93264 33738
rect 93264 33686 93316 33738
rect 93316 33686 93318 33738
rect 93262 33684 93318 33686
rect 93366 33738 93422 33740
rect 93366 33686 93368 33738
rect 93368 33686 93420 33738
rect 93420 33686 93422 33738
rect 93366 33684 93422 33686
rect 93470 33738 93526 33740
rect 93470 33686 93472 33738
rect 93472 33686 93524 33738
rect 93524 33686 93526 33738
rect 93470 33684 93526 33686
rect 93772 35644 93828 35700
rect 93772 34354 93828 34356
rect 93772 34302 93774 34354
rect 93774 34302 93826 34354
rect 93826 34302 93828 34354
rect 93772 34300 93828 34302
rect 94332 37324 94388 37380
rect 94332 35868 94388 35924
rect 94556 36876 94612 36932
rect 94220 35084 94276 35140
rect 93996 33404 94052 33460
rect 94108 33628 94164 33684
rect 93548 32396 93604 32452
rect 93996 33068 94052 33124
rect 93262 32170 93318 32172
rect 93262 32118 93264 32170
rect 93264 32118 93316 32170
rect 93316 32118 93318 32170
rect 93262 32116 93318 32118
rect 93366 32170 93422 32172
rect 93366 32118 93368 32170
rect 93368 32118 93420 32170
rect 93420 32118 93422 32170
rect 93366 32116 93422 32118
rect 93470 32170 93526 32172
rect 93470 32118 93472 32170
rect 93472 32118 93524 32170
rect 93524 32118 93526 32170
rect 93470 32116 93526 32118
rect 93996 31612 94052 31668
rect 93262 30602 93318 30604
rect 93262 30550 93264 30602
rect 93264 30550 93316 30602
rect 93316 30550 93318 30602
rect 93262 30548 93318 30550
rect 93366 30602 93422 30604
rect 93366 30550 93368 30602
rect 93368 30550 93420 30602
rect 93420 30550 93422 30602
rect 93366 30548 93422 30550
rect 93470 30602 93526 30604
rect 93470 30550 93472 30602
rect 93472 30550 93524 30602
rect 93524 30550 93526 30602
rect 93470 30548 93526 30550
rect 93262 29034 93318 29036
rect 93262 28982 93264 29034
rect 93264 28982 93316 29034
rect 93316 28982 93318 29034
rect 93262 28980 93318 28982
rect 93366 29034 93422 29036
rect 93366 28982 93368 29034
rect 93368 28982 93420 29034
rect 93420 28982 93422 29034
rect 93366 28980 93422 28982
rect 93470 29034 93526 29036
rect 93470 28982 93472 29034
rect 93472 28982 93524 29034
rect 93524 28982 93526 29034
rect 93470 28980 93526 28982
rect 93262 27466 93318 27468
rect 93262 27414 93264 27466
rect 93264 27414 93316 27466
rect 93316 27414 93318 27466
rect 93262 27412 93318 27414
rect 93366 27466 93422 27468
rect 93366 27414 93368 27466
rect 93368 27414 93420 27466
rect 93420 27414 93422 27466
rect 93366 27412 93422 27414
rect 93470 27466 93526 27468
rect 93470 27414 93472 27466
rect 93472 27414 93524 27466
rect 93524 27414 93526 27466
rect 93470 27412 93526 27414
rect 94220 26236 94276 26292
rect 93262 25898 93318 25900
rect 93262 25846 93264 25898
rect 93264 25846 93316 25898
rect 93316 25846 93318 25898
rect 93262 25844 93318 25846
rect 93366 25898 93422 25900
rect 93366 25846 93368 25898
rect 93368 25846 93420 25898
rect 93420 25846 93422 25898
rect 93366 25844 93422 25846
rect 93470 25898 93526 25900
rect 93470 25846 93472 25898
rect 93472 25846 93524 25898
rect 93524 25846 93526 25898
rect 93470 25844 93526 25846
rect 93262 24330 93318 24332
rect 93262 24278 93264 24330
rect 93264 24278 93316 24330
rect 93316 24278 93318 24330
rect 93262 24276 93318 24278
rect 93366 24330 93422 24332
rect 93366 24278 93368 24330
rect 93368 24278 93420 24330
rect 93420 24278 93422 24330
rect 93366 24276 93422 24278
rect 93470 24330 93526 24332
rect 93470 24278 93472 24330
rect 93472 24278 93524 24330
rect 93524 24278 93526 24330
rect 93470 24276 93526 24278
rect 93262 22762 93318 22764
rect 93262 22710 93264 22762
rect 93264 22710 93316 22762
rect 93316 22710 93318 22762
rect 93262 22708 93318 22710
rect 93366 22762 93422 22764
rect 93366 22710 93368 22762
rect 93368 22710 93420 22762
rect 93420 22710 93422 22762
rect 93366 22708 93422 22710
rect 93470 22762 93526 22764
rect 93470 22710 93472 22762
rect 93472 22710 93524 22762
rect 93524 22710 93526 22762
rect 93470 22708 93526 22710
rect 93262 21194 93318 21196
rect 93262 21142 93264 21194
rect 93264 21142 93316 21194
rect 93316 21142 93318 21194
rect 93262 21140 93318 21142
rect 93366 21194 93422 21196
rect 93366 21142 93368 21194
rect 93368 21142 93420 21194
rect 93420 21142 93422 21194
rect 93366 21140 93422 21142
rect 93470 21194 93526 21196
rect 93470 21142 93472 21194
rect 93472 21142 93524 21194
rect 93524 21142 93526 21194
rect 93470 21140 93526 21142
rect 92988 20076 93044 20132
rect 93262 19626 93318 19628
rect 93262 19574 93264 19626
rect 93264 19574 93316 19626
rect 93316 19574 93318 19626
rect 93262 19572 93318 19574
rect 93366 19626 93422 19628
rect 93366 19574 93368 19626
rect 93368 19574 93420 19626
rect 93420 19574 93422 19626
rect 93366 19572 93422 19574
rect 93470 19626 93526 19628
rect 93470 19574 93472 19626
rect 93472 19574 93524 19626
rect 93524 19574 93526 19626
rect 93470 19572 93526 19574
rect 93262 18058 93318 18060
rect 93262 18006 93264 18058
rect 93264 18006 93316 18058
rect 93316 18006 93318 18058
rect 93262 18004 93318 18006
rect 93366 18058 93422 18060
rect 93366 18006 93368 18058
rect 93368 18006 93420 18058
rect 93420 18006 93422 18058
rect 93366 18004 93422 18006
rect 93470 18058 93526 18060
rect 93470 18006 93472 18058
rect 93472 18006 93524 18058
rect 93524 18006 93526 18058
rect 93470 18004 93526 18006
rect 91420 11116 91476 11172
rect 92428 17612 92484 17668
rect 93262 16490 93318 16492
rect 93262 16438 93264 16490
rect 93264 16438 93316 16490
rect 93316 16438 93318 16490
rect 93262 16436 93318 16438
rect 93366 16490 93422 16492
rect 93366 16438 93368 16490
rect 93368 16438 93420 16490
rect 93420 16438 93422 16490
rect 93366 16436 93422 16438
rect 93470 16490 93526 16492
rect 93470 16438 93472 16490
rect 93472 16438 93524 16490
rect 93524 16438 93526 16490
rect 93470 16436 93526 16438
rect 93262 14922 93318 14924
rect 93262 14870 93264 14922
rect 93264 14870 93316 14922
rect 93316 14870 93318 14922
rect 93262 14868 93318 14870
rect 93366 14922 93422 14924
rect 93366 14870 93368 14922
rect 93368 14870 93420 14922
rect 93420 14870 93422 14922
rect 93366 14868 93422 14870
rect 93470 14922 93526 14924
rect 93470 14870 93472 14922
rect 93472 14870 93524 14922
rect 93524 14870 93526 14922
rect 93470 14868 93526 14870
rect 93262 13354 93318 13356
rect 93262 13302 93264 13354
rect 93264 13302 93316 13354
rect 93316 13302 93318 13354
rect 93262 13300 93318 13302
rect 93366 13354 93422 13356
rect 93366 13302 93368 13354
rect 93368 13302 93420 13354
rect 93420 13302 93422 13354
rect 93366 13300 93422 13302
rect 93470 13354 93526 13356
rect 93470 13302 93472 13354
rect 93472 13302 93524 13354
rect 93524 13302 93526 13354
rect 93470 13300 93526 13302
rect 93262 11786 93318 11788
rect 93262 11734 93264 11786
rect 93264 11734 93316 11786
rect 93316 11734 93318 11786
rect 93262 11732 93318 11734
rect 93366 11786 93422 11788
rect 93366 11734 93368 11786
rect 93368 11734 93420 11786
rect 93420 11734 93422 11786
rect 93366 11732 93422 11734
rect 93470 11786 93526 11788
rect 93470 11734 93472 11786
rect 93472 11734 93524 11786
rect 93524 11734 93526 11786
rect 93470 11732 93526 11734
rect 93262 10218 93318 10220
rect 93262 10166 93264 10218
rect 93264 10166 93316 10218
rect 93316 10166 93318 10218
rect 93262 10164 93318 10166
rect 93366 10218 93422 10220
rect 93366 10166 93368 10218
rect 93368 10166 93420 10218
rect 93420 10166 93422 10218
rect 93366 10164 93422 10166
rect 93470 10218 93526 10220
rect 93470 10166 93472 10218
rect 93472 10166 93524 10218
rect 93524 10166 93526 10218
rect 93470 10164 93526 10166
rect 93262 8650 93318 8652
rect 93262 8598 93264 8650
rect 93264 8598 93316 8650
rect 93316 8598 93318 8650
rect 93262 8596 93318 8598
rect 93366 8650 93422 8652
rect 93366 8598 93368 8650
rect 93368 8598 93420 8650
rect 93420 8598 93422 8650
rect 93366 8596 93422 8598
rect 93470 8650 93526 8652
rect 93470 8598 93472 8650
rect 93472 8598 93524 8650
rect 93524 8598 93526 8650
rect 93470 8596 93526 8598
rect 89740 7420 89796 7476
rect 88956 6524 89012 6580
rect 89068 7308 89124 7364
rect 89180 7196 89236 7252
rect 89628 7196 89684 7252
rect 92540 8316 92596 8372
rect 90860 7698 90916 7700
rect 90860 7646 90862 7698
rect 90862 7646 90914 7698
rect 90914 7646 90916 7698
rect 90860 7644 90916 7646
rect 90860 7420 90916 7476
rect 91420 7362 91476 7364
rect 91420 7310 91422 7362
rect 91422 7310 91474 7362
rect 91474 7310 91476 7362
rect 91420 7308 91476 7310
rect 90412 6860 90468 6916
rect 91196 6914 91252 6916
rect 91196 6862 91198 6914
rect 91198 6862 91250 6914
rect 91250 6862 91252 6914
rect 91196 6860 91252 6862
rect 91980 6690 92036 6692
rect 91980 6638 91982 6690
rect 91982 6638 92034 6690
rect 92034 6638 92036 6690
rect 91980 6636 92036 6638
rect 91868 6578 91924 6580
rect 91868 6526 91870 6578
rect 91870 6526 91922 6578
rect 91922 6526 91924 6578
rect 91868 6524 91924 6526
rect 90076 6076 90132 6132
rect 89404 5234 89460 5236
rect 89404 5182 89406 5234
rect 89406 5182 89458 5234
rect 89458 5182 89460 5234
rect 89404 5180 89460 5182
rect 89516 4620 89572 4676
rect 89180 4338 89236 4340
rect 89180 4286 89182 4338
rect 89182 4286 89234 4338
rect 89234 4286 89236 4338
rect 89180 4284 89236 4286
rect 90412 6130 90468 6132
rect 90412 6078 90414 6130
rect 90414 6078 90466 6130
rect 90466 6078 90468 6130
rect 90412 6076 90468 6078
rect 91868 6018 91924 6020
rect 91868 5966 91870 6018
rect 91870 5966 91922 6018
rect 91922 5966 91924 6018
rect 91868 5964 91924 5966
rect 90972 5906 91028 5908
rect 90972 5854 90974 5906
rect 90974 5854 91026 5906
rect 91026 5854 91028 5906
rect 90972 5852 91028 5854
rect 91980 5852 92036 5908
rect 90748 5180 90804 5236
rect 91644 5234 91700 5236
rect 91644 5182 91646 5234
rect 91646 5182 91698 5234
rect 91698 5182 91700 5234
rect 91644 5180 91700 5182
rect 92204 5234 92260 5236
rect 92204 5182 92206 5234
rect 92206 5182 92258 5234
rect 92258 5182 92260 5234
rect 92204 5180 92260 5182
rect 91084 5010 91140 5012
rect 91084 4958 91086 5010
rect 91086 4958 91138 5010
rect 91138 4958 91140 5010
rect 91084 4956 91140 4958
rect 92428 4956 92484 5012
rect 90748 4620 90804 4676
rect 91756 4172 91812 4228
rect 87948 3442 88004 3444
rect 87948 3390 87950 3442
rect 87950 3390 88002 3442
rect 88002 3390 88004 3442
rect 87948 3388 88004 3390
rect 89068 3388 89124 3444
rect 91084 3442 91140 3444
rect 91084 3390 91086 3442
rect 91086 3390 91138 3442
rect 91138 3390 91140 3442
rect 91084 3388 91140 3390
rect 94780 35532 94836 35588
rect 94556 33628 94612 33684
rect 94780 33122 94836 33124
rect 94780 33070 94782 33122
rect 94782 33070 94834 33122
rect 94834 33070 94836 33122
rect 94780 33068 94836 33070
rect 96236 36652 96292 36708
rect 96012 36316 96068 36372
rect 96460 36092 96516 36148
rect 95116 35196 95172 35252
rect 95564 35644 95620 35700
rect 95788 35084 95844 35140
rect 95900 34860 95956 34916
rect 96460 35308 96516 35364
rect 95116 33292 95172 33348
rect 95228 33458 95284 33460
rect 95228 33406 95230 33458
rect 95230 33406 95282 33458
rect 95282 33406 95284 33458
rect 95228 33404 95284 33406
rect 95004 33068 95060 33124
rect 97468 36370 97524 36372
rect 97468 36318 97470 36370
rect 97470 36318 97522 36370
rect 97522 36318 97524 36370
rect 97468 36316 97524 36318
rect 97244 35308 97300 35364
rect 96908 33964 96964 34020
rect 97580 35196 97636 35252
rect 97804 35084 97860 35140
rect 98028 34076 98084 34132
rect 98252 35756 98308 35812
rect 97916 34018 97972 34020
rect 97916 33966 97918 34018
rect 97918 33966 97970 34018
rect 97970 33966 97972 34018
rect 97916 33964 97972 33966
rect 96012 32732 96068 32788
rect 98700 36428 98756 36484
rect 99036 36370 99092 36372
rect 99036 36318 99038 36370
rect 99038 36318 99090 36370
rect 99090 36318 99092 36370
rect 99036 36316 99092 36318
rect 98700 35810 98756 35812
rect 98700 35758 98702 35810
rect 98702 35758 98754 35810
rect 98754 35758 98756 35810
rect 98700 35756 98756 35758
rect 98588 35698 98644 35700
rect 98588 35646 98590 35698
rect 98590 35646 98642 35698
rect 98642 35646 98644 35698
rect 98588 35644 98644 35646
rect 100156 37212 100212 37268
rect 99372 35474 99428 35476
rect 99372 35422 99374 35474
rect 99374 35422 99426 35474
rect 99426 35422 99428 35474
rect 99372 35420 99428 35422
rect 99260 35084 99316 35140
rect 98812 34860 98868 34916
rect 98588 34748 98644 34804
rect 98924 34748 98980 34804
rect 99484 33964 99540 34020
rect 95228 32508 95284 32564
rect 94892 31612 94948 31668
rect 94332 7644 94388 7700
rect 98252 26236 98308 26292
rect 99036 30940 99092 30996
rect 98588 23324 98644 23380
rect 100380 35980 100436 36036
rect 100828 36428 100884 36484
rect 100492 35084 100548 35140
rect 100940 35698 100996 35700
rect 100940 35646 100942 35698
rect 100942 35646 100994 35698
rect 100994 35646 100996 35698
rect 100940 35644 100996 35646
rect 100492 34018 100548 34020
rect 100492 33966 100494 34018
rect 100494 33966 100546 34018
rect 100546 33966 100548 34018
rect 100492 33964 100548 33966
rect 101612 36540 101668 36596
rect 101388 35196 101444 35252
rect 101500 35980 101556 36036
rect 101164 34914 101220 34916
rect 101164 34862 101166 34914
rect 101166 34862 101218 34914
rect 101218 34862 101220 34914
rect 101164 34860 101220 34862
rect 102172 35980 102228 36036
rect 102060 35420 102116 35476
rect 101612 35196 101668 35252
rect 101836 35084 101892 35140
rect 102396 35420 102452 35476
rect 102620 35420 102676 35476
rect 102396 35196 102452 35252
rect 102732 35196 102788 35252
rect 102284 34748 102340 34804
rect 102620 34242 102676 34244
rect 102620 34190 102622 34242
rect 102622 34190 102674 34242
rect 102674 34190 102676 34242
rect 102620 34188 102676 34190
rect 103628 36482 103684 36484
rect 103628 36430 103630 36482
rect 103630 36430 103682 36482
rect 103682 36430 103684 36482
rect 103628 36428 103684 36430
rect 104748 37772 104804 37828
rect 104076 36316 104132 36372
rect 103740 35698 103796 35700
rect 103740 35646 103742 35698
rect 103742 35646 103794 35698
rect 103794 35646 103796 35698
rect 103740 35644 103796 35646
rect 103628 34748 103684 34804
rect 103180 34412 103236 34468
rect 103180 34188 103236 34244
rect 100268 32732 100324 32788
rect 102396 32732 102452 32788
rect 99708 26348 99764 26404
rect 98252 8316 98308 8372
rect 101836 24332 101892 24388
rect 97244 7532 97300 7588
rect 92876 7308 92932 7364
rect 93262 7082 93318 7084
rect 93262 7030 93264 7082
rect 93264 7030 93316 7082
rect 93316 7030 93318 7082
rect 93262 7028 93318 7030
rect 93366 7082 93422 7084
rect 93366 7030 93368 7082
rect 93368 7030 93420 7082
rect 93420 7030 93422 7082
rect 93366 7028 93422 7030
rect 93470 7082 93526 7084
rect 93470 7030 93472 7082
rect 93472 7030 93524 7082
rect 93524 7030 93526 7082
rect 93470 7028 93526 7030
rect 101724 7644 101780 7700
rect 99484 6914 99540 6916
rect 99484 6862 99486 6914
rect 99486 6862 99538 6914
rect 99538 6862 99540 6914
rect 99484 6860 99540 6862
rect 97132 6748 97188 6804
rect 93100 6690 93156 6692
rect 93100 6638 93102 6690
rect 93102 6638 93154 6690
rect 93154 6638 93156 6690
rect 93100 6636 93156 6638
rect 93660 6524 93716 6580
rect 93262 5514 93318 5516
rect 93262 5462 93264 5514
rect 93264 5462 93316 5514
rect 93316 5462 93318 5514
rect 93262 5460 93318 5462
rect 93366 5514 93422 5516
rect 93366 5462 93368 5514
rect 93368 5462 93420 5514
rect 93420 5462 93422 5514
rect 93366 5460 93422 5462
rect 93470 5514 93526 5516
rect 93470 5462 93472 5514
rect 93472 5462 93524 5514
rect 93524 5462 93526 5514
rect 93470 5460 93526 5462
rect 95564 5964 95620 6020
rect 93660 5292 93716 5348
rect 93100 5234 93156 5236
rect 93100 5182 93102 5234
rect 93102 5182 93154 5234
rect 93154 5182 93156 5234
rect 93100 5180 93156 5182
rect 94556 5180 94612 5236
rect 93660 4956 93716 5012
rect 94220 5010 94276 5012
rect 94220 4958 94222 5010
rect 94222 4958 94274 5010
rect 94274 4958 94276 5010
rect 94220 4956 94276 4958
rect 94892 5068 94948 5124
rect 95228 5122 95284 5124
rect 95228 5070 95230 5122
rect 95230 5070 95282 5122
rect 95282 5070 95284 5122
rect 95228 5068 95284 5070
rect 98476 6690 98532 6692
rect 98476 6638 98478 6690
rect 98478 6638 98530 6690
rect 98530 6638 98532 6690
rect 98476 6636 98532 6638
rect 98700 5346 98756 5348
rect 98700 5294 98702 5346
rect 98702 5294 98754 5346
rect 98754 5294 98756 5346
rect 98700 5292 98756 5294
rect 93436 4226 93492 4228
rect 93436 4174 93438 4226
rect 93438 4174 93490 4226
rect 93490 4174 93492 4226
rect 93436 4172 93492 4174
rect 93262 3946 93318 3948
rect 93262 3894 93264 3946
rect 93264 3894 93316 3946
rect 93316 3894 93318 3946
rect 93262 3892 93318 3894
rect 93366 3946 93422 3948
rect 93366 3894 93368 3946
rect 93368 3894 93420 3946
rect 93420 3894 93422 3946
rect 93366 3892 93422 3894
rect 93470 3946 93526 3948
rect 93470 3894 93472 3946
rect 93472 3894 93524 3946
rect 93524 3894 93526 3946
rect 93470 3892 93526 3894
rect 97804 5180 97860 5236
rect 98364 5180 98420 5236
rect 99036 4338 99092 4340
rect 99036 4286 99038 4338
rect 99038 4286 99090 4338
rect 99090 4286 99092 4338
rect 99036 4284 99092 4286
rect 99484 4338 99540 4340
rect 99484 4286 99486 4338
rect 99486 4286 99538 4338
rect 99538 4286 99540 4338
rect 99484 4284 99540 4286
rect 100268 7308 100324 7364
rect 100268 6690 100324 6692
rect 100268 6638 100270 6690
rect 100270 6638 100322 6690
rect 100322 6638 100324 6690
rect 100268 6636 100324 6638
rect 101052 6860 101108 6916
rect 100044 4508 100100 4564
rect 94556 3836 94612 3892
rect 91868 3442 91924 3444
rect 91868 3390 91870 3442
rect 91870 3390 91922 3442
rect 91922 3390 91924 3442
rect 91868 3388 91924 3390
rect 93100 3388 93156 3444
rect 94668 3442 94724 3444
rect 94668 3390 94670 3442
rect 94670 3390 94722 3442
rect 94722 3390 94724 3442
rect 94668 3388 94724 3390
rect 95900 3836 95956 3892
rect 98812 3666 98868 3668
rect 98812 3614 98814 3666
rect 98814 3614 98866 3666
rect 98866 3614 98868 3666
rect 98812 3612 98868 3614
rect 96236 3442 96292 3444
rect 96236 3390 96238 3442
rect 96238 3390 96290 3442
rect 96290 3390 96292 3442
rect 96236 3388 96292 3390
rect 101612 4396 101668 4452
rect 102732 31276 102788 31332
rect 102396 22652 102452 22708
rect 103852 34412 103908 34468
rect 104076 35420 104132 35476
rect 104748 34748 104804 34804
rect 104860 36204 104916 36260
rect 105756 37660 105812 37716
rect 105644 37212 105700 37268
rect 105308 36370 105364 36372
rect 105308 36318 105310 36370
rect 105310 36318 105362 36370
rect 105362 36318 105364 36370
rect 105308 36316 105364 36318
rect 105084 35980 105140 36036
rect 105532 35698 105588 35700
rect 105532 35646 105534 35698
rect 105534 35646 105586 35698
rect 105586 35646 105588 35698
rect 105532 35644 105588 35646
rect 104972 33964 105028 34020
rect 105196 34524 105252 34580
rect 105420 34188 105476 34244
rect 105756 36428 105812 36484
rect 106316 36258 106372 36260
rect 106316 36206 106318 36258
rect 106318 36206 106370 36258
rect 106370 36206 106372 36258
rect 106316 36204 106372 36206
rect 105868 35756 105924 35812
rect 106092 35308 106148 35364
rect 106092 34802 106148 34804
rect 106092 34750 106094 34802
rect 106094 34750 106146 34802
rect 106146 34750 106148 34802
rect 106092 34748 106148 34750
rect 105868 34018 105924 34020
rect 105868 33966 105870 34018
rect 105870 33966 105922 34018
rect 105922 33966 105924 34018
rect 105868 33964 105924 33966
rect 105644 33740 105700 33796
rect 104300 30044 104356 30100
rect 103740 12684 103796 12740
rect 104972 28588 105028 28644
rect 101948 5234 102004 5236
rect 101948 5182 101950 5234
rect 101950 5182 102002 5234
rect 102002 5182 102004 5234
rect 101948 5180 102004 5182
rect 102508 5234 102564 5236
rect 102508 5182 102510 5234
rect 102510 5182 102562 5234
rect 102562 5182 102564 5234
rect 102508 5180 102564 5182
rect 102060 4508 102116 4564
rect 102508 4562 102564 4564
rect 102508 4510 102510 4562
rect 102510 4510 102562 4562
rect 102562 4510 102564 4562
rect 102508 4508 102564 4510
rect 103180 4450 103236 4452
rect 103180 4398 103182 4450
rect 103182 4398 103234 4450
rect 103234 4398 103236 4450
rect 103180 4396 103236 4398
rect 101836 3612 101892 3668
rect 102844 3666 102900 3668
rect 102844 3614 102846 3666
rect 102846 3614 102898 3666
rect 102898 3614 102900 3666
rect 102844 3612 102900 3614
rect 106316 34188 106372 34244
rect 106652 34188 106708 34244
rect 106988 37100 107044 37156
rect 106876 35084 106932 35140
rect 106764 33964 106820 34020
rect 106876 33516 106932 33572
rect 107884 37884 107940 37940
rect 107660 36316 107716 36372
rect 107100 35810 107156 35812
rect 107100 35758 107102 35810
rect 107102 35758 107154 35810
rect 107154 35758 107156 35810
rect 107100 35756 107156 35758
rect 107436 35084 107492 35140
rect 106652 32956 106708 33012
rect 105756 32284 105812 32340
rect 105756 28588 105812 28644
rect 105420 23212 105476 23268
rect 106652 26124 106708 26180
rect 105756 7084 105812 7140
rect 104972 3612 105028 3668
rect 107436 34412 107492 34468
rect 107660 34018 107716 34020
rect 107660 33966 107662 34018
rect 107662 33966 107714 34018
rect 107714 33966 107716 34018
rect 107660 33964 107716 33966
rect 107884 33964 107940 34020
rect 107660 33516 107716 33572
rect 107548 31500 107604 31556
rect 107548 24332 107604 24388
rect 108444 35308 108500 35364
rect 108892 36370 108948 36372
rect 108892 36318 108894 36370
rect 108894 36318 108946 36370
rect 108946 36318 108948 36370
rect 108892 36316 108948 36318
rect 108892 35810 108948 35812
rect 108892 35758 108894 35810
rect 108894 35758 108946 35810
rect 108946 35758 108948 35810
rect 108892 35756 108948 35758
rect 108556 35084 108612 35140
rect 109452 35756 109508 35812
rect 109676 38444 109732 38500
rect 109900 36428 109956 36484
rect 110124 35756 110180 35812
rect 109788 35084 109844 35140
rect 109004 34300 109060 34356
rect 109564 34354 109620 34356
rect 109564 34302 109566 34354
rect 109566 34302 109618 34354
rect 109618 34302 109620 34354
rect 109564 34300 109620 34302
rect 109228 34076 109284 34132
rect 110348 35084 110404 35140
rect 110572 36988 110628 37044
rect 110236 34076 110292 34132
rect 110460 34130 110516 34132
rect 110460 34078 110462 34130
rect 110462 34078 110514 34130
rect 110514 34078 110516 34130
rect 110460 34076 110516 34078
rect 108668 34018 108724 34020
rect 108668 33966 108670 34018
rect 108670 33966 108722 34018
rect 108722 33966 108724 34018
rect 108668 33964 108724 33966
rect 108220 33292 108276 33348
rect 107996 31948 108052 32004
rect 107884 22988 107940 23044
rect 108556 24444 108612 24500
rect 108556 12684 108612 12740
rect 111580 37996 111636 38052
rect 111244 36316 111300 36372
rect 110684 36258 110740 36260
rect 110684 36206 110686 36258
rect 110686 36206 110738 36258
rect 110738 36206 110740 36258
rect 110684 36204 110740 36206
rect 111672 36090 111728 36092
rect 111672 36038 111674 36090
rect 111674 36038 111726 36090
rect 111726 36038 111728 36090
rect 111672 36036 111728 36038
rect 111776 36090 111832 36092
rect 111776 36038 111778 36090
rect 111778 36038 111830 36090
rect 111830 36038 111832 36090
rect 111776 36036 111832 36038
rect 111880 36090 111936 36092
rect 111880 36038 111882 36090
rect 111882 36038 111934 36090
rect 111934 36038 111936 36090
rect 111880 36036 111936 36038
rect 111356 35868 111412 35924
rect 110908 35810 110964 35812
rect 110908 35758 110910 35810
rect 110910 35758 110962 35810
rect 110962 35758 110964 35810
rect 110908 35756 110964 35758
rect 110908 35420 110964 35476
rect 110908 34354 110964 34356
rect 110908 34302 110910 34354
rect 110910 34302 110962 34354
rect 110962 34302 110964 34354
rect 110908 34300 110964 34302
rect 111692 35868 111748 35924
rect 112028 35196 112084 35252
rect 111580 35084 111636 35140
rect 111672 34522 111728 34524
rect 111672 34470 111674 34522
rect 111674 34470 111726 34522
rect 111726 34470 111728 34522
rect 111672 34468 111728 34470
rect 111776 34522 111832 34524
rect 111776 34470 111778 34522
rect 111778 34470 111830 34522
rect 111830 34470 111832 34522
rect 111776 34468 111832 34470
rect 111880 34522 111936 34524
rect 111880 34470 111882 34522
rect 111882 34470 111934 34522
rect 111934 34470 111936 34522
rect 111880 34468 111936 34470
rect 111916 34188 111972 34244
rect 110572 33852 110628 33908
rect 111916 33852 111972 33908
rect 112028 33740 112084 33796
rect 112588 36370 112644 36372
rect 112588 36318 112590 36370
rect 112590 36318 112642 36370
rect 112642 36318 112644 36370
rect 112588 36316 112644 36318
rect 113260 38668 113316 38724
rect 113036 35756 113092 35812
rect 113148 37548 113204 37604
rect 112140 33516 112196 33572
rect 112476 34018 112532 34020
rect 112476 33966 112478 34018
rect 112478 33966 112530 34018
rect 112530 33966 112532 34018
rect 112476 33964 112532 33966
rect 112364 33346 112420 33348
rect 112364 33294 112366 33346
rect 112366 33294 112418 33346
rect 112418 33294 112420 33346
rect 112364 33292 112420 33294
rect 111672 32954 111728 32956
rect 111672 32902 111674 32954
rect 111674 32902 111726 32954
rect 111726 32902 111728 32954
rect 111672 32900 111728 32902
rect 111776 32954 111832 32956
rect 111776 32902 111778 32954
rect 111778 32902 111830 32954
rect 111830 32902 111832 32954
rect 111776 32900 111832 32902
rect 111880 32954 111936 32956
rect 111880 32902 111882 32954
rect 111882 32902 111934 32954
rect 111934 32902 111936 32954
rect 111880 32900 111936 32902
rect 111672 31386 111728 31388
rect 111672 31334 111674 31386
rect 111674 31334 111726 31386
rect 111726 31334 111728 31386
rect 111672 31332 111728 31334
rect 111776 31386 111832 31388
rect 111776 31334 111778 31386
rect 111778 31334 111830 31386
rect 111830 31334 111832 31386
rect 111776 31332 111832 31334
rect 111880 31386 111936 31388
rect 111880 31334 111882 31386
rect 111882 31334 111934 31386
rect 111934 31334 111936 31386
rect 111880 31332 111936 31334
rect 111672 29818 111728 29820
rect 111672 29766 111674 29818
rect 111674 29766 111726 29818
rect 111726 29766 111728 29818
rect 111672 29764 111728 29766
rect 111776 29818 111832 29820
rect 111776 29766 111778 29818
rect 111778 29766 111830 29818
rect 111830 29766 111832 29818
rect 111776 29764 111832 29766
rect 111880 29818 111936 29820
rect 111880 29766 111882 29818
rect 111882 29766 111934 29818
rect 111934 29766 111936 29818
rect 111880 29764 111936 29766
rect 113484 34524 113540 34580
rect 113372 33964 113428 34020
rect 113148 33852 113204 33908
rect 113036 33516 113092 33572
rect 113932 35868 113988 35924
rect 114380 36370 114436 36372
rect 114380 36318 114382 36370
rect 114382 36318 114434 36370
rect 114434 36318 114436 36370
rect 114380 36316 114436 36318
rect 114828 36316 114884 36372
rect 115052 36092 115108 36148
rect 114268 35810 114324 35812
rect 114268 35758 114270 35810
rect 114270 35758 114322 35810
rect 114322 35758 114324 35810
rect 114268 35756 114324 35758
rect 114044 35084 114100 35140
rect 114828 35196 114884 35252
rect 113820 34914 113876 34916
rect 113820 34862 113822 34914
rect 113822 34862 113874 34914
rect 113874 34862 113876 34914
rect 113820 34860 113876 34862
rect 114604 34860 114660 34916
rect 113820 34242 113876 34244
rect 113820 34190 113822 34242
rect 113822 34190 113874 34242
rect 113874 34190 113876 34242
rect 113820 34188 113876 34190
rect 113820 33740 113876 33796
rect 113596 32284 113652 32340
rect 112476 29484 112532 29540
rect 111672 28250 111728 28252
rect 111672 28198 111674 28250
rect 111674 28198 111726 28250
rect 111726 28198 111728 28250
rect 111672 28196 111728 28198
rect 111776 28250 111832 28252
rect 111776 28198 111778 28250
rect 111778 28198 111830 28250
rect 111830 28198 111832 28250
rect 111776 28196 111832 28198
rect 111880 28250 111936 28252
rect 111880 28198 111882 28250
rect 111882 28198 111934 28250
rect 111934 28198 111936 28250
rect 111880 28196 111936 28198
rect 111672 26682 111728 26684
rect 111672 26630 111674 26682
rect 111674 26630 111726 26682
rect 111726 26630 111728 26682
rect 111672 26628 111728 26630
rect 111776 26682 111832 26684
rect 111776 26630 111778 26682
rect 111778 26630 111830 26682
rect 111830 26630 111832 26682
rect 111776 26628 111832 26630
rect 111880 26682 111936 26684
rect 111880 26630 111882 26682
rect 111882 26630 111934 26682
rect 111934 26630 111936 26682
rect 111880 26628 111936 26630
rect 111672 25114 111728 25116
rect 111672 25062 111674 25114
rect 111674 25062 111726 25114
rect 111726 25062 111728 25114
rect 111672 25060 111728 25062
rect 111776 25114 111832 25116
rect 111776 25062 111778 25114
rect 111778 25062 111830 25114
rect 111830 25062 111832 25114
rect 111776 25060 111832 25062
rect 111880 25114 111936 25116
rect 111880 25062 111882 25114
rect 111882 25062 111934 25114
rect 111934 25062 111936 25114
rect 111880 25060 111936 25062
rect 111672 23546 111728 23548
rect 111672 23494 111674 23546
rect 111674 23494 111726 23546
rect 111726 23494 111728 23546
rect 111672 23492 111728 23494
rect 111776 23546 111832 23548
rect 111776 23494 111778 23546
rect 111778 23494 111830 23546
rect 111830 23494 111832 23546
rect 111776 23492 111832 23494
rect 111880 23546 111936 23548
rect 111880 23494 111882 23546
rect 111882 23494 111934 23546
rect 111934 23494 111936 23546
rect 111880 23492 111936 23494
rect 113260 22652 113316 22708
rect 111672 21978 111728 21980
rect 111672 21926 111674 21978
rect 111674 21926 111726 21978
rect 111726 21926 111728 21978
rect 111672 21924 111728 21926
rect 111776 21978 111832 21980
rect 111776 21926 111778 21978
rect 111778 21926 111830 21978
rect 111830 21926 111832 21978
rect 111776 21924 111832 21926
rect 111880 21978 111936 21980
rect 111880 21926 111882 21978
rect 111882 21926 111934 21978
rect 111934 21926 111936 21978
rect 111880 21924 111936 21926
rect 111672 20410 111728 20412
rect 111672 20358 111674 20410
rect 111674 20358 111726 20410
rect 111726 20358 111728 20410
rect 111672 20356 111728 20358
rect 111776 20410 111832 20412
rect 111776 20358 111778 20410
rect 111778 20358 111830 20410
rect 111830 20358 111832 20410
rect 111776 20356 111832 20358
rect 111880 20410 111936 20412
rect 111880 20358 111882 20410
rect 111882 20358 111934 20410
rect 111934 20358 111936 20410
rect 111880 20356 111936 20358
rect 111672 18842 111728 18844
rect 111672 18790 111674 18842
rect 111674 18790 111726 18842
rect 111726 18790 111728 18842
rect 111672 18788 111728 18790
rect 111776 18842 111832 18844
rect 111776 18790 111778 18842
rect 111778 18790 111830 18842
rect 111830 18790 111832 18842
rect 111776 18788 111832 18790
rect 111880 18842 111936 18844
rect 111880 18790 111882 18842
rect 111882 18790 111934 18842
rect 111934 18790 111936 18842
rect 111880 18788 111936 18790
rect 111672 17274 111728 17276
rect 111672 17222 111674 17274
rect 111674 17222 111726 17274
rect 111726 17222 111728 17274
rect 111672 17220 111728 17222
rect 111776 17274 111832 17276
rect 111776 17222 111778 17274
rect 111778 17222 111830 17274
rect 111830 17222 111832 17274
rect 111776 17220 111832 17222
rect 111880 17274 111936 17276
rect 111880 17222 111882 17274
rect 111882 17222 111934 17274
rect 111934 17222 111936 17274
rect 111880 17220 111936 17222
rect 111672 15706 111728 15708
rect 111672 15654 111674 15706
rect 111674 15654 111726 15706
rect 111726 15654 111728 15706
rect 111672 15652 111728 15654
rect 111776 15706 111832 15708
rect 111776 15654 111778 15706
rect 111778 15654 111830 15706
rect 111830 15654 111832 15706
rect 111776 15652 111832 15654
rect 111880 15706 111936 15708
rect 111880 15654 111882 15706
rect 111882 15654 111934 15706
rect 111934 15654 111936 15706
rect 111880 15652 111936 15654
rect 111672 14138 111728 14140
rect 111672 14086 111674 14138
rect 111674 14086 111726 14138
rect 111726 14086 111728 14138
rect 111672 14084 111728 14086
rect 111776 14138 111832 14140
rect 111776 14086 111778 14138
rect 111778 14086 111830 14138
rect 111830 14086 111832 14138
rect 111776 14084 111832 14086
rect 111880 14138 111936 14140
rect 111880 14086 111882 14138
rect 111882 14086 111934 14138
rect 111934 14086 111936 14138
rect 111880 14084 111936 14086
rect 111672 12570 111728 12572
rect 111672 12518 111674 12570
rect 111674 12518 111726 12570
rect 111726 12518 111728 12570
rect 111672 12516 111728 12518
rect 111776 12570 111832 12572
rect 111776 12518 111778 12570
rect 111778 12518 111830 12570
rect 111830 12518 111832 12570
rect 111776 12516 111832 12518
rect 111880 12570 111936 12572
rect 111880 12518 111882 12570
rect 111882 12518 111934 12570
rect 111934 12518 111936 12570
rect 111880 12516 111936 12518
rect 111672 11002 111728 11004
rect 111672 10950 111674 11002
rect 111674 10950 111726 11002
rect 111726 10950 111728 11002
rect 111672 10948 111728 10950
rect 111776 11002 111832 11004
rect 111776 10950 111778 11002
rect 111778 10950 111830 11002
rect 111830 10950 111832 11002
rect 111776 10948 111832 10950
rect 111880 11002 111936 11004
rect 111880 10950 111882 11002
rect 111882 10950 111934 11002
rect 111934 10950 111936 11002
rect 111880 10948 111936 10950
rect 111672 9434 111728 9436
rect 111672 9382 111674 9434
rect 111674 9382 111726 9434
rect 111726 9382 111728 9434
rect 111672 9380 111728 9382
rect 111776 9434 111832 9436
rect 111776 9382 111778 9434
rect 111778 9382 111830 9434
rect 111830 9382 111832 9434
rect 111776 9380 111832 9382
rect 111880 9434 111936 9436
rect 111880 9382 111882 9434
rect 111882 9382 111934 9434
rect 111934 9382 111936 9434
rect 111880 9380 111936 9382
rect 110460 8652 110516 8708
rect 110460 8428 110516 8484
rect 107212 6076 107268 6132
rect 107884 6130 107940 6132
rect 107884 6078 107886 6130
rect 107886 6078 107938 6130
rect 107938 6078 107940 6130
rect 107884 6076 107940 6078
rect 107548 5180 107604 5236
rect 107884 5068 107940 5124
rect 108220 5740 108276 5796
rect 108220 5180 108276 5236
rect 108332 4060 108388 4116
rect 110348 6524 110404 6580
rect 108892 6076 108948 6132
rect 109564 5906 109620 5908
rect 109564 5854 109566 5906
rect 109566 5854 109618 5906
rect 109618 5854 109620 5906
rect 109564 5852 109620 5854
rect 109228 5122 109284 5124
rect 109228 5070 109230 5122
rect 109230 5070 109282 5122
rect 109282 5070 109284 5122
rect 109228 5068 109284 5070
rect 111672 7866 111728 7868
rect 111672 7814 111674 7866
rect 111674 7814 111726 7866
rect 111726 7814 111728 7866
rect 111672 7812 111728 7814
rect 111776 7866 111832 7868
rect 111776 7814 111778 7866
rect 111778 7814 111830 7866
rect 111830 7814 111832 7866
rect 111776 7812 111832 7814
rect 111880 7866 111936 7868
rect 111880 7814 111882 7866
rect 111882 7814 111934 7866
rect 111934 7814 111936 7866
rect 111880 7812 111936 7814
rect 113036 6636 113092 6692
rect 111580 6524 111636 6580
rect 110460 6076 110516 6132
rect 111672 6298 111728 6300
rect 111672 6246 111674 6298
rect 111674 6246 111726 6298
rect 111726 6246 111728 6298
rect 111672 6244 111728 6246
rect 111776 6298 111832 6300
rect 111776 6246 111778 6298
rect 111778 6246 111830 6298
rect 111830 6246 111832 6298
rect 111776 6244 111832 6246
rect 111880 6298 111936 6300
rect 111880 6246 111882 6298
rect 111882 6246 111934 6298
rect 111934 6246 111936 6298
rect 111880 6244 111936 6246
rect 111020 6076 111076 6132
rect 112028 6018 112084 6020
rect 112028 5966 112030 6018
rect 112030 5966 112082 6018
rect 112082 5966 112084 6018
rect 112028 5964 112084 5966
rect 110348 5852 110404 5908
rect 110348 5516 110404 5572
rect 109676 4956 109732 5012
rect 110684 4956 110740 5012
rect 111020 5628 111076 5684
rect 111132 5516 111188 5572
rect 111356 4898 111412 4900
rect 111356 4846 111358 4898
rect 111358 4846 111410 4898
rect 111410 4846 111412 4898
rect 111356 4844 111412 4846
rect 111672 4730 111728 4732
rect 111672 4678 111674 4730
rect 111674 4678 111726 4730
rect 111726 4678 111728 4730
rect 111672 4676 111728 4678
rect 111776 4730 111832 4732
rect 111776 4678 111778 4730
rect 111778 4678 111830 4730
rect 111830 4678 111832 4730
rect 111776 4676 111832 4678
rect 111880 4730 111936 4732
rect 111880 4678 111882 4730
rect 111882 4678 111934 4730
rect 111934 4678 111936 4730
rect 111880 4676 111936 4678
rect 110684 4172 110740 4228
rect 112028 4338 112084 4340
rect 112028 4286 112030 4338
rect 112030 4286 112082 4338
rect 112082 4286 112084 4338
rect 112028 4284 112084 4286
rect 111692 4226 111748 4228
rect 111692 4174 111694 4226
rect 111694 4174 111746 4226
rect 111746 4174 111748 4226
rect 111692 4172 111748 4174
rect 108780 3612 108836 3668
rect 110572 3666 110628 3668
rect 110572 3614 110574 3666
rect 110574 3614 110626 3666
rect 110626 3614 110628 3666
rect 110572 3612 110628 3614
rect 111804 3554 111860 3556
rect 111804 3502 111806 3554
rect 111806 3502 111858 3554
rect 111858 3502 111860 3554
rect 111804 3500 111860 3502
rect 111672 3162 111728 3164
rect 111672 3110 111674 3162
rect 111674 3110 111726 3162
rect 111726 3110 111728 3162
rect 111672 3108 111728 3110
rect 111776 3162 111832 3164
rect 111776 3110 111778 3162
rect 111778 3110 111830 3162
rect 111830 3110 111832 3162
rect 111776 3108 111832 3110
rect 111880 3162 111936 3164
rect 111880 3110 111882 3162
rect 111882 3110 111934 3162
rect 111934 3110 111936 3162
rect 111880 3108 111936 3110
rect 113036 4338 113092 4340
rect 113036 4286 113038 4338
rect 113038 4286 113090 4338
rect 113090 4286 113092 4338
rect 113036 4284 113092 4286
rect 112588 4060 112644 4116
rect 112588 3724 112644 3780
rect 112364 3500 112420 3556
rect 114156 34130 114212 34132
rect 114156 34078 114158 34130
rect 114158 34078 114210 34130
rect 114210 34078 114212 34130
rect 114156 34076 114212 34078
rect 114044 32284 114100 32340
rect 113932 13356 113988 13412
rect 115388 35980 115444 36036
rect 115052 34076 115108 34132
rect 115612 35644 115668 35700
rect 115500 35084 115556 35140
rect 115388 34860 115444 34916
rect 115276 34636 115332 34692
rect 116508 36370 116564 36372
rect 116508 36318 116510 36370
rect 116510 36318 116562 36370
rect 116562 36318 116564 36370
rect 116508 36316 116564 36318
rect 116060 35810 116116 35812
rect 116060 35758 116062 35810
rect 116062 35758 116114 35810
rect 116114 35758 116116 35810
rect 116060 35756 116116 35758
rect 115948 35644 116004 35700
rect 117180 37436 117236 37492
rect 116620 35084 116676 35140
rect 115724 33964 115780 34020
rect 116620 34018 116676 34020
rect 116620 33966 116622 34018
rect 116622 33966 116674 34018
rect 116674 33966 116676 34018
rect 116620 33964 116676 33966
rect 117068 35084 117124 35140
rect 116956 34690 117012 34692
rect 116956 34638 116958 34690
rect 116958 34638 117010 34690
rect 117010 34638 117012 34690
rect 116956 34636 117012 34638
rect 117628 38332 117684 38388
rect 117628 37100 117684 37156
rect 118412 36652 118468 36708
rect 119196 37100 119252 37156
rect 117292 35196 117348 35252
rect 117180 34300 117236 34356
rect 116844 32620 116900 32676
rect 118300 36370 118356 36372
rect 118300 36318 118302 36370
rect 118302 36318 118354 36370
rect 118354 36318 118356 36370
rect 118300 36316 118356 36318
rect 117852 35084 117908 35140
rect 118412 35196 118468 35252
rect 119084 34524 119140 34580
rect 117740 34354 117796 34356
rect 117740 34302 117742 34354
rect 117742 34302 117794 34354
rect 117794 34302 117796 34354
rect 117740 34300 117796 34302
rect 118524 33516 118580 33572
rect 119420 36594 119476 36596
rect 119420 36542 119422 36594
rect 119422 36542 119474 36594
rect 119474 36542 119476 36594
rect 119420 36540 119476 36542
rect 120092 36204 120148 36260
rect 119868 35474 119924 35476
rect 119868 35422 119870 35474
rect 119870 35422 119922 35474
rect 119922 35422 119924 35474
rect 119868 35420 119924 35422
rect 119420 35084 119476 35140
rect 119980 35084 120036 35140
rect 119420 34748 119476 34804
rect 115612 32508 115668 32564
rect 117852 33180 117908 33236
rect 118412 33234 118468 33236
rect 118412 33182 118414 33234
rect 118414 33182 118466 33234
rect 118466 33182 118468 33234
rect 118412 33180 118468 33182
rect 118748 33234 118804 33236
rect 118748 33182 118750 33234
rect 118750 33182 118802 33234
rect 118802 33182 118804 33234
rect 118748 33180 118804 33182
rect 118748 32450 118804 32452
rect 118748 32398 118750 32450
rect 118750 32398 118802 32450
rect 118802 32398 118804 32450
rect 118748 32396 118804 32398
rect 118972 32396 119028 32452
rect 119084 33516 119140 33572
rect 119084 33292 119140 33348
rect 119196 31724 119252 31780
rect 119644 33068 119700 33124
rect 120428 36652 120484 36708
rect 120652 36540 120708 36596
rect 120092 33122 120148 33124
rect 120092 33070 120094 33122
rect 120094 33070 120146 33122
rect 120146 33070 120148 33122
rect 120092 33068 120148 33070
rect 117628 26124 117684 26180
rect 117404 22876 117460 22932
rect 115276 20972 115332 21028
rect 115724 13356 115780 13412
rect 113596 8092 113652 8148
rect 113484 6524 113540 6580
rect 114156 6188 114212 6244
rect 114044 5964 114100 6020
rect 115164 8092 115220 8148
rect 114380 6802 114436 6804
rect 114380 6750 114382 6802
rect 114382 6750 114434 6802
rect 114434 6750 114436 6802
rect 114380 6748 114436 6750
rect 120316 35196 120372 35252
rect 120540 35420 120596 35476
rect 121548 37100 121604 37156
rect 121436 36258 121492 36260
rect 121436 36206 121438 36258
rect 121438 36206 121490 36258
rect 121490 36206 121492 36258
rect 121436 36204 121492 36206
rect 121100 35586 121156 35588
rect 121100 35534 121102 35586
rect 121102 35534 121154 35586
rect 121154 35534 121156 35586
rect 121100 35532 121156 35534
rect 121100 35196 121156 35252
rect 120092 26124 120148 26180
rect 119308 24556 119364 24612
rect 122220 36652 122276 36708
rect 120988 26012 121044 26068
rect 121996 36316 122052 36372
rect 122108 35196 122164 35252
rect 122556 35756 122612 35812
rect 122668 35084 122724 35140
rect 123340 36594 123396 36596
rect 123340 36542 123342 36594
rect 123342 36542 123394 36594
rect 123394 36542 123396 36594
rect 123340 36540 123396 36542
rect 123116 35810 123172 35812
rect 123116 35758 123118 35810
rect 123118 35758 123170 35810
rect 123170 35758 123172 35810
rect 123116 35756 123172 35758
rect 125356 38556 125412 38612
rect 124348 36370 124404 36372
rect 124348 36318 124350 36370
rect 124350 36318 124402 36370
rect 124402 36318 124404 36370
rect 124348 36316 124404 36318
rect 123452 35532 123508 35588
rect 122892 33964 122948 34020
rect 124796 35532 124852 35588
rect 123004 35308 123060 35364
rect 124012 35084 124068 35140
rect 124012 34860 124068 34916
rect 121772 22540 121828 22596
rect 119196 9996 119252 10052
rect 115724 6802 115780 6804
rect 115724 6750 115726 6802
rect 115726 6750 115778 6802
rect 115778 6750 115780 6802
rect 115724 6748 115780 6750
rect 115836 8652 115892 8708
rect 115052 6578 115108 6580
rect 115052 6526 115054 6578
rect 115054 6526 115106 6578
rect 115106 6526 115108 6578
rect 115052 6524 115108 6526
rect 115724 6524 115780 6580
rect 114380 5964 114436 6020
rect 113932 5682 113988 5684
rect 113932 5630 113934 5682
rect 113934 5630 113986 5682
rect 113986 5630 113988 5682
rect 113932 5628 113988 5630
rect 115612 6018 115668 6020
rect 115612 5966 115614 6018
rect 115614 5966 115666 6018
rect 115666 5966 115668 6018
rect 115612 5964 115668 5966
rect 115052 5180 115108 5236
rect 113596 4844 113652 4900
rect 119196 8258 119252 8260
rect 119196 8206 119198 8258
rect 119198 8206 119250 8258
rect 119250 8206 119252 8258
rect 119196 8204 119252 8206
rect 122108 15932 122164 15988
rect 122444 26012 122500 26068
rect 120540 8258 120596 8260
rect 120540 8206 120542 8258
rect 120542 8206 120594 8258
rect 120594 8206 120596 8258
rect 120540 8204 120596 8206
rect 120988 9996 121044 10052
rect 118300 8146 118356 8148
rect 118300 8094 118302 8146
rect 118302 8094 118354 8146
rect 118354 8094 118356 8146
rect 118300 8092 118356 8094
rect 119420 8146 119476 8148
rect 119420 8094 119422 8146
rect 119422 8094 119474 8146
rect 119474 8094 119476 8146
rect 119420 8092 119476 8094
rect 116508 6860 116564 6916
rect 116284 6524 116340 6580
rect 116284 6300 116340 6356
rect 117516 7362 117572 7364
rect 117516 7310 117518 7362
rect 117518 7310 117570 7362
rect 117570 7310 117572 7362
rect 117516 7308 117572 7310
rect 116732 6636 116788 6692
rect 116172 5794 116228 5796
rect 116172 5742 116174 5794
rect 116174 5742 116226 5794
rect 116226 5742 116228 5794
rect 116172 5740 116228 5742
rect 115948 5292 116004 5348
rect 116172 5292 116228 5348
rect 116732 5180 116788 5236
rect 115836 4844 115892 4900
rect 115948 4172 116004 4228
rect 114604 3612 114660 3668
rect 113260 3388 113316 3444
rect 114604 3442 114660 3444
rect 114604 3390 114606 3442
rect 114606 3390 114658 3442
rect 114658 3390 114660 3442
rect 114604 3388 114660 3390
rect 115612 3442 115668 3444
rect 115612 3390 115614 3442
rect 115614 3390 115666 3442
rect 115666 3390 115668 3442
rect 115612 3388 115668 3390
rect 117180 5122 117236 5124
rect 117180 5070 117182 5122
rect 117182 5070 117234 5122
rect 117234 5070 117236 5122
rect 117180 5068 117236 5070
rect 117180 4844 117236 4900
rect 119420 7474 119476 7476
rect 119420 7422 119422 7474
rect 119422 7422 119474 7474
rect 119474 7422 119476 7474
rect 119420 7420 119476 7422
rect 119644 7308 119700 7364
rect 119868 6412 119924 6468
rect 119644 5906 119700 5908
rect 119644 5854 119646 5906
rect 119646 5854 119698 5906
rect 119698 5854 119700 5906
rect 119644 5852 119700 5854
rect 119980 5740 120036 5796
rect 119868 5292 119924 5348
rect 119980 4508 120036 4564
rect 117292 4226 117348 4228
rect 117292 4174 117294 4226
rect 117294 4174 117346 4226
rect 117346 4174 117348 4226
rect 117292 4172 117348 4174
rect 118188 4060 118244 4116
rect 120428 4060 120484 4116
rect 119980 3666 120036 3668
rect 119980 3614 119982 3666
rect 119982 3614 120034 3666
rect 120034 3614 120036 3666
rect 119980 3612 120036 3614
rect 121212 7308 121268 7364
rect 121436 8034 121492 8036
rect 121436 7982 121438 8034
rect 121438 7982 121490 8034
rect 121490 7982 121492 8034
rect 121436 7980 121492 7982
rect 123788 34018 123844 34020
rect 123788 33966 123790 34018
rect 123790 33966 123842 34018
rect 123842 33966 123844 34018
rect 123788 33964 123844 33966
rect 125692 36204 125748 36260
rect 125804 35868 125860 35924
rect 125580 35644 125636 35700
rect 123900 33068 123956 33124
rect 123564 31836 123620 31892
rect 124908 33122 124964 33124
rect 124908 33070 124910 33122
rect 124910 33070 124962 33122
rect 124962 33070 124964 33122
rect 124908 33068 124964 33070
rect 126140 36370 126196 36372
rect 126140 36318 126142 36370
rect 126142 36318 126194 36370
rect 126194 36318 126196 36370
rect 126140 36316 126196 36318
rect 127708 36370 127764 36372
rect 127708 36318 127710 36370
rect 127710 36318 127762 36370
rect 127762 36318 127764 36370
rect 127708 36316 127764 36318
rect 127932 36204 127988 36260
rect 126476 35084 126532 35140
rect 125580 32732 125636 32788
rect 126028 33964 126084 34020
rect 124796 26236 124852 26292
rect 122444 7980 122500 8036
rect 125132 26124 125188 26180
rect 121436 7420 121492 7476
rect 121996 7474 122052 7476
rect 121996 7422 121998 7474
rect 121998 7422 122050 7474
rect 122050 7422 122052 7474
rect 121996 7420 122052 7422
rect 123340 7420 123396 7476
rect 122892 7362 122948 7364
rect 122892 7310 122894 7362
rect 122894 7310 122946 7362
rect 122946 7310 122948 7362
rect 122892 7308 122948 7310
rect 121324 6860 121380 6916
rect 121324 6466 121380 6468
rect 121324 6414 121326 6466
rect 121326 6414 121378 6466
rect 121378 6414 121380 6466
rect 121324 6412 121380 6414
rect 120988 5292 121044 5348
rect 121100 5180 121156 5236
rect 120652 3836 120708 3892
rect 121772 5852 121828 5908
rect 125020 6412 125076 6468
rect 124236 4562 124292 4564
rect 124236 4510 124238 4562
rect 124238 4510 124290 4562
rect 124290 4510 124292 4562
rect 124236 4508 124292 4510
rect 124684 4508 124740 4564
rect 117292 3500 117348 3556
rect 116284 3442 116340 3444
rect 116284 3390 116286 3442
rect 116286 3390 116338 3442
rect 116338 3390 116340 3442
rect 116284 3388 116340 3390
rect 118524 3500 118580 3556
rect 119420 3442 119476 3444
rect 119420 3390 119422 3442
rect 119422 3390 119474 3442
rect 119474 3390 119476 3442
rect 119420 3388 119476 3390
rect 120092 3388 120148 3444
rect 127932 35420 127988 35476
rect 127708 35084 127764 35140
rect 127484 34076 127540 34132
rect 127596 34636 127652 34692
rect 126588 33180 126644 33236
rect 128940 36428 128996 36484
rect 128828 34914 128884 34916
rect 128828 34862 128830 34914
rect 128830 34862 128882 34914
rect 128882 34862 128884 34914
rect 128828 34860 128884 34862
rect 129052 35756 129108 35812
rect 129836 36482 129892 36484
rect 129836 36430 129838 36482
rect 129838 36430 129890 36482
rect 129890 36430 129892 36482
rect 129836 36428 129892 36430
rect 129500 35868 129556 35924
rect 127596 30156 127652 30212
rect 126028 25676 126084 25732
rect 126812 27692 126868 27748
rect 126364 11116 126420 11172
rect 129164 35420 129220 35476
rect 129388 34860 129444 34916
rect 129276 34690 129332 34692
rect 129276 34638 129278 34690
rect 129278 34638 129330 34690
rect 129330 34638 129332 34690
rect 129276 34636 129332 34638
rect 130082 36874 130138 36876
rect 130082 36822 130084 36874
rect 130084 36822 130136 36874
rect 130136 36822 130138 36874
rect 130082 36820 130138 36822
rect 130186 36874 130242 36876
rect 130186 36822 130188 36874
rect 130188 36822 130240 36874
rect 130240 36822 130242 36874
rect 130186 36820 130242 36822
rect 130290 36874 130346 36876
rect 130290 36822 130292 36874
rect 130292 36822 130344 36874
rect 130344 36822 130346 36874
rect 130290 36820 130346 36822
rect 130396 36370 130452 36372
rect 130396 36318 130398 36370
rect 130398 36318 130450 36370
rect 130450 36318 130452 36370
rect 130396 36316 130452 36318
rect 130732 35756 130788 35812
rect 130082 35306 130138 35308
rect 130082 35254 130084 35306
rect 130084 35254 130136 35306
rect 130136 35254 130138 35306
rect 130082 35252 130138 35254
rect 130186 35306 130242 35308
rect 130186 35254 130188 35306
rect 130188 35254 130240 35306
rect 130240 35254 130242 35306
rect 130186 35252 130242 35254
rect 130290 35306 130346 35308
rect 130290 35254 130292 35306
rect 130292 35254 130344 35306
rect 130344 35254 130346 35306
rect 130290 35252 130346 35254
rect 130060 34914 130116 34916
rect 130060 34862 130062 34914
rect 130062 34862 130114 34914
rect 130114 34862 130116 34914
rect 130060 34860 130116 34862
rect 129948 34636 130004 34692
rect 129948 34018 130004 34020
rect 129948 33966 129950 34018
rect 129950 33966 130002 34018
rect 130002 33966 130004 34018
rect 129948 33964 130004 33966
rect 130508 34860 130564 34916
rect 130620 33964 130676 34020
rect 130082 33738 130138 33740
rect 130082 33686 130084 33738
rect 130084 33686 130136 33738
rect 130136 33686 130138 33738
rect 130082 33684 130138 33686
rect 130186 33738 130242 33740
rect 130186 33686 130188 33738
rect 130188 33686 130240 33738
rect 130240 33686 130242 33738
rect 130186 33684 130242 33686
rect 130290 33738 130346 33740
rect 130290 33686 130292 33738
rect 130292 33686 130344 33738
rect 130344 33686 130346 33738
rect 130290 33684 130346 33686
rect 130732 33852 130788 33908
rect 131628 36204 131684 36260
rect 131292 34130 131348 34132
rect 131292 34078 131294 34130
rect 131294 34078 131346 34130
rect 131346 34078 131348 34130
rect 131292 34076 131348 34078
rect 131628 35698 131684 35700
rect 131628 35646 131630 35698
rect 131630 35646 131682 35698
rect 131682 35646 131684 35698
rect 131628 35644 131684 35646
rect 132748 36764 132804 36820
rect 132188 35922 132244 35924
rect 132188 35870 132190 35922
rect 132190 35870 132242 35922
rect 132242 35870 132244 35922
rect 132188 35868 132244 35870
rect 131852 35084 131908 35140
rect 132636 35644 132692 35700
rect 131516 34412 131572 34468
rect 131068 32732 131124 32788
rect 132076 34802 132132 34804
rect 132076 34750 132078 34802
rect 132078 34750 132130 34802
rect 132130 34750 132132 34802
rect 132076 34748 132132 34750
rect 131740 34412 131796 34468
rect 132748 35196 132804 35252
rect 130082 32170 130138 32172
rect 130082 32118 130084 32170
rect 130084 32118 130136 32170
rect 130136 32118 130138 32170
rect 130082 32116 130138 32118
rect 130186 32170 130242 32172
rect 130186 32118 130188 32170
rect 130188 32118 130240 32170
rect 130240 32118 130242 32170
rect 130186 32116 130242 32118
rect 130290 32170 130346 32172
rect 130290 32118 130292 32170
rect 130292 32118 130344 32170
rect 130344 32118 130346 32170
rect 130290 32116 130346 32118
rect 131964 33346 132020 33348
rect 131964 33294 131966 33346
rect 131966 33294 132018 33346
rect 132018 33294 132020 33346
rect 131964 33292 132020 33294
rect 132972 34748 133028 34804
rect 132860 33404 132916 33460
rect 132300 33292 132356 33348
rect 131628 31052 131684 31108
rect 130082 30602 130138 30604
rect 130082 30550 130084 30602
rect 130084 30550 130136 30602
rect 130136 30550 130138 30602
rect 130082 30548 130138 30550
rect 130186 30602 130242 30604
rect 130186 30550 130188 30602
rect 130188 30550 130240 30602
rect 130240 30550 130242 30602
rect 130186 30548 130242 30550
rect 130290 30602 130346 30604
rect 130290 30550 130292 30602
rect 130292 30550 130344 30602
rect 130344 30550 130346 30602
rect 130290 30548 130346 30550
rect 130082 29034 130138 29036
rect 130082 28982 130084 29034
rect 130084 28982 130136 29034
rect 130136 28982 130138 29034
rect 130082 28980 130138 28982
rect 130186 29034 130242 29036
rect 130186 28982 130188 29034
rect 130188 28982 130240 29034
rect 130240 28982 130242 29034
rect 130186 28980 130242 28982
rect 130290 29034 130346 29036
rect 130290 28982 130292 29034
rect 130292 28982 130344 29034
rect 130344 28982 130346 29034
rect 130290 28980 130346 28982
rect 133532 35980 133588 36036
rect 133644 35756 133700 35812
rect 133868 36764 133924 36820
rect 135100 36428 135156 36484
rect 134540 36316 134596 36372
rect 135324 36316 135380 36372
rect 133980 36258 134036 36260
rect 133980 36206 133982 36258
rect 133982 36206 134034 36258
rect 134034 36206 134036 36258
rect 133980 36204 134036 36206
rect 133644 35084 133700 35140
rect 133084 28364 133140 28420
rect 130082 27466 130138 27468
rect 130082 27414 130084 27466
rect 130084 27414 130136 27466
rect 130136 27414 130138 27466
rect 130082 27412 130138 27414
rect 130186 27466 130242 27468
rect 130186 27414 130188 27466
rect 130188 27414 130240 27466
rect 130240 27414 130242 27466
rect 130186 27412 130242 27414
rect 130290 27466 130346 27468
rect 130290 27414 130292 27466
rect 130292 27414 130344 27466
rect 130344 27414 130346 27466
rect 130290 27412 130346 27414
rect 133196 26124 133252 26180
rect 130082 25898 130138 25900
rect 130082 25846 130084 25898
rect 130084 25846 130136 25898
rect 130136 25846 130138 25898
rect 130082 25844 130138 25846
rect 130186 25898 130242 25900
rect 130186 25846 130188 25898
rect 130188 25846 130240 25898
rect 130240 25846 130242 25898
rect 130186 25844 130242 25846
rect 130290 25898 130346 25900
rect 130290 25846 130292 25898
rect 130292 25846 130344 25898
rect 130344 25846 130346 25898
rect 130290 25844 130346 25846
rect 130082 24330 130138 24332
rect 130082 24278 130084 24330
rect 130084 24278 130136 24330
rect 130136 24278 130138 24330
rect 130082 24276 130138 24278
rect 130186 24330 130242 24332
rect 130186 24278 130188 24330
rect 130188 24278 130240 24330
rect 130240 24278 130242 24330
rect 130186 24276 130242 24278
rect 130290 24330 130346 24332
rect 130290 24278 130292 24330
rect 130292 24278 130344 24330
rect 130344 24278 130346 24330
rect 130290 24276 130346 24278
rect 130082 22762 130138 22764
rect 130082 22710 130084 22762
rect 130084 22710 130136 22762
rect 130136 22710 130138 22762
rect 130082 22708 130138 22710
rect 130186 22762 130242 22764
rect 130186 22710 130188 22762
rect 130188 22710 130240 22762
rect 130240 22710 130242 22762
rect 130186 22708 130242 22710
rect 130290 22762 130346 22764
rect 130290 22710 130292 22762
rect 130292 22710 130344 22762
rect 130344 22710 130346 22762
rect 130290 22708 130346 22710
rect 133868 34354 133924 34356
rect 133868 34302 133870 34354
rect 133870 34302 133922 34354
rect 133922 34302 133924 34354
rect 133868 34300 133924 34302
rect 134988 35698 135044 35700
rect 134988 35646 134990 35698
rect 134990 35646 135042 35698
rect 135042 35646 135044 35698
rect 134988 35644 135044 35646
rect 134764 35420 134820 35476
rect 136108 36370 136164 36372
rect 136108 36318 136110 36370
rect 136110 36318 136162 36370
rect 136162 36318 136164 36370
rect 136108 36316 136164 36318
rect 135660 35756 135716 35812
rect 137116 36204 137172 36260
rect 137116 35980 137172 36036
rect 137004 35586 137060 35588
rect 137004 35534 137006 35586
rect 137006 35534 137058 35586
rect 137058 35534 137060 35586
rect 137004 35532 137060 35534
rect 136332 35308 136388 35364
rect 136780 35308 136836 35364
rect 135436 35084 135492 35140
rect 136332 35084 136388 35140
rect 136332 34748 136388 34804
rect 135660 34300 135716 34356
rect 135100 33292 135156 33348
rect 137004 34242 137060 34244
rect 137004 34190 137006 34242
rect 137006 34190 137058 34242
rect 137058 34190 137060 34242
rect 137004 34188 137060 34190
rect 138124 36316 138180 36372
rect 137340 34690 137396 34692
rect 137340 34638 137342 34690
rect 137342 34638 137394 34690
rect 137394 34638 137396 34690
rect 137340 34636 137396 34638
rect 137340 34412 137396 34468
rect 138012 36258 138068 36260
rect 138012 36206 138014 36258
rect 138014 36206 138066 36258
rect 138066 36206 138068 36258
rect 138012 36204 138068 36206
rect 139020 36092 139076 36148
rect 138012 35308 138068 35364
rect 138796 35196 138852 35252
rect 140028 36370 140084 36372
rect 140028 36318 140030 36370
rect 140030 36318 140082 36370
rect 140082 36318 140084 36370
rect 140028 36316 140084 36318
rect 139356 35196 139412 35252
rect 139132 35084 139188 35140
rect 138012 34802 138068 34804
rect 138012 34750 138014 34802
rect 138014 34750 138066 34802
rect 138066 34750 138068 34802
rect 138012 34748 138068 34750
rect 138572 34802 138628 34804
rect 138572 34750 138574 34802
rect 138574 34750 138626 34802
rect 138626 34750 138628 34802
rect 138572 34748 138628 34750
rect 138348 34242 138404 34244
rect 138348 34190 138350 34242
rect 138350 34190 138402 34242
rect 138402 34190 138404 34242
rect 138348 34188 138404 34190
rect 137452 34076 137508 34132
rect 137340 33852 137396 33908
rect 137228 33404 137284 33460
rect 138124 33458 138180 33460
rect 138124 33406 138126 33458
rect 138126 33406 138178 33458
rect 138178 33406 138180 33458
rect 138124 33404 138180 33406
rect 137452 33346 137508 33348
rect 137452 33294 137454 33346
rect 137454 33294 137506 33346
rect 137506 33294 137508 33346
rect 137452 33292 137508 33294
rect 139020 34412 139076 34468
rect 139692 34802 139748 34804
rect 139692 34750 139694 34802
rect 139694 34750 139746 34802
rect 139746 34750 139748 34802
rect 139692 34748 139748 34750
rect 140028 34130 140084 34132
rect 140028 34078 140030 34130
rect 140030 34078 140082 34130
rect 140082 34078 140084 34130
rect 140028 34076 140084 34078
rect 139244 33404 139300 33460
rect 137004 26796 137060 26852
rect 138796 33068 138852 33124
rect 135996 24108 136052 24164
rect 133644 21756 133700 21812
rect 134428 21756 134484 21812
rect 130082 21194 130138 21196
rect 130082 21142 130084 21194
rect 130084 21142 130136 21194
rect 130136 21142 130138 21194
rect 130082 21140 130138 21142
rect 130186 21194 130242 21196
rect 130186 21142 130188 21194
rect 130188 21142 130240 21194
rect 130240 21142 130242 21194
rect 130186 21140 130242 21142
rect 130290 21194 130346 21196
rect 130290 21142 130292 21194
rect 130292 21142 130344 21194
rect 130344 21142 130346 21194
rect 130290 21140 130346 21142
rect 128828 12572 128884 12628
rect 126812 9884 126868 9940
rect 128716 9938 128772 9940
rect 128716 9886 128718 9938
rect 128718 9886 128770 9938
rect 128770 9886 128772 9938
rect 128716 9884 128772 9886
rect 128044 9042 128100 9044
rect 128044 8990 128046 9042
rect 128046 8990 128098 9042
rect 128098 8990 128100 9042
rect 128044 8988 128100 8990
rect 126028 7586 126084 7588
rect 126028 7534 126030 7586
rect 126030 7534 126082 7586
rect 126082 7534 126084 7586
rect 126028 7532 126084 7534
rect 127036 7420 127092 7476
rect 128156 7756 128212 7812
rect 128044 7644 128100 7700
rect 128156 7474 128212 7476
rect 128156 7422 128158 7474
rect 128158 7422 128210 7474
rect 128210 7422 128212 7474
rect 128156 7420 128212 7422
rect 126924 6412 126980 6468
rect 126476 6300 126532 6356
rect 125356 4338 125412 4340
rect 125356 4286 125358 4338
rect 125358 4286 125410 4338
rect 125410 4286 125412 4338
rect 125356 4284 125412 4286
rect 123228 3554 123284 3556
rect 123228 3502 123230 3554
rect 123230 3502 123282 3554
rect 123282 3502 123284 3554
rect 123228 3500 123284 3502
rect 121772 3388 121828 3444
rect 122108 3442 122164 3444
rect 122108 3390 122110 3442
rect 122110 3390 122162 3442
rect 122162 3390 122164 3442
rect 122108 3388 122164 3390
rect 123676 3442 123732 3444
rect 123676 3390 123678 3442
rect 123678 3390 123730 3442
rect 123730 3390 123732 3442
rect 123676 3388 123732 3390
rect 124012 3388 124068 3444
rect 127372 6466 127428 6468
rect 127372 6414 127374 6466
rect 127374 6414 127426 6466
rect 127426 6414 127428 6466
rect 127372 6412 127428 6414
rect 128044 6412 128100 6468
rect 127148 6300 127204 6356
rect 126924 5068 126980 5124
rect 127372 4508 127428 4564
rect 127820 3724 127876 3780
rect 125692 3388 125748 3444
rect 126028 3388 126084 3444
rect 126364 3442 126420 3444
rect 126364 3390 126366 3442
rect 126366 3390 126418 3442
rect 126418 3390 126420 3442
rect 126364 3388 126420 3390
rect 127148 3442 127204 3444
rect 127148 3390 127150 3442
rect 127150 3390 127202 3442
rect 127202 3390 127204 3442
rect 127148 3388 127204 3390
rect 128940 8034 128996 8036
rect 128940 7982 128942 8034
rect 128942 7982 128994 8034
rect 128994 7982 128996 8034
rect 128940 7980 128996 7982
rect 128940 7250 128996 7252
rect 128940 7198 128942 7250
rect 128942 7198 128994 7250
rect 128994 7198 128996 7250
rect 128940 7196 128996 7198
rect 128492 5292 128548 5348
rect 128604 4844 128660 4900
rect 128604 4284 128660 4340
rect 130082 19626 130138 19628
rect 130082 19574 130084 19626
rect 130084 19574 130136 19626
rect 130136 19574 130138 19626
rect 130082 19572 130138 19574
rect 130186 19626 130242 19628
rect 130186 19574 130188 19626
rect 130188 19574 130240 19626
rect 130240 19574 130242 19626
rect 130186 19572 130242 19574
rect 130290 19626 130346 19628
rect 130290 19574 130292 19626
rect 130292 19574 130344 19626
rect 130344 19574 130346 19626
rect 130290 19572 130346 19574
rect 130082 18058 130138 18060
rect 130082 18006 130084 18058
rect 130084 18006 130136 18058
rect 130136 18006 130138 18058
rect 130082 18004 130138 18006
rect 130186 18058 130242 18060
rect 130186 18006 130188 18058
rect 130188 18006 130240 18058
rect 130240 18006 130242 18058
rect 130186 18004 130242 18006
rect 130290 18058 130346 18060
rect 130290 18006 130292 18058
rect 130292 18006 130344 18058
rect 130344 18006 130346 18058
rect 130290 18004 130346 18006
rect 130082 16490 130138 16492
rect 130082 16438 130084 16490
rect 130084 16438 130136 16490
rect 130136 16438 130138 16490
rect 130082 16436 130138 16438
rect 130186 16490 130242 16492
rect 130186 16438 130188 16490
rect 130188 16438 130240 16490
rect 130240 16438 130242 16490
rect 130186 16436 130242 16438
rect 130290 16490 130346 16492
rect 130290 16438 130292 16490
rect 130292 16438 130344 16490
rect 130344 16438 130346 16490
rect 130290 16436 130346 16438
rect 130082 14922 130138 14924
rect 130082 14870 130084 14922
rect 130084 14870 130136 14922
rect 130136 14870 130138 14922
rect 130082 14868 130138 14870
rect 130186 14922 130242 14924
rect 130186 14870 130188 14922
rect 130188 14870 130240 14922
rect 130240 14870 130242 14922
rect 130186 14868 130242 14870
rect 130290 14922 130346 14924
rect 130290 14870 130292 14922
rect 130292 14870 130344 14922
rect 130344 14870 130346 14922
rect 130290 14868 130346 14870
rect 130082 13354 130138 13356
rect 130082 13302 130084 13354
rect 130084 13302 130136 13354
rect 130136 13302 130138 13354
rect 130082 13300 130138 13302
rect 130186 13354 130242 13356
rect 130186 13302 130188 13354
rect 130188 13302 130240 13354
rect 130240 13302 130242 13354
rect 130186 13300 130242 13302
rect 130290 13354 130346 13356
rect 130290 13302 130292 13354
rect 130292 13302 130344 13354
rect 130344 13302 130346 13354
rect 130290 13300 130346 13302
rect 130082 11786 130138 11788
rect 130082 11734 130084 11786
rect 130084 11734 130136 11786
rect 130136 11734 130138 11786
rect 130082 11732 130138 11734
rect 130186 11786 130242 11788
rect 130186 11734 130188 11786
rect 130188 11734 130240 11786
rect 130240 11734 130242 11786
rect 130186 11732 130242 11734
rect 130290 11786 130346 11788
rect 130290 11734 130292 11786
rect 130292 11734 130344 11786
rect 130344 11734 130346 11786
rect 130290 11732 130346 11734
rect 130082 10218 130138 10220
rect 130082 10166 130084 10218
rect 130084 10166 130136 10218
rect 130136 10166 130138 10218
rect 130082 10164 130138 10166
rect 130186 10218 130242 10220
rect 130186 10166 130188 10218
rect 130188 10166 130240 10218
rect 130240 10166 130242 10218
rect 130186 10164 130242 10166
rect 130290 10218 130346 10220
rect 130290 10166 130292 10218
rect 130292 10166 130344 10218
rect 130344 10166 130346 10218
rect 130290 10164 130346 10166
rect 129500 9884 129556 9940
rect 129164 9042 129220 9044
rect 129164 8990 129166 9042
rect 129166 8990 129218 9042
rect 129218 8990 129220 9042
rect 129164 8988 129220 8990
rect 130172 9154 130228 9156
rect 130172 9102 130174 9154
rect 130174 9102 130226 9154
rect 130226 9102 130228 9154
rect 130172 9100 130228 9102
rect 131292 9154 131348 9156
rect 131292 9102 131294 9154
rect 131294 9102 131346 9154
rect 131346 9102 131348 9154
rect 131292 9100 131348 9102
rect 130082 8650 130138 8652
rect 130082 8598 130084 8650
rect 130084 8598 130136 8650
rect 130136 8598 130138 8650
rect 130082 8596 130138 8598
rect 130186 8650 130242 8652
rect 130186 8598 130188 8650
rect 130188 8598 130240 8650
rect 130240 8598 130242 8650
rect 130186 8596 130242 8598
rect 130290 8650 130346 8652
rect 130290 8598 130292 8650
rect 130292 8598 130344 8650
rect 130344 8598 130346 8650
rect 130290 8596 130346 8598
rect 129724 7586 129780 7588
rect 129724 7534 129726 7586
rect 129726 7534 129778 7586
rect 129778 7534 129780 7586
rect 129724 7532 129780 7534
rect 131292 7868 131348 7924
rect 130844 7420 130900 7476
rect 129164 6412 129220 6468
rect 129612 7308 129668 7364
rect 130082 7082 130138 7084
rect 130082 7030 130084 7082
rect 130084 7030 130136 7082
rect 130136 7030 130138 7082
rect 130082 7028 130138 7030
rect 130186 7082 130242 7084
rect 130186 7030 130188 7082
rect 130188 7030 130240 7082
rect 130240 7030 130242 7082
rect 130186 7028 130242 7030
rect 130290 7082 130346 7084
rect 130290 7030 130292 7082
rect 130292 7030 130344 7082
rect 130344 7030 130346 7082
rect 130290 7028 130346 7030
rect 130956 6524 131012 6580
rect 131516 6300 131572 6356
rect 131628 7644 131684 7700
rect 131628 6748 131684 6804
rect 130082 5514 130138 5516
rect 130082 5462 130084 5514
rect 130084 5462 130136 5514
rect 130136 5462 130138 5514
rect 130082 5460 130138 5462
rect 130186 5514 130242 5516
rect 130186 5462 130188 5514
rect 130188 5462 130240 5514
rect 130240 5462 130242 5514
rect 130186 5460 130242 5462
rect 130290 5514 130346 5516
rect 130290 5462 130292 5514
rect 130292 5462 130344 5514
rect 130344 5462 130346 5514
rect 130290 5460 130346 5462
rect 132300 8034 132356 8036
rect 132300 7982 132302 8034
rect 132302 7982 132354 8034
rect 132354 7982 132356 8034
rect 132300 7980 132356 7982
rect 132860 7868 132916 7924
rect 133644 7532 133700 7588
rect 132076 7084 132132 7140
rect 131964 6578 132020 6580
rect 131964 6526 131966 6578
rect 131966 6526 132018 6578
rect 132018 6526 132020 6578
rect 131964 6524 132020 6526
rect 131852 6412 131908 6468
rect 132076 6130 132132 6132
rect 132076 6078 132078 6130
rect 132078 6078 132130 6130
rect 132130 6078 132132 6130
rect 132076 6076 132132 6078
rect 133532 7362 133588 7364
rect 133532 7310 133534 7362
rect 133534 7310 133586 7362
rect 133586 7310 133588 7362
rect 133532 7308 133588 7310
rect 133084 7084 133140 7140
rect 132636 6412 132692 6468
rect 132188 5964 132244 6020
rect 131852 5628 131908 5684
rect 130956 5068 131012 5124
rect 132860 6188 132916 6244
rect 131964 5122 132020 5124
rect 131964 5070 131966 5122
rect 131966 5070 132018 5122
rect 132018 5070 132020 5122
rect 131964 5068 132020 5070
rect 132188 4508 132244 4564
rect 129612 4338 129668 4340
rect 129612 4286 129614 4338
rect 129614 4286 129666 4338
rect 129666 4286 129668 4338
rect 129612 4284 129668 4286
rect 132076 4172 132132 4228
rect 130082 3946 130138 3948
rect 130082 3894 130084 3946
rect 130084 3894 130136 3946
rect 130136 3894 130138 3946
rect 130082 3892 130138 3894
rect 130186 3946 130242 3948
rect 130186 3894 130188 3946
rect 130188 3894 130240 3946
rect 130240 3894 130242 3946
rect 130186 3892 130242 3894
rect 130290 3946 130346 3948
rect 130290 3894 130292 3946
rect 130292 3894 130344 3946
rect 130344 3894 130346 3946
rect 130290 3892 130346 3894
rect 131516 3778 131572 3780
rect 131516 3726 131518 3778
rect 131518 3726 131570 3778
rect 131570 3726 131572 3778
rect 131516 3724 131572 3726
rect 131628 3666 131684 3668
rect 131628 3614 131630 3666
rect 131630 3614 131682 3666
rect 131682 3614 131684 3666
rect 131628 3612 131684 3614
rect 129388 3500 129444 3556
rect 130284 3500 130340 3556
rect 132972 6076 133028 6132
rect 133084 6018 133140 6020
rect 133084 5966 133086 6018
rect 133086 5966 133138 6018
rect 133138 5966 133140 6018
rect 133084 5964 133140 5966
rect 132860 5404 132916 5460
rect 132636 4396 132692 4452
rect 133308 4956 133364 5012
rect 133196 4226 133252 4228
rect 133196 4174 133198 4226
rect 133198 4174 133250 4226
rect 133250 4174 133252 4226
rect 133196 4172 133252 4174
rect 132636 4114 132692 4116
rect 132636 4062 132638 4114
rect 132638 4062 132690 4114
rect 132690 4062 132692 4114
rect 132636 4060 132692 4062
rect 133308 3948 133364 4004
rect 132300 3778 132356 3780
rect 132300 3726 132302 3778
rect 132302 3726 132354 3778
rect 132354 3726 132356 3778
rect 132300 3724 132356 3726
rect 134204 6466 134260 6468
rect 134204 6414 134206 6466
rect 134206 6414 134258 6466
rect 134258 6414 134260 6466
rect 134204 6412 134260 6414
rect 134092 6018 134148 6020
rect 134092 5966 134094 6018
rect 134094 5966 134146 6018
rect 134146 5966 134148 6018
rect 134092 5964 134148 5966
rect 133980 5682 134036 5684
rect 133980 5630 133982 5682
rect 133982 5630 134034 5682
rect 134034 5630 134036 5682
rect 133980 5628 134036 5630
rect 134204 5068 134260 5124
rect 134316 5740 134372 5796
rect 133756 4508 133812 4564
rect 134316 4060 134372 4116
rect 133420 3724 133476 3780
rect 132188 3666 132244 3668
rect 132188 3614 132190 3666
rect 132190 3614 132242 3666
rect 132242 3614 132244 3666
rect 132188 3612 132244 3614
rect 134764 7980 134820 8036
rect 134540 4956 134596 5012
rect 137900 6018 137956 6020
rect 137900 5966 137902 6018
rect 137902 5966 137954 6018
rect 137954 5966 137956 6018
rect 137900 5964 137956 5966
rect 134988 5794 135044 5796
rect 134988 5742 134990 5794
rect 134990 5742 135042 5794
rect 135042 5742 135044 5794
rect 134988 5740 135044 5742
rect 137340 5628 137396 5684
rect 136220 5180 136276 5236
rect 135212 4956 135268 5012
rect 134876 4562 134932 4564
rect 134876 4510 134878 4562
rect 134878 4510 134930 4562
rect 134930 4510 134932 4562
rect 134876 4508 134932 4510
rect 136332 5122 136388 5124
rect 136332 5070 136334 5122
rect 136334 5070 136386 5122
rect 136386 5070 136388 5122
rect 136332 5068 136388 5070
rect 137004 4898 137060 4900
rect 137004 4846 137006 4898
rect 137006 4846 137058 4898
rect 137058 4846 137060 4898
rect 137004 4844 137060 4846
rect 137340 4396 137396 4452
rect 136892 4338 136948 4340
rect 136892 4286 136894 4338
rect 136894 4286 136946 4338
rect 136946 4286 136948 4338
rect 136892 4284 136948 4286
rect 137340 3612 137396 3668
rect 135660 3554 135716 3556
rect 135660 3502 135662 3554
rect 135662 3502 135714 3554
rect 135714 3502 135716 3554
rect 135660 3500 135716 3502
rect 137900 5292 137956 5348
rect 138684 6018 138740 6020
rect 138684 5966 138686 6018
rect 138686 5966 138738 6018
rect 138738 5966 138740 6018
rect 138684 5964 138740 5966
rect 138012 5234 138068 5236
rect 138012 5182 138014 5234
rect 138014 5182 138066 5234
rect 138066 5182 138068 5234
rect 138012 5180 138068 5182
rect 138348 5180 138404 5236
rect 133308 3442 133364 3444
rect 133308 3390 133310 3442
rect 133310 3390 133362 3442
rect 133362 3390 133364 3442
rect 133308 3388 133364 3390
rect 139244 33068 139300 33124
rect 139580 33458 139636 33460
rect 139580 33406 139582 33458
rect 139582 33406 139634 33458
rect 139634 33406 139636 33458
rect 139580 33404 139636 33406
rect 140700 35084 140756 35140
rect 141036 38220 141092 38276
rect 140924 36258 140980 36260
rect 140924 36206 140926 36258
rect 140926 36206 140978 36258
rect 140978 36206 140980 36258
rect 140924 36204 140980 36206
rect 141820 37212 141876 37268
rect 141820 36482 141876 36484
rect 141820 36430 141822 36482
rect 141822 36430 141874 36482
rect 141874 36430 141876 36482
rect 141820 36428 141876 36430
rect 142604 36540 142660 36596
rect 142156 36370 142212 36372
rect 142156 36318 142158 36370
rect 142158 36318 142210 36370
rect 142210 36318 142212 36370
rect 142156 36316 142212 36318
rect 143276 36428 143332 36484
rect 141036 35756 141092 35812
rect 140812 34972 140868 35028
rect 141148 35196 141204 35252
rect 141708 35026 141764 35028
rect 141708 34974 141710 35026
rect 141710 34974 141762 35026
rect 141762 34974 141764 35026
rect 141708 34972 141764 34974
rect 141820 34076 141876 34132
rect 141820 32396 141876 32452
rect 139356 6076 139412 6132
rect 138908 5404 138964 5460
rect 139916 6748 139972 6804
rect 139692 5682 139748 5684
rect 139692 5630 139694 5682
rect 139694 5630 139746 5682
rect 139746 5630 139748 5682
rect 139692 5628 139748 5630
rect 139692 5404 139748 5460
rect 139132 4956 139188 5012
rect 139020 4844 139076 4900
rect 139020 3666 139076 3668
rect 139020 3614 139022 3666
rect 139022 3614 139074 3666
rect 139074 3614 139076 3666
rect 139020 3612 139076 3614
rect 141260 6524 141316 6580
rect 140252 6130 140308 6132
rect 140252 6078 140254 6130
rect 140254 6078 140306 6130
rect 140306 6078 140308 6130
rect 140252 6076 140308 6078
rect 140812 5906 140868 5908
rect 140812 5854 140814 5906
rect 140814 5854 140866 5906
rect 140866 5854 140868 5906
rect 140812 5852 140868 5854
rect 140140 5234 140196 5236
rect 140140 5182 140142 5234
rect 140142 5182 140194 5234
rect 140194 5182 140196 5234
rect 140140 5180 140196 5182
rect 141372 5906 141428 5908
rect 141372 5854 141374 5906
rect 141374 5854 141426 5906
rect 141426 5854 141428 5906
rect 141372 5852 141428 5854
rect 141260 5740 141316 5796
rect 141372 5628 141428 5684
rect 142380 34188 142436 34244
rect 142828 35756 142884 35812
rect 143164 35810 143220 35812
rect 143164 35758 143166 35810
rect 143166 35758 143218 35810
rect 143218 35758 143220 35810
rect 143164 35756 143220 35758
rect 142940 35196 142996 35252
rect 143052 34242 143108 34244
rect 143052 34190 143054 34242
rect 143054 34190 143106 34242
rect 143106 34190 143108 34242
rect 143052 34188 143108 34190
rect 142940 34130 142996 34132
rect 142940 34078 142942 34130
rect 142942 34078 142994 34130
rect 142994 34078 142996 34130
rect 142940 34076 142996 34078
rect 143724 36988 143780 37044
rect 143500 34748 143556 34804
rect 143948 35196 144004 35252
rect 145292 36652 145348 36708
rect 146188 36652 146244 36708
rect 145740 36482 145796 36484
rect 145740 36430 145742 36482
rect 145742 36430 145794 36482
rect 145794 36430 145796 36482
rect 145740 36428 145796 36430
rect 144732 34802 144788 34804
rect 144732 34750 144734 34802
rect 144734 34750 144786 34802
rect 144786 34750 144788 34802
rect 144732 34748 144788 34750
rect 144396 33964 144452 34020
rect 144620 34636 144676 34692
rect 142380 28476 142436 28532
rect 142380 7308 142436 7364
rect 142492 7420 142548 7476
rect 142268 6860 142324 6916
rect 142492 6412 142548 6468
rect 142268 5852 142324 5908
rect 141932 5794 141988 5796
rect 141932 5742 141934 5794
rect 141934 5742 141986 5794
rect 141986 5742 141988 5794
rect 141932 5740 141988 5742
rect 143164 7196 143220 7252
rect 142716 6578 142772 6580
rect 142716 6526 142718 6578
rect 142718 6526 142770 6578
rect 142770 6526 142772 6578
rect 142716 6524 142772 6526
rect 142604 6076 142660 6132
rect 142492 5740 142548 5796
rect 141708 4844 141764 4900
rect 142716 4956 142772 5012
rect 142604 4844 142660 4900
rect 143164 4844 143220 4900
rect 141484 4396 141540 4452
rect 143836 7868 143892 7924
rect 143612 7084 143668 7140
rect 143500 6466 143556 6468
rect 143500 6414 143502 6466
rect 143502 6414 143554 6466
rect 143554 6414 143556 6466
rect 143500 6412 143556 6414
rect 143388 5964 143444 6020
rect 143500 4844 143556 4900
rect 143724 6130 143780 6132
rect 143724 6078 143726 6130
rect 143726 6078 143778 6130
rect 143778 6078 143780 6130
rect 143724 6076 143780 6078
rect 140140 3612 140196 3668
rect 138012 3442 138068 3444
rect 138012 3390 138014 3442
rect 138014 3390 138066 3442
rect 138066 3390 138068 3442
rect 138012 3388 138068 3390
rect 141036 3666 141092 3668
rect 141036 3614 141038 3666
rect 141038 3614 141090 3666
rect 141090 3614 141092 3666
rect 141036 3612 141092 3614
rect 143948 6860 144004 6916
rect 144508 5234 144564 5236
rect 144508 5182 144510 5234
rect 144510 5182 144562 5234
rect 144562 5182 144564 5234
rect 144508 5180 144564 5182
rect 144172 3612 144228 3668
rect 144060 3554 144116 3556
rect 144060 3502 144062 3554
rect 144062 3502 144114 3554
rect 144114 3502 144116 3554
rect 144060 3500 144116 3502
rect 147532 36594 147588 36596
rect 147532 36542 147534 36594
rect 147534 36542 147586 36594
rect 147586 36542 147588 36594
rect 147532 36540 147588 36542
rect 146860 36316 146916 36372
rect 148492 36090 148548 36092
rect 148492 36038 148494 36090
rect 148494 36038 148546 36090
rect 148546 36038 148548 36090
rect 148492 36036 148548 36038
rect 148596 36090 148652 36092
rect 148596 36038 148598 36090
rect 148598 36038 148650 36090
rect 148650 36038 148652 36090
rect 148596 36036 148652 36038
rect 148700 36090 148756 36092
rect 148700 36038 148702 36090
rect 148702 36038 148754 36090
rect 148754 36038 148756 36090
rect 148700 36036 148756 36038
rect 146188 35868 146244 35924
rect 146860 35922 146916 35924
rect 146860 35870 146862 35922
rect 146862 35870 146914 35922
rect 146914 35870 146916 35922
rect 146860 35868 146916 35870
rect 145292 34636 145348 34692
rect 145628 34690 145684 34692
rect 145628 34638 145630 34690
rect 145630 34638 145682 34690
rect 145682 34638 145684 34690
rect 145628 34636 145684 34638
rect 148492 34522 148548 34524
rect 148492 34470 148494 34522
rect 148494 34470 148546 34522
rect 148546 34470 148548 34522
rect 148492 34468 148548 34470
rect 148596 34522 148652 34524
rect 148596 34470 148598 34522
rect 148598 34470 148650 34522
rect 148650 34470 148652 34522
rect 148596 34468 148652 34470
rect 148700 34522 148756 34524
rect 148700 34470 148702 34522
rect 148702 34470 148754 34522
rect 148754 34470 148756 34522
rect 148700 34468 148756 34470
rect 145628 34018 145684 34020
rect 145628 33966 145630 34018
rect 145630 33966 145682 34018
rect 145682 33966 145684 34018
rect 145628 33964 145684 33966
rect 148492 32954 148548 32956
rect 148492 32902 148494 32954
rect 148494 32902 148546 32954
rect 148546 32902 148548 32954
rect 148492 32900 148548 32902
rect 148596 32954 148652 32956
rect 148596 32902 148598 32954
rect 148598 32902 148650 32954
rect 148650 32902 148652 32954
rect 148596 32900 148652 32902
rect 148700 32954 148756 32956
rect 148700 32902 148702 32954
rect 148702 32902 148754 32954
rect 148754 32902 148756 32954
rect 148700 32900 148756 32902
rect 147868 32732 147924 32788
rect 144844 31612 144900 31668
rect 145964 7756 146020 7812
rect 145292 6130 145348 6132
rect 145292 6078 145294 6130
rect 145294 6078 145346 6130
rect 145346 6078 145348 6130
rect 145292 6076 145348 6078
rect 144844 6018 144900 6020
rect 144844 5966 144846 6018
rect 144846 5966 144898 6018
rect 144898 5966 144900 6018
rect 144844 5964 144900 5966
rect 145068 4844 145124 4900
rect 145180 4956 145236 5012
rect 145180 4396 145236 4452
rect 145852 5234 145908 5236
rect 145852 5182 145854 5234
rect 145854 5182 145906 5234
rect 145906 5182 145908 5234
rect 145852 5180 145908 5182
rect 145964 4508 146020 4564
rect 145628 4450 145684 4452
rect 145628 4398 145630 4450
rect 145630 4398 145682 4450
rect 145682 4398 145684 4450
rect 145628 4396 145684 4398
rect 146524 6300 146580 6356
rect 145628 4172 145684 4228
rect 145068 3500 145124 3556
rect 148492 31386 148548 31388
rect 148492 31334 148494 31386
rect 148494 31334 148546 31386
rect 148546 31334 148548 31386
rect 148492 31332 148548 31334
rect 148596 31386 148652 31388
rect 148596 31334 148598 31386
rect 148598 31334 148650 31386
rect 148650 31334 148652 31386
rect 148596 31332 148652 31334
rect 148700 31386 148756 31388
rect 148700 31334 148702 31386
rect 148702 31334 148754 31386
rect 148754 31334 148756 31386
rect 148700 31332 148756 31334
rect 147980 31052 148036 31108
rect 148492 29818 148548 29820
rect 148492 29766 148494 29818
rect 148494 29766 148546 29818
rect 148546 29766 148548 29818
rect 148492 29764 148548 29766
rect 148596 29818 148652 29820
rect 148596 29766 148598 29818
rect 148598 29766 148650 29818
rect 148650 29766 148652 29818
rect 148596 29764 148652 29766
rect 148700 29818 148756 29820
rect 148700 29766 148702 29818
rect 148702 29766 148754 29818
rect 148754 29766 148756 29818
rect 148700 29764 148756 29766
rect 148492 28250 148548 28252
rect 148492 28198 148494 28250
rect 148494 28198 148546 28250
rect 148546 28198 148548 28250
rect 148492 28196 148548 28198
rect 148596 28250 148652 28252
rect 148596 28198 148598 28250
rect 148598 28198 148650 28250
rect 148650 28198 148652 28250
rect 148596 28196 148652 28198
rect 148700 28250 148756 28252
rect 148700 28198 148702 28250
rect 148702 28198 148754 28250
rect 148754 28198 148756 28250
rect 148700 28196 148756 28198
rect 148492 26682 148548 26684
rect 148492 26630 148494 26682
rect 148494 26630 148546 26682
rect 148546 26630 148548 26682
rect 148492 26628 148548 26630
rect 148596 26682 148652 26684
rect 148596 26630 148598 26682
rect 148598 26630 148650 26682
rect 148650 26630 148652 26682
rect 148596 26628 148652 26630
rect 148700 26682 148756 26684
rect 148700 26630 148702 26682
rect 148702 26630 148754 26682
rect 148754 26630 148756 26682
rect 148700 26628 148756 26630
rect 148492 25114 148548 25116
rect 148492 25062 148494 25114
rect 148494 25062 148546 25114
rect 148546 25062 148548 25114
rect 148492 25060 148548 25062
rect 148596 25114 148652 25116
rect 148596 25062 148598 25114
rect 148598 25062 148650 25114
rect 148650 25062 148652 25114
rect 148596 25060 148652 25062
rect 148700 25114 148756 25116
rect 148700 25062 148702 25114
rect 148702 25062 148754 25114
rect 148754 25062 148756 25114
rect 148700 25060 148756 25062
rect 148492 23546 148548 23548
rect 148492 23494 148494 23546
rect 148494 23494 148546 23546
rect 148546 23494 148548 23546
rect 148492 23492 148548 23494
rect 148596 23546 148652 23548
rect 148596 23494 148598 23546
rect 148598 23494 148650 23546
rect 148650 23494 148652 23546
rect 148596 23492 148652 23494
rect 148700 23546 148756 23548
rect 148700 23494 148702 23546
rect 148702 23494 148754 23546
rect 148754 23494 148756 23546
rect 148700 23492 148756 23494
rect 148492 21978 148548 21980
rect 148492 21926 148494 21978
rect 148494 21926 148546 21978
rect 148546 21926 148548 21978
rect 148492 21924 148548 21926
rect 148596 21978 148652 21980
rect 148596 21926 148598 21978
rect 148598 21926 148650 21978
rect 148650 21926 148652 21978
rect 148596 21924 148652 21926
rect 148700 21978 148756 21980
rect 148700 21926 148702 21978
rect 148702 21926 148754 21978
rect 148754 21926 148756 21978
rect 148700 21924 148756 21926
rect 148492 20410 148548 20412
rect 148492 20358 148494 20410
rect 148494 20358 148546 20410
rect 148546 20358 148548 20410
rect 148492 20356 148548 20358
rect 148596 20410 148652 20412
rect 148596 20358 148598 20410
rect 148598 20358 148650 20410
rect 148650 20358 148652 20410
rect 148596 20356 148652 20358
rect 148700 20410 148756 20412
rect 148700 20358 148702 20410
rect 148702 20358 148754 20410
rect 148754 20358 148756 20410
rect 148700 20356 148756 20358
rect 148492 18842 148548 18844
rect 148492 18790 148494 18842
rect 148494 18790 148546 18842
rect 148546 18790 148548 18842
rect 148492 18788 148548 18790
rect 148596 18842 148652 18844
rect 148596 18790 148598 18842
rect 148598 18790 148650 18842
rect 148650 18790 148652 18842
rect 148596 18788 148652 18790
rect 148700 18842 148756 18844
rect 148700 18790 148702 18842
rect 148702 18790 148754 18842
rect 148754 18790 148756 18842
rect 148700 18788 148756 18790
rect 148492 17274 148548 17276
rect 148492 17222 148494 17274
rect 148494 17222 148546 17274
rect 148546 17222 148548 17274
rect 148492 17220 148548 17222
rect 148596 17274 148652 17276
rect 148596 17222 148598 17274
rect 148598 17222 148650 17274
rect 148650 17222 148652 17274
rect 148596 17220 148652 17222
rect 148700 17274 148756 17276
rect 148700 17222 148702 17274
rect 148702 17222 148754 17274
rect 148754 17222 148756 17274
rect 148700 17220 148756 17222
rect 148492 15706 148548 15708
rect 148492 15654 148494 15706
rect 148494 15654 148546 15706
rect 148546 15654 148548 15706
rect 148492 15652 148548 15654
rect 148596 15706 148652 15708
rect 148596 15654 148598 15706
rect 148598 15654 148650 15706
rect 148650 15654 148652 15706
rect 148596 15652 148652 15654
rect 148700 15706 148756 15708
rect 148700 15654 148702 15706
rect 148702 15654 148754 15706
rect 148754 15654 148756 15706
rect 148700 15652 148756 15654
rect 148492 14138 148548 14140
rect 148492 14086 148494 14138
rect 148494 14086 148546 14138
rect 148546 14086 148548 14138
rect 148492 14084 148548 14086
rect 148596 14138 148652 14140
rect 148596 14086 148598 14138
rect 148598 14086 148650 14138
rect 148650 14086 148652 14138
rect 148596 14084 148652 14086
rect 148700 14138 148756 14140
rect 148700 14086 148702 14138
rect 148702 14086 148754 14138
rect 148754 14086 148756 14138
rect 148700 14084 148756 14086
rect 148492 12570 148548 12572
rect 148492 12518 148494 12570
rect 148494 12518 148546 12570
rect 148546 12518 148548 12570
rect 148492 12516 148548 12518
rect 148596 12570 148652 12572
rect 148596 12518 148598 12570
rect 148598 12518 148650 12570
rect 148650 12518 148652 12570
rect 148596 12516 148652 12518
rect 148700 12570 148756 12572
rect 148700 12518 148702 12570
rect 148702 12518 148754 12570
rect 148754 12518 148756 12570
rect 148700 12516 148756 12518
rect 148492 11002 148548 11004
rect 148492 10950 148494 11002
rect 148494 10950 148546 11002
rect 148546 10950 148548 11002
rect 148492 10948 148548 10950
rect 148596 11002 148652 11004
rect 148596 10950 148598 11002
rect 148598 10950 148650 11002
rect 148650 10950 148652 11002
rect 148596 10948 148652 10950
rect 148700 11002 148756 11004
rect 148700 10950 148702 11002
rect 148702 10950 148754 11002
rect 148754 10950 148756 11002
rect 148700 10948 148756 10950
rect 148492 9434 148548 9436
rect 148492 9382 148494 9434
rect 148494 9382 148546 9434
rect 148546 9382 148548 9434
rect 148492 9380 148548 9382
rect 148596 9434 148652 9436
rect 148596 9382 148598 9434
rect 148598 9382 148650 9434
rect 148650 9382 148652 9434
rect 148596 9380 148652 9382
rect 148700 9434 148756 9436
rect 148700 9382 148702 9434
rect 148702 9382 148754 9434
rect 148754 9382 148756 9434
rect 148700 9380 148756 9382
rect 148492 7866 148548 7868
rect 148492 7814 148494 7866
rect 148494 7814 148546 7866
rect 148546 7814 148548 7866
rect 148492 7812 148548 7814
rect 148596 7866 148652 7868
rect 148596 7814 148598 7866
rect 148598 7814 148650 7866
rect 148650 7814 148652 7866
rect 148596 7812 148652 7814
rect 148700 7866 148756 7868
rect 148700 7814 148702 7866
rect 148702 7814 148754 7866
rect 148754 7814 148756 7866
rect 148700 7812 148756 7814
rect 148492 6298 148548 6300
rect 148492 6246 148494 6298
rect 148494 6246 148546 6298
rect 148546 6246 148548 6298
rect 148492 6244 148548 6246
rect 148596 6298 148652 6300
rect 148596 6246 148598 6298
rect 148598 6246 148650 6298
rect 148650 6246 148652 6298
rect 148596 6244 148652 6246
rect 148700 6298 148756 6300
rect 148700 6246 148702 6298
rect 148702 6246 148754 6298
rect 148754 6246 148756 6298
rect 148700 6244 148756 6246
rect 147980 6076 148036 6132
rect 147868 5180 147924 5236
rect 148492 4730 148548 4732
rect 148492 4678 148494 4730
rect 148494 4678 148546 4730
rect 148546 4678 148548 4730
rect 148492 4676 148548 4678
rect 148596 4730 148652 4732
rect 148596 4678 148598 4730
rect 148598 4678 148650 4730
rect 148650 4678 148652 4730
rect 148596 4676 148652 4678
rect 148700 4730 148756 4732
rect 148700 4678 148702 4730
rect 148702 4678 148754 4730
rect 148754 4678 148756 4730
rect 148700 4676 148756 4678
rect 146748 4562 146804 4564
rect 146748 4510 146750 4562
rect 146750 4510 146802 4562
rect 146802 4510 146804 4562
rect 146748 4508 146804 4510
rect 147196 4226 147252 4228
rect 147196 4174 147198 4226
rect 147198 4174 147250 4226
rect 147250 4174 147252 4226
rect 147196 4172 147252 4174
rect 147532 3666 147588 3668
rect 147532 3614 147534 3666
rect 147534 3614 147586 3666
rect 147586 3614 147588 3666
rect 147532 3612 147588 3614
rect 148492 3162 148548 3164
rect 148492 3110 148494 3162
rect 148494 3110 148546 3162
rect 148546 3110 148548 3162
rect 148492 3108 148548 3110
rect 148596 3162 148652 3164
rect 148596 3110 148598 3162
rect 148598 3110 148650 3162
rect 148650 3110 148652 3162
rect 148596 3108 148652 3110
rect 148700 3162 148756 3164
rect 148700 3110 148702 3162
rect 148702 3110 148754 3162
rect 148754 3110 148756 3162
rect 148700 3108 148756 3110
<< metal3 >>
rect 22754 38892 22764 38948
rect 22820 38892 82796 38948
rect 82852 38892 82862 38948
rect 30034 38780 30044 38836
rect 30100 38780 85820 38836
rect 85876 38780 85886 38836
rect 43922 38668 43932 38724
rect 43988 38668 75292 38724
rect 75348 38668 75358 38724
rect 78754 38668 78764 38724
rect 78820 38668 113260 38724
rect 113316 38668 113326 38724
rect 71138 38556 71148 38612
rect 71204 38556 125356 38612
rect 125412 38556 125422 38612
rect 69906 38444 69916 38500
rect 69972 38444 109676 38500
rect 109732 38444 109742 38500
rect 67218 38332 67228 38388
rect 67284 38332 117628 38388
rect 117684 38332 117694 38388
rect 70802 38220 70812 38276
rect 70868 38220 141036 38276
rect 141092 38220 141102 38276
rect 56242 38108 56252 38164
rect 56308 38108 84028 38164
rect 84084 38108 84094 38164
rect 43026 37996 43036 38052
rect 43092 37996 76412 38052
rect 76468 37996 76478 38052
rect 77298 37996 77308 38052
rect 77364 37996 78652 38052
rect 78708 37996 111580 38052
rect 111636 37996 111646 38052
rect 36306 37884 36316 37940
rect 36372 37884 65660 37940
rect 65716 37884 65726 37940
rect 69794 37884 69804 37940
rect 69860 37884 107884 37940
rect 107940 37884 107950 37940
rect 63634 37772 63644 37828
rect 63700 37772 104748 37828
rect 104804 37772 104814 37828
rect 62514 37660 62524 37716
rect 62580 37660 105756 37716
rect 105812 37660 105822 37716
rect 38994 37548 39004 37604
rect 39060 37548 68012 37604
rect 68068 37548 68078 37604
rect 69010 37548 69020 37604
rect 69076 37548 113148 37604
rect 113204 37548 113214 37604
rect 64082 37436 64092 37492
rect 64148 37436 65436 37492
rect 65492 37436 117180 37492
rect 117236 37436 117246 37492
rect 73490 37324 73500 37380
rect 73556 37324 73724 37380
rect 73780 37324 94332 37380
rect 94388 37324 94398 37380
rect 44594 37212 44604 37268
rect 44660 37212 73164 37268
rect 73220 37212 73230 37268
rect 81554 37212 81564 37268
rect 81620 37212 100156 37268
rect 100212 37212 100222 37268
rect 105634 37212 105644 37268
rect 105700 37212 141820 37268
rect 141876 37212 141886 37268
rect 82562 37100 82572 37156
rect 82628 37100 106988 37156
rect 107044 37100 107054 37156
rect 117618 37100 117628 37156
rect 117684 37100 119196 37156
rect 119252 37100 121548 37156
rect 121604 37100 121614 37156
rect 16594 36988 16604 37044
rect 16660 36988 45276 37044
rect 45332 36988 45342 37044
rect 75618 36988 75628 37044
rect 75684 36988 91420 37044
rect 91476 36988 92764 37044
rect 92820 36988 92830 37044
rect 93314 36988 93324 37044
rect 93380 36988 94612 37044
rect 110562 36988 110572 37044
rect 110628 36988 143724 37044
rect 143780 36988 143790 37044
rect 94556 36932 94612 36988
rect 8418 36876 8428 36932
rect 8484 36876 9100 36932
rect 9156 36876 9166 36932
rect 66546 36876 66556 36932
rect 66612 36876 85708 36932
rect 94546 36876 94556 36932
rect 94612 36876 94622 36932
rect 19612 36820 19622 36876
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19886 36820 19896 36876
rect 56432 36820 56442 36876
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56706 36820 56716 36876
rect 77186 36764 77196 36820
rect 77252 36764 78988 36820
rect 79044 36764 79054 36820
rect 85652 36708 85708 36876
rect 93252 36820 93262 36876
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93526 36820 93536 36876
rect 130072 36820 130082 36876
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130346 36820 130356 36876
rect 93650 36764 93660 36820
rect 93716 36764 102508 36820
rect 132738 36764 132748 36820
rect 132804 36764 133868 36820
rect 133924 36764 133934 36820
rect 24210 36652 24220 36708
rect 24276 36652 35756 36708
rect 35812 36652 35822 36708
rect 49522 36652 49532 36708
rect 49588 36652 78988 36708
rect 85652 36652 96236 36708
rect 96292 36652 96302 36708
rect 78932 36596 78988 36652
rect 102452 36596 102508 36764
rect 118402 36652 118412 36708
rect 118468 36652 120428 36708
rect 120484 36652 122220 36708
rect 122276 36652 122286 36708
rect 145282 36652 145292 36708
rect 145348 36652 146188 36708
rect 146244 36652 146254 36708
rect 13906 36540 13916 36596
rect 13972 36540 15372 36596
rect 15428 36540 15438 36596
rect 27682 36540 27692 36596
rect 27748 36540 30940 36596
rect 30996 36540 31006 36596
rect 32274 36540 32284 36596
rect 32340 36540 47404 36596
rect 47460 36540 47470 36596
rect 48066 36540 48076 36596
rect 48132 36540 55468 36596
rect 68450 36540 68460 36596
rect 68516 36540 69132 36596
rect 69188 36540 69198 36596
rect 71698 36540 71708 36596
rect 71764 36540 74508 36596
rect 74564 36540 74574 36596
rect 78932 36540 101612 36596
rect 101668 36540 101678 36596
rect 102452 36540 119420 36596
rect 119476 36540 119486 36596
rect 120642 36540 120652 36596
rect 120708 36540 123340 36596
rect 123396 36540 123406 36596
rect 142594 36540 142604 36596
rect 142660 36540 147532 36596
rect 147588 36540 147598 36596
rect 55412 36484 55468 36540
rect 20626 36428 20636 36484
rect 20692 36428 26740 36484
rect 26898 36428 26908 36484
rect 26964 36428 31948 36484
rect 33506 36428 33516 36484
rect 33572 36428 35084 36484
rect 35140 36428 35150 36484
rect 37426 36428 37436 36484
rect 37492 36428 38892 36484
rect 38948 36428 38958 36484
rect 40338 36428 40348 36484
rect 40404 36428 47908 36484
rect 49186 36428 49196 36484
rect 49252 36428 50988 36484
rect 51044 36428 51054 36484
rect 53106 36428 53116 36484
rect 53172 36428 54796 36484
rect 54852 36428 54862 36484
rect 55412 36428 85708 36484
rect 86146 36428 86156 36484
rect 86212 36428 86828 36484
rect 86884 36428 89068 36484
rect 89124 36428 89134 36484
rect 98690 36428 98700 36484
rect 98756 36428 100828 36484
rect 100884 36428 103628 36484
rect 103684 36428 103694 36484
rect 105746 36428 105756 36484
rect 105812 36428 109900 36484
rect 109956 36428 109966 36484
rect 128930 36428 128940 36484
rect 128996 36428 129836 36484
rect 129892 36428 129902 36484
rect 130620 36428 135100 36484
rect 135156 36428 135166 36484
rect 141810 36428 141820 36484
rect 141876 36428 143276 36484
rect 143332 36428 145740 36484
rect 145796 36428 145806 36484
rect 26684 36372 26740 36428
rect 31892 36372 31948 36428
rect 47852 36372 47908 36428
rect 85652 36372 85708 36428
rect 11778 36316 11788 36372
rect 11844 36316 12908 36372
rect 12964 36316 12974 36372
rect 21410 36316 21420 36372
rect 21476 36316 22204 36372
rect 22260 36316 22270 36372
rect 22530 36316 22540 36372
rect 22596 36316 22876 36372
rect 22932 36316 22942 36372
rect 26684 36316 29260 36372
rect 29316 36316 30604 36372
rect 30660 36316 30670 36372
rect 31892 36316 36652 36372
rect 36708 36316 36718 36372
rect 45266 36316 45276 36372
rect 45332 36316 46116 36372
rect 46834 36316 46844 36372
rect 46900 36316 47628 36372
rect 47684 36316 47694 36372
rect 47852 36316 52892 36372
rect 52948 36316 52958 36372
rect 60834 36316 60844 36372
rect 60900 36316 65548 36372
rect 65604 36316 65884 36372
rect 65940 36316 65950 36372
rect 68898 36316 68908 36372
rect 68964 36316 72380 36372
rect 72436 36316 75628 36372
rect 75684 36316 75694 36372
rect 79090 36316 79100 36372
rect 79156 36316 81228 36372
rect 81284 36316 83020 36372
rect 83076 36316 83086 36372
rect 85652 36316 89180 36372
rect 89236 36316 89516 36372
rect 89572 36316 89582 36372
rect 89842 36316 89852 36372
rect 89908 36316 90748 36372
rect 90804 36316 90814 36372
rect 96002 36316 96012 36372
rect 96068 36316 97468 36372
rect 97524 36316 99036 36372
rect 99092 36316 99102 36372
rect 104066 36316 104076 36372
rect 104132 36316 105308 36372
rect 105364 36316 105374 36372
rect 107650 36316 107660 36372
rect 107716 36316 108892 36372
rect 108948 36316 108958 36372
rect 111234 36316 111244 36372
rect 111300 36316 112588 36372
rect 112644 36316 114380 36372
rect 114436 36316 114446 36372
rect 114818 36316 114828 36372
rect 114884 36316 116508 36372
rect 116564 36316 118300 36372
rect 118356 36316 118366 36372
rect 121986 36316 121996 36372
rect 122052 36316 124348 36372
rect 124404 36316 126140 36372
rect 126196 36316 126206 36372
rect 127698 36316 127708 36372
rect 127764 36316 130396 36372
rect 130452 36316 130462 36372
rect 46060 36260 46116 36316
rect 6066 36204 6076 36260
rect 6132 36204 6636 36260
rect 6692 36204 6702 36260
rect 9986 36204 9996 36260
rect 10052 36204 10780 36260
rect 10836 36204 10846 36260
rect 18610 36204 18620 36260
rect 18676 36204 20188 36260
rect 20244 36204 20254 36260
rect 27570 36204 27580 36260
rect 27636 36204 33964 36260
rect 34020 36204 34030 36260
rect 37772 36204 38500 36260
rect 41122 36204 41132 36260
rect 41188 36204 45836 36260
rect 45892 36204 45902 36260
rect 46060 36204 49644 36260
rect 49700 36204 49710 36260
rect 49970 36204 49980 36260
rect 50036 36204 51548 36260
rect 51604 36204 51614 36260
rect 69682 36204 69692 36260
rect 69748 36204 72492 36260
rect 72548 36204 72558 36260
rect 82226 36204 82236 36260
rect 82292 36204 84924 36260
rect 84980 36204 84990 36260
rect 90178 36204 90188 36260
rect 90244 36204 93660 36260
rect 93716 36204 93726 36260
rect 104850 36204 104860 36260
rect 104916 36204 106316 36260
rect 106372 36204 110684 36260
rect 110740 36204 110750 36260
rect 120082 36204 120092 36260
rect 120148 36204 121436 36260
rect 121492 36204 121502 36260
rect 125682 36204 125692 36260
rect 125748 36204 127932 36260
rect 127988 36204 127998 36260
rect 37772 36148 37828 36204
rect 29586 36092 29596 36148
rect 29652 36092 37828 36148
rect 38444 36148 38500 36204
rect 130620 36148 130676 36428
rect 134530 36316 134540 36372
rect 134596 36316 135324 36372
rect 135380 36316 136108 36372
rect 136164 36316 136174 36372
rect 138114 36316 138124 36372
rect 138180 36316 140028 36372
rect 140084 36316 140094 36372
rect 142146 36316 142156 36372
rect 142212 36316 146860 36372
rect 146916 36316 146926 36372
rect 131618 36204 131628 36260
rect 131684 36204 133980 36260
rect 134036 36204 134046 36260
rect 137106 36204 137116 36260
rect 137172 36204 138012 36260
rect 138068 36204 140924 36260
rect 140980 36204 140990 36260
rect 38444 36092 44716 36148
rect 44772 36092 44782 36148
rect 46274 36092 46284 36148
rect 46340 36092 59500 36148
rect 59556 36092 59566 36148
rect 84466 36092 84476 36148
rect 84532 36092 96460 36148
rect 96516 36092 96526 36148
rect 115042 36092 115052 36148
rect 115108 36092 130676 36148
rect 132692 36092 139020 36148
rect 139076 36092 139086 36148
rect 38022 36036 38032 36092
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38296 36036 38306 36092
rect 74842 36036 74852 36092
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 75116 36036 75126 36092
rect 111662 36036 111672 36092
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111936 36036 111946 36092
rect 132692 36036 132748 36092
rect 148482 36036 148492 36092
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148756 36036 148766 36092
rect 18274 35980 18284 36036
rect 18340 35980 21868 36036
rect 21924 35980 21934 36036
rect 39106 35980 39116 36036
rect 39172 35980 45724 36036
rect 45780 35980 45790 36036
rect 51090 35980 51100 36036
rect 51156 35980 73108 36036
rect 73052 35924 73108 35980
rect 78932 35980 91420 36036
rect 91476 35980 91486 36036
rect 91756 35980 100380 36036
rect 100436 35980 101500 36036
rect 101556 35980 102172 36036
rect 102228 35980 105084 36036
rect 105140 35980 105150 36036
rect 115378 35980 115388 36036
rect 115444 35980 132748 36036
rect 133522 35980 133532 36036
rect 133588 35980 137116 36036
rect 137172 35980 137182 36036
rect 78932 35924 78988 35980
rect 91756 35924 91812 35980
rect 7858 35868 7868 35924
rect 7924 35868 9660 35924
rect 9716 35868 9726 35924
rect 21410 35868 21420 35924
rect 21476 35868 22540 35924
rect 22596 35868 22606 35924
rect 27010 35868 27020 35924
rect 27076 35868 48412 35924
rect 48468 35868 48478 35924
rect 52770 35868 52780 35924
rect 52836 35868 69692 35924
rect 69748 35868 69758 35924
rect 73052 35868 78988 35924
rect 82226 35868 82236 35924
rect 82292 35868 91812 35924
rect 92418 35868 92428 35924
rect 92484 35868 92988 35924
rect 93044 35868 93054 35924
rect 94322 35868 94332 35924
rect 94388 35868 111356 35924
rect 111412 35868 111692 35924
rect 111748 35868 111758 35924
rect 113922 35868 113932 35924
rect 113988 35868 125804 35924
rect 125860 35868 125870 35924
rect 129490 35868 129500 35924
rect 129556 35868 132188 35924
rect 132244 35868 132254 35924
rect 146178 35868 146188 35924
rect 146244 35868 146860 35924
rect 146916 35868 146926 35924
rect 12786 35756 12796 35812
rect 12852 35756 19740 35812
rect 19796 35756 19806 35812
rect 35746 35756 35756 35812
rect 35812 35756 39340 35812
rect 39396 35756 39406 35812
rect 52210 35756 52220 35812
rect 52276 35756 52668 35812
rect 52724 35756 52734 35812
rect 56802 35756 56812 35812
rect 56868 35756 57596 35812
rect 57652 35756 57662 35812
rect 74722 35756 74732 35812
rect 74788 35756 75292 35812
rect 75348 35756 75628 35812
rect 75684 35756 75694 35812
rect 76290 35756 76300 35812
rect 76356 35756 78092 35812
rect 78148 35756 78158 35812
rect 83458 35756 83468 35812
rect 83524 35756 84924 35812
rect 84980 35756 84990 35812
rect 85250 35756 85260 35812
rect 85316 35756 86716 35812
rect 86772 35756 86782 35812
rect 91522 35756 91532 35812
rect 91588 35756 98252 35812
rect 98308 35756 98700 35812
rect 98756 35756 98766 35812
rect 105858 35756 105868 35812
rect 105924 35756 107100 35812
rect 107156 35756 108892 35812
rect 108948 35756 108958 35812
rect 109442 35756 109452 35812
rect 109508 35756 110124 35812
rect 110180 35756 110908 35812
rect 110964 35756 110974 35812
rect 113026 35756 113036 35812
rect 113092 35756 114268 35812
rect 114324 35756 116060 35812
rect 116116 35756 116126 35812
rect 122546 35756 122556 35812
rect 122612 35756 123116 35812
rect 123172 35756 123182 35812
rect 129042 35756 129052 35812
rect 129108 35756 130732 35812
rect 130788 35756 130798 35812
rect 133634 35756 133644 35812
rect 133700 35756 135660 35812
rect 135716 35756 135726 35812
rect 141026 35756 141036 35812
rect 141092 35756 142828 35812
rect 142884 35756 143164 35812
rect 143220 35756 143230 35812
rect 20402 35644 20412 35700
rect 20468 35644 22764 35700
rect 22820 35644 22830 35700
rect 48738 35644 48748 35700
rect 48804 35644 54572 35700
rect 54628 35644 54638 35700
rect 72706 35644 72716 35700
rect 72772 35644 77308 35700
rect 77364 35644 77374 35700
rect 89954 35644 89964 35700
rect 90020 35644 90412 35700
rect 90468 35644 91196 35700
rect 91252 35644 93772 35700
rect 93828 35644 95564 35700
rect 95620 35644 98588 35700
rect 98644 35644 100940 35700
rect 100996 35644 101006 35700
rect 103730 35644 103740 35700
rect 103796 35644 105532 35700
rect 105588 35644 105598 35700
rect 115602 35644 115612 35700
rect 115668 35644 115948 35700
rect 116004 35644 116014 35700
rect 125570 35644 125580 35700
rect 125636 35644 131628 35700
rect 131684 35644 131694 35700
rect 132626 35644 132636 35700
rect 132692 35644 134988 35700
rect 135044 35644 135054 35700
rect 23090 35532 23100 35588
rect 23156 35532 23884 35588
rect 23940 35532 32508 35588
rect 32564 35532 32574 35588
rect 50418 35532 50428 35588
rect 50484 35532 62636 35588
rect 62692 35532 62702 35588
rect 63074 35532 63084 35588
rect 63140 35532 68908 35588
rect 68964 35532 68974 35588
rect 74834 35532 74844 35588
rect 74900 35532 77084 35588
rect 77140 35532 77150 35588
rect 78418 35532 78428 35588
rect 78484 35532 79772 35588
rect 79828 35532 79838 35588
rect 92082 35532 92092 35588
rect 92148 35532 94780 35588
rect 94836 35532 94846 35588
rect 102060 35532 121100 35588
rect 121156 35532 121166 35588
rect 123442 35532 123452 35588
rect 123508 35532 124796 35588
rect 124852 35532 124862 35588
rect 126812 35532 137004 35588
rect 137060 35532 137070 35588
rect 62636 35476 62692 35532
rect 102060 35476 102116 35532
rect 126812 35476 126868 35532
rect 19058 35420 19068 35476
rect 19124 35420 19628 35476
rect 19684 35420 19694 35476
rect 40002 35420 40012 35476
rect 40068 35420 42028 35476
rect 42084 35420 42094 35476
rect 50194 35420 50204 35476
rect 50260 35420 51660 35476
rect 51716 35420 51726 35476
rect 51996 35420 62412 35476
rect 62468 35420 62478 35476
rect 62636 35420 64876 35476
rect 64932 35420 65548 35476
rect 65604 35420 65614 35476
rect 66322 35420 66332 35476
rect 66388 35420 67004 35476
rect 67060 35420 67228 35476
rect 76290 35420 76300 35476
rect 76356 35420 78764 35476
rect 78820 35420 78830 35476
rect 78932 35420 97468 35476
rect 99362 35420 99372 35476
rect 99428 35420 102060 35476
rect 102116 35420 102126 35476
rect 102386 35420 102396 35476
rect 102452 35420 102620 35476
rect 102676 35420 102686 35476
rect 104066 35420 104076 35476
rect 104132 35420 110908 35476
rect 110964 35420 110974 35476
rect 119858 35420 119868 35476
rect 119924 35420 120540 35476
rect 120596 35420 126868 35476
rect 127922 35420 127932 35476
rect 127988 35420 129164 35476
rect 129220 35420 134764 35476
rect 134820 35420 134830 35476
rect 51996 35364 52052 35420
rect 13346 35308 13356 35364
rect 13412 35308 14252 35364
rect 14308 35308 14318 35364
rect 24882 35308 24892 35364
rect 24948 35308 25564 35364
rect 25620 35308 41580 35364
rect 41636 35308 41646 35364
rect 46386 35308 46396 35364
rect 46452 35308 52052 35364
rect 65548 35364 65604 35420
rect 67172 35364 67228 35420
rect 78932 35364 78988 35420
rect 97412 35364 97468 35420
rect 65548 35308 66220 35364
rect 66276 35308 66286 35364
rect 67172 35308 78988 35364
rect 96450 35308 96460 35364
rect 96516 35308 97244 35364
rect 97300 35308 97310 35364
rect 97412 35308 106092 35364
rect 106148 35308 106158 35364
rect 108434 35308 108444 35364
rect 108500 35308 123004 35364
rect 123060 35308 123070 35364
rect 136322 35308 136332 35364
rect 136388 35308 136780 35364
rect 136836 35308 138012 35364
rect 138068 35308 138078 35364
rect 19612 35252 19622 35308
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19886 35252 19896 35308
rect 56432 35252 56442 35308
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56706 35252 56716 35308
rect 93252 35252 93262 35308
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93526 35252 93536 35308
rect 130072 35252 130082 35308
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130346 35252 130356 35308
rect 20132 35196 27804 35252
rect 27860 35196 28364 35252
rect 28420 35196 28430 35252
rect 57026 35196 57036 35252
rect 57092 35196 62300 35252
rect 62356 35196 62366 35252
rect 78932 35196 88956 35252
rect 89012 35196 90300 35252
rect 90356 35196 90366 35252
rect 90738 35196 90748 35252
rect 90804 35196 92764 35252
rect 92820 35196 92830 35252
rect 95106 35196 95116 35252
rect 95172 35196 97580 35252
rect 97636 35196 97646 35252
rect 101378 35196 101388 35252
rect 101444 35196 101612 35252
rect 101668 35196 102396 35252
rect 102452 35196 102462 35252
rect 102722 35196 102732 35252
rect 102788 35196 111860 35252
rect 112018 35196 112028 35252
rect 112084 35196 114828 35252
rect 114884 35196 114894 35252
rect 117282 35196 117292 35252
rect 117348 35196 118412 35252
rect 118468 35196 118478 35252
rect 120306 35196 120316 35252
rect 120372 35196 121100 35252
rect 121156 35196 122108 35252
rect 122164 35196 122174 35252
rect 132738 35196 132748 35252
rect 132804 35196 138796 35252
rect 138852 35196 138862 35252
rect 139346 35196 139356 35252
rect 139412 35196 141148 35252
rect 141204 35196 141214 35252
rect 142930 35196 142940 35252
rect 142996 35196 143948 35252
rect 144004 35196 144014 35252
rect 20132 35140 20188 35196
rect 78932 35140 78988 35196
rect 90300 35140 90356 35196
rect 111804 35140 111860 35196
rect 7298 35084 7308 35140
rect 7364 35084 8428 35140
rect 8484 35084 8494 35140
rect 18610 35084 18620 35140
rect 18676 35084 20188 35140
rect 20626 35084 20636 35140
rect 20692 35084 21868 35140
rect 21924 35084 21934 35140
rect 28130 35084 28140 35140
rect 28196 35084 28812 35140
rect 28868 35084 28878 35140
rect 42802 35084 42812 35140
rect 42868 35084 43148 35140
rect 43204 35084 53564 35140
rect 53620 35084 53630 35140
rect 68114 35084 68124 35140
rect 68180 35084 69356 35140
rect 69412 35084 69916 35140
rect 69972 35084 69982 35140
rect 75618 35084 75628 35140
rect 75684 35084 78988 35140
rect 80882 35084 80892 35140
rect 80948 35084 82572 35140
rect 82628 35084 82638 35140
rect 84354 35084 84364 35140
rect 84420 35084 85932 35140
rect 85988 35084 85998 35140
rect 87042 35084 87052 35140
rect 87108 35084 87948 35140
rect 88004 35084 88014 35140
rect 90300 35084 91308 35140
rect 91364 35084 91374 35140
rect 91522 35084 91532 35140
rect 91588 35084 93324 35140
rect 93380 35084 93390 35140
rect 94210 35084 94220 35140
rect 94276 35084 95788 35140
rect 95844 35084 95854 35140
rect 97794 35084 97804 35140
rect 97860 35084 99260 35140
rect 99316 35084 99326 35140
rect 100482 35084 100492 35140
rect 100548 35084 101836 35140
rect 101892 35084 101902 35140
rect 106866 35084 106876 35140
rect 106932 35084 107436 35140
rect 107492 35084 107502 35140
rect 108546 35084 108556 35140
rect 108612 35084 109788 35140
rect 109844 35084 109854 35140
rect 110338 35084 110348 35140
rect 110404 35084 111580 35140
rect 111636 35084 111646 35140
rect 111804 35084 113428 35140
rect 114034 35084 114044 35140
rect 114100 35084 115500 35140
rect 115556 35084 115566 35140
rect 116610 35084 116620 35140
rect 116676 35084 117068 35140
rect 117124 35084 117852 35140
rect 117908 35084 117918 35140
rect 119410 35084 119420 35140
rect 119476 35084 119980 35140
rect 120036 35084 122668 35140
rect 122724 35084 124012 35140
rect 124068 35084 124078 35140
rect 126466 35084 126476 35140
rect 126532 35084 127708 35140
rect 127764 35084 127774 35140
rect 131842 35084 131852 35140
rect 131908 35084 133644 35140
rect 133700 35084 133710 35140
rect 135426 35084 135436 35140
rect 135492 35084 136332 35140
rect 136388 35084 136398 35140
rect 139122 35084 139132 35140
rect 139188 35084 140700 35140
rect 140756 35084 140766 35140
rect 9874 34972 9884 35028
rect 9940 34972 10332 35028
rect 10388 34972 10398 35028
rect 11666 34972 11676 35028
rect 11732 34972 31948 35028
rect 36978 34972 36988 35028
rect 37044 34972 37884 35028
rect 37940 34972 37950 35028
rect 38434 34972 38444 35028
rect 38500 34972 39452 35028
rect 39508 34972 43708 35028
rect 47506 34972 47516 35028
rect 47572 34972 48300 35028
rect 48356 34972 49588 35028
rect 50306 34972 50316 35028
rect 50372 34972 50876 35028
rect 50932 34972 50942 35028
rect 73602 34972 73612 35028
rect 73668 34972 74508 35028
rect 74564 34972 74574 35028
rect 78932 34972 109228 35028
rect 31892 34916 31948 34972
rect 10770 34860 10780 34916
rect 10836 34860 19852 34916
rect 19908 34860 19918 34916
rect 31892 34860 39788 34916
rect 39844 34860 39854 34916
rect 43652 34804 43708 34972
rect 49532 34916 49588 34972
rect 78932 34916 78988 34972
rect 45602 34860 45612 34916
rect 45668 34860 47292 34916
rect 47348 34860 47852 34916
rect 47908 34860 47918 34916
rect 49522 34860 49532 34916
rect 49588 34860 50428 34916
rect 50484 34860 50494 34916
rect 55346 34860 55356 34916
rect 55412 34860 61292 34916
rect 61348 34860 61358 34916
rect 74162 34860 74172 34916
rect 74228 34860 78988 34916
rect 92978 34860 92988 34916
rect 93044 34860 95900 34916
rect 95956 34860 95966 34916
rect 98802 34860 98812 34916
rect 98868 34860 101164 34916
rect 101220 34860 101230 34916
rect 8866 34748 8876 34804
rect 8932 34748 17836 34804
rect 17892 34748 18956 34804
rect 19012 34748 19022 34804
rect 31490 34748 31500 34804
rect 31556 34748 32844 34804
rect 32900 34748 33292 34804
rect 33348 34748 33358 34804
rect 36642 34748 36652 34804
rect 36708 34748 37660 34804
rect 37716 34748 37726 34804
rect 43652 34748 49588 34804
rect 51986 34748 51996 34804
rect 52052 34748 56700 34804
rect 56756 34748 56766 34804
rect 59490 34748 59500 34804
rect 59556 34748 59836 34804
rect 59892 34748 59902 34804
rect 66556 34748 67116 34804
rect 67172 34748 67340 34804
rect 67396 34748 67406 34804
rect 73266 34748 73276 34804
rect 73332 34748 78204 34804
rect 78260 34748 78270 34804
rect 78530 34748 78540 34804
rect 78596 34748 79436 34804
rect 79492 34748 80444 34804
rect 80500 34748 80510 34804
rect 82562 34748 82572 34804
rect 82628 34748 83804 34804
rect 83860 34748 83870 34804
rect 88610 34748 88620 34804
rect 88676 34748 98588 34804
rect 98644 34748 98924 34804
rect 98980 34748 98990 34804
rect 102274 34748 102284 34804
rect 102340 34748 103628 34804
rect 103684 34748 103694 34804
rect 104738 34748 104748 34804
rect 104804 34748 106092 34804
rect 106148 34748 106158 34804
rect 6626 34636 6636 34692
rect 6692 34636 15596 34692
rect 15652 34636 16156 34692
rect 16212 34636 16222 34692
rect 16482 34636 16492 34692
rect 16548 34636 18396 34692
rect 18452 34636 18462 34692
rect 19730 34636 19740 34692
rect 19796 34636 20748 34692
rect 20804 34636 24220 34692
rect 24276 34636 24286 34692
rect 33170 34636 33180 34692
rect 33236 34636 33964 34692
rect 34020 34636 43708 34692
rect 44706 34636 44716 34692
rect 44772 34636 47068 34692
rect 47124 34636 47134 34692
rect 47394 34636 47404 34692
rect 47460 34636 48972 34692
rect 49028 34636 49038 34692
rect 14914 34524 14924 34580
rect 14980 34524 35644 34580
rect 35700 34524 36204 34580
rect 36260 34524 36270 34580
rect 38022 34468 38032 34524
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38296 34468 38306 34524
rect 43652 34468 43708 34636
rect 49532 34468 49588 34748
rect 56242 34636 56252 34692
rect 56308 34636 57036 34692
rect 57092 34636 57102 34692
rect 66556 34580 66612 34748
rect 109172 34692 109228 34972
rect 113372 34804 113428 35084
rect 115042 34972 115052 35028
rect 115108 34972 140644 35028
rect 140802 34972 140812 35028
rect 140868 34972 141708 35028
rect 141764 34972 141774 35028
rect 113810 34860 113820 34916
rect 113876 34860 114604 34916
rect 114660 34860 115388 34916
rect 115444 34860 115454 34916
rect 124002 34860 124012 34916
rect 124068 34860 128828 34916
rect 128884 34860 129388 34916
rect 129444 34860 130060 34916
rect 130116 34860 130508 34916
rect 130564 34860 130574 34916
rect 113372 34748 119420 34804
rect 119476 34748 119486 34804
rect 132066 34748 132076 34804
rect 132132 34748 132972 34804
rect 133028 34748 133038 34804
rect 136322 34748 136332 34804
rect 136388 34748 138012 34804
rect 138068 34748 138078 34804
rect 138562 34748 138572 34804
rect 138628 34748 139692 34804
rect 139748 34748 139758 34804
rect 138572 34692 138628 34748
rect 66770 34636 66780 34692
rect 66836 34636 67900 34692
rect 67956 34636 68572 34692
rect 68628 34636 69468 34692
rect 69524 34636 76076 34692
rect 76132 34636 76142 34692
rect 88498 34636 88508 34692
rect 88564 34636 89628 34692
rect 89684 34636 89694 34692
rect 109172 34636 115052 34692
rect 115108 34636 115118 34692
rect 115266 34636 115276 34692
rect 115332 34636 116956 34692
rect 117012 34636 117022 34692
rect 127586 34636 127596 34692
rect 127652 34636 129276 34692
rect 129332 34636 129948 34692
rect 130004 34636 130014 34692
rect 133644 34636 137340 34692
rect 137396 34636 138628 34692
rect 140588 34692 140644 34972
rect 143490 34748 143500 34804
rect 143556 34748 144732 34804
rect 144788 34748 144798 34804
rect 140588 34636 144620 34692
rect 144676 34636 145292 34692
rect 145348 34636 145628 34692
rect 145684 34636 145694 34692
rect 52882 34524 52892 34580
rect 52948 34524 66612 34580
rect 76178 34524 76188 34580
rect 76244 34524 76860 34580
rect 76916 34524 78988 34580
rect 79044 34524 79054 34580
rect 88946 34524 88956 34580
rect 89012 34524 90524 34580
rect 90580 34524 91308 34580
rect 91364 34524 91374 34580
rect 92418 34524 92428 34580
rect 92484 34524 105196 34580
rect 105252 34524 105262 34580
rect 113474 34524 113484 34580
rect 113540 34524 119084 34580
rect 119140 34524 119150 34580
rect 74842 34468 74852 34524
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 75116 34468 75126 34524
rect 111662 34468 111672 34524
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111936 34468 111946 34524
rect 16818 34412 16828 34468
rect 16884 34412 18564 34468
rect 19842 34412 19852 34468
rect 19908 34412 21532 34468
rect 21588 34412 21868 34468
rect 21924 34412 21934 34468
rect 24434 34412 24444 34468
rect 24500 34412 24780 34468
rect 24836 34412 37100 34468
rect 37156 34412 37166 34468
rect 43652 34412 46396 34468
rect 46452 34412 46462 34468
rect 49532 34412 61348 34468
rect 62402 34412 62412 34468
rect 62468 34412 73556 34468
rect 75730 34412 75740 34468
rect 75796 34412 82236 34468
rect 82292 34412 82302 34468
rect 103170 34412 103180 34468
rect 103236 34412 103852 34468
rect 103908 34412 103918 34468
rect 107426 34412 107436 34468
rect 107492 34412 110964 34468
rect 18508 34356 18564 34412
rect 61292 34356 61348 34412
rect 73500 34356 73556 34412
rect 110908 34356 110964 34412
rect 113484 34356 113540 34524
rect 15026 34300 15036 34356
rect 15092 34300 15932 34356
rect 15988 34300 15998 34356
rect 16930 34300 16940 34356
rect 16996 34300 18284 34356
rect 18340 34300 18350 34356
rect 18508 34300 29372 34356
rect 29428 34300 30604 34356
rect 30660 34300 30670 34356
rect 32834 34300 32844 34356
rect 32900 34300 33516 34356
rect 33572 34300 46060 34356
rect 46116 34300 46126 34356
rect 48178 34300 48188 34356
rect 48244 34300 48748 34356
rect 48804 34300 57484 34356
rect 57540 34300 57550 34356
rect 61292 34300 66556 34356
rect 66612 34300 66622 34356
rect 68226 34300 68236 34356
rect 68292 34300 69916 34356
rect 69972 34300 69982 34356
rect 73500 34300 76300 34356
rect 76356 34300 76860 34356
rect 76916 34300 76926 34356
rect 77074 34300 77084 34356
rect 77140 34300 81620 34356
rect 81778 34300 81788 34356
rect 81844 34300 82684 34356
rect 82740 34300 82750 34356
rect 87602 34300 87612 34356
rect 87668 34300 88396 34356
rect 88452 34300 88462 34356
rect 90290 34300 90300 34356
rect 90356 34300 93772 34356
rect 93828 34300 93838 34356
rect 108994 34300 109004 34356
rect 109060 34300 109564 34356
rect 109620 34300 109630 34356
rect 110898 34300 110908 34356
rect 110964 34300 113540 34356
rect 113596 34412 131516 34468
rect 131572 34412 131740 34468
rect 131796 34412 131806 34468
rect 81564 34244 81620 34300
rect 19954 34188 19964 34244
rect 20020 34188 20748 34244
rect 20804 34188 20814 34244
rect 22866 34188 22876 34244
rect 22932 34188 23212 34244
rect 23268 34188 36988 34244
rect 37044 34188 37054 34244
rect 39890 34188 39900 34244
rect 39956 34188 40460 34244
rect 40516 34188 40526 34244
rect 48514 34188 48524 34244
rect 48580 34188 49644 34244
rect 49700 34188 49710 34244
rect 50754 34188 50764 34244
rect 50820 34188 54124 34244
rect 54180 34188 54190 34244
rect 54562 34188 54572 34244
rect 54628 34188 78988 34244
rect 81564 34188 88620 34244
rect 88676 34188 90412 34244
rect 90468 34188 90478 34244
rect 92306 34188 92316 34244
rect 92372 34188 102620 34244
rect 102676 34188 103180 34244
rect 103236 34188 103246 34244
rect 105410 34188 105420 34244
rect 105476 34188 106316 34244
rect 106372 34188 106652 34244
rect 106708 34188 111916 34244
rect 111972 34188 111982 34244
rect 78932 34132 78988 34188
rect 113596 34132 113652 34412
rect 117170 34300 117180 34356
rect 117236 34300 117740 34356
rect 117796 34300 117806 34356
rect 133644 34244 133700 34636
rect 148482 34468 148492 34524
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148756 34468 148766 34524
rect 137330 34412 137340 34468
rect 137396 34412 139020 34468
rect 139076 34412 139086 34468
rect 133858 34300 133868 34356
rect 133924 34300 135660 34356
rect 135716 34300 135726 34356
rect 113810 34188 113820 34244
rect 113876 34188 133700 34244
rect 136994 34188 137004 34244
rect 137060 34188 138348 34244
rect 138404 34188 138414 34244
rect 142370 34188 142380 34244
rect 142436 34188 143052 34244
rect 143108 34188 143118 34244
rect 40786 34076 40796 34132
rect 40852 34076 44604 34132
rect 44660 34076 44670 34132
rect 67330 34076 67340 34132
rect 67396 34076 68236 34132
rect 68292 34076 71148 34132
rect 71204 34076 71214 34132
rect 73490 34076 73500 34132
rect 73556 34076 74172 34132
rect 74228 34076 74238 34132
rect 78932 34076 83804 34132
rect 83860 34076 84140 34132
rect 84196 34076 84206 34132
rect 90850 34076 90860 34132
rect 90916 34076 92428 34132
rect 92484 34076 92494 34132
rect 98018 34076 98028 34132
rect 98084 34076 109228 34132
rect 109284 34076 109294 34132
rect 110226 34076 110236 34132
rect 110292 34076 110460 34132
rect 110516 34076 113652 34132
rect 114146 34076 114156 34132
rect 114212 34076 115052 34132
rect 115108 34076 115118 34132
rect 127474 34076 127484 34132
rect 127540 34076 131292 34132
rect 131348 34076 131358 34132
rect 137442 34076 137452 34132
rect 137508 34076 140028 34132
rect 140084 34076 140094 34132
rect 141810 34076 141820 34132
rect 141876 34076 142940 34132
rect 142996 34076 143006 34132
rect 14578 33964 14588 34020
rect 14644 33964 15036 34020
rect 15092 33964 23884 34020
rect 23940 33964 24892 34020
rect 24948 33964 25788 34020
rect 25844 33964 25854 34020
rect 28354 33964 28364 34020
rect 28420 33964 28588 34020
rect 28644 33964 28654 34020
rect 33282 33964 33292 34020
rect 33348 33964 58268 34020
rect 58324 33964 58604 34020
rect 58660 33964 58670 34020
rect 65650 33964 65660 34020
rect 65716 33964 69468 34020
rect 69524 33964 69534 34020
rect 88162 33964 88172 34020
rect 88228 33964 89628 34020
rect 89684 33964 89694 34020
rect 91074 33964 91084 34020
rect 91140 33964 91868 34020
rect 91924 33964 93828 34020
rect 96898 33964 96908 34020
rect 96964 33964 97916 34020
rect 97972 33964 97982 34020
rect 99474 33964 99484 34020
rect 99540 33964 100492 34020
rect 100548 33964 100558 34020
rect 104962 33964 104972 34020
rect 105028 33964 105868 34020
rect 105924 33964 105934 34020
rect 106754 33964 106764 34020
rect 106820 33964 107660 34020
rect 107716 33964 107726 34020
rect 107874 33964 107884 34020
rect 107940 33964 108668 34020
rect 108724 33964 108734 34020
rect 112466 33964 112476 34020
rect 112532 33964 113372 34020
rect 113428 33964 113438 34020
rect 115714 33964 115724 34020
rect 115780 33964 116620 34020
rect 116676 33964 116686 34020
rect 122882 33964 122892 34020
rect 122948 33964 123788 34020
rect 123844 33964 123854 34020
rect 126018 33964 126028 34020
rect 126084 33964 129948 34020
rect 130004 33964 130620 34020
rect 130676 33964 130686 34020
rect 144386 33964 144396 34020
rect 144452 33964 145628 34020
rect 145684 33964 145694 34020
rect 93772 33908 93828 33964
rect 8082 33852 8092 33908
rect 8148 33852 8540 33908
rect 8596 33852 29484 33908
rect 29540 33852 29820 33908
rect 29876 33852 29886 33908
rect 34514 33852 34524 33908
rect 34580 33852 43596 33908
rect 43652 33852 43662 33908
rect 49746 33852 49756 33908
rect 49812 33852 50764 33908
rect 50820 33852 50830 33908
rect 55412 33852 56868 33908
rect 59490 33852 59500 33908
rect 59556 33852 61964 33908
rect 62020 33852 62030 33908
rect 63634 33852 63644 33908
rect 63700 33852 63980 33908
rect 64036 33852 65100 33908
rect 65156 33852 75068 33908
rect 75124 33852 75740 33908
rect 75796 33852 75806 33908
rect 80434 33852 80444 33908
rect 80500 33852 93716 33908
rect 93772 33852 110572 33908
rect 110628 33852 110638 33908
rect 111906 33852 111916 33908
rect 111972 33852 113148 33908
rect 113204 33852 113214 33908
rect 130722 33852 130732 33908
rect 130788 33852 137340 33908
rect 137396 33852 137406 33908
rect 26002 33740 26012 33796
rect 26068 33740 41580 33796
rect 41636 33740 42140 33796
rect 42196 33740 42206 33796
rect 43586 33740 43596 33796
rect 43652 33740 51436 33796
rect 51492 33740 51502 33796
rect 51762 33740 51772 33796
rect 51828 33740 52444 33796
rect 52500 33740 52510 33796
rect 19612 33684 19622 33740
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19886 33684 19896 33740
rect 55412 33684 55468 33852
rect 56432 33684 56442 33740
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56706 33684 56716 33740
rect 56812 33684 56868 33852
rect 93660 33796 93716 33852
rect 58482 33740 58492 33796
rect 58548 33740 59612 33796
rect 59668 33740 59678 33796
rect 93660 33740 105644 33796
rect 105700 33740 105710 33796
rect 112018 33740 112028 33796
rect 112084 33740 113820 33796
rect 113876 33740 113886 33796
rect 93252 33684 93262 33740
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93526 33684 93536 33740
rect 130072 33684 130082 33740
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130346 33684 130356 33740
rect 41010 33628 41020 33684
rect 41076 33628 41804 33684
rect 41860 33628 43148 33684
rect 43204 33628 43214 33684
rect 43586 33628 43596 33684
rect 43652 33628 55468 33684
rect 56812 33628 87612 33684
rect 87668 33628 87678 33684
rect 94098 33628 94108 33684
rect 94164 33628 94556 33684
rect 94612 33628 94622 33684
rect 32610 33516 32620 33572
rect 32676 33516 38444 33572
rect 38500 33516 38510 33572
rect 41906 33516 41916 33572
rect 41972 33516 42140 33572
rect 42196 33516 42206 33572
rect 42354 33516 42364 33572
rect 42420 33516 47964 33572
rect 48020 33516 48030 33572
rect 51314 33516 51324 33572
rect 51380 33516 52556 33572
rect 52612 33516 52622 33572
rect 58706 33516 58716 33572
rect 58772 33516 59164 33572
rect 59220 33516 59230 33572
rect 64418 33516 64428 33572
rect 64484 33516 64764 33572
rect 64820 33516 64830 33572
rect 88834 33516 88844 33572
rect 88900 33516 90748 33572
rect 90804 33516 90814 33572
rect 106866 33516 106876 33572
rect 106932 33516 107660 33572
rect 107716 33516 109228 33572
rect 112130 33516 112140 33572
rect 112196 33516 113036 33572
rect 113092 33516 113102 33572
rect 118514 33516 118524 33572
rect 118580 33516 119084 33572
rect 119140 33516 119150 33572
rect 109172 33460 109228 33516
rect 30034 33404 30044 33460
rect 30100 33404 31836 33460
rect 31892 33404 31902 33460
rect 36082 33404 36092 33460
rect 36148 33404 36764 33460
rect 36820 33404 51212 33460
rect 51268 33404 51278 33460
rect 53554 33404 53564 33460
rect 53620 33404 53900 33460
rect 53956 33404 70252 33460
rect 70308 33404 70318 33460
rect 77746 33404 77756 33460
rect 77812 33404 85708 33460
rect 88050 33404 88060 33460
rect 88116 33404 89068 33460
rect 89124 33404 89134 33460
rect 93986 33404 93996 33460
rect 94052 33404 95228 33460
rect 95284 33404 95294 33460
rect 109172 33404 132860 33460
rect 132916 33404 132926 33460
rect 137218 33404 137228 33460
rect 137284 33404 138124 33460
rect 138180 33404 138190 33460
rect 139234 33404 139244 33460
rect 139300 33404 139580 33460
rect 139636 33404 139646 33460
rect 85652 33348 85708 33404
rect 28802 33292 28812 33348
rect 28868 33292 48860 33348
rect 48916 33292 48926 33348
rect 65986 33292 65996 33348
rect 66052 33292 66668 33348
rect 66724 33292 66734 33348
rect 85652 33292 95116 33348
rect 95172 33292 95182 33348
rect 108210 33292 108220 33348
rect 108276 33292 112364 33348
rect 112420 33292 112430 33348
rect 119074 33292 119084 33348
rect 119140 33292 131964 33348
rect 132020 33292 132300 33348
rect 132356 33292 132366 33348
rect 135090 33292 135100 33348
rect 135156 33292 137452 33348
rect 137508 33292 137518 33348
rect 18162 33180 18172 33236
rect 18228 33180 35028 33236
rect 38098 33180 38108 33236
rect 38164 33180 38668 33236
rect 38724 33180 38734 33236
rect 49186 33180 49196 33236
rect 49252 33180 49420 33236
rect 49476 33180 80556 33236
rect 80612 33180 81340 33236
rect 81396 33180 81406 33236
rect 117842 33180 117852 33236
rect 117908 33180 118412 33236
rect 118468 33180 118478 33236
rect 118738 33180 118748 33236
rect 118804 33180 126588 33236
rect 126644 33180 126654 33236
rect 19730 33068 19740 33124
rect 19796 33068 26012 33124
rect 26068 33068 26078 33124
rect 30818 33068 30828 33124
rect 30884 33068 32620 33124
rect 32676 33068 32686 33124
rect 19058 32956 19068 33012
rect 19124 32956 20524 33012
rect 20580 32956 22092 33012
rect 22148 32956 31948 33012
rect 32004 32956 32014 33012
rect 31266 32844 31276 32900
rect 31332 32844 31836 32900
rect 31892 32844 32284 32900
rect 32340 32844 32350 32900
rect 34972 32788 35028 33180
rect 35186 33068 35196 33124
rect 35252 33068 42364 33124
rect 42420 33068 42430 33124
rect 45378 33068 45388 33124
rect 45444 33068 49868 33124
rect 49924 33068 49934 33124
rect 63410 33068 63420 33124
rect 63476 33068 63868 33124
rect 63924 33068 63934 33124
rect 65874 33068 65884 33124
rect 65940 33068 66668 33124
rect 66724 33068 66734 33124
rect 67172 33068 77644 33124
rect 77700 33068 77710 33124
rect 93986 33068 93996 33124
rect 94052 33068 94780 33124
rect 94836 33068 95004 33124
rect 95060 33068 95070 33124
rect 119634 33068 119644 33124
rect 119700 33068 120092 33124
rect 120148 33068 120158 33124
rect 123890 33068 123900 33124
rect 123956 33068 124908 33124
rect 124964 33068 138796 33124
rect 138852 33068 139244 33124
rect 139300 33068 139310 33124
rect 67172 33012 67228 33068
rect 42130 32956 42140 33012
rect 42196 32956 67228 33012
rect 67330 32956 67340 33012
rect 67396 32956 73332 33012
rect 84578 32956 84588 33012
rect 84644 32956 106652 33012
rect 106708 32956 106718 33012
rect 38022 32900 38032 32956
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38296 32900 38306 32956
rect 38434 32844 38444 32900
rect 38500 32844 39004 32900
rect 39060 32844 39228 32900
rect 39284 32844 39294 32900
rect 51538 32844 51548 32900
rect 51604 32844 51996 32900
rect 52052 32844 58828 32900
rect 58884 32844 72884 32900
rect 34972 32732 40460 32788
rect 40516 32732 41244 32788
rect 41300 32732 41310 32788
rect 41468 32732 57148 32788
rect 57204 32732 57214 32788
rect 62290 32732 62300 32788
rect 62356 32732 63196 32788
rect 63252 32732 63262 32788
rect 64530 32732 64540 32788
rect 64596 32732 67228 32788
rect 67284 32732 67294 32788
rect 41468 32676 41524 32732
rect 72828 32676 72884 32844
rect 73276 32788 73332 32956
rect 74842 32900 74852 32956
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 75116 32900 75126 32956
rect 111662 32900 111672 32956
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111936 32900 111946 32956
rect 148482 32900 148492 32956
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148756 32900 148766 32956
rect 73276 32732 96012 32788
rect 96068 32732 96078 32788
rect 100258 32732 100268 32788
rect 100324 32732 102396 32788
rect 102452 32732 125580 32788
rect 125636 32732 125646 32788
rect 131058 32732 131068 32788
rect 131124 32732 147868 32788
rect 147924 32732 147934 32788
rect 9874 32620 9884 32676
rect 9940 32620 11676 32676
rect 11732 32620 37884 32676
rect 37940 32620 37950 32676
rect 38434 32620 38444 32676
rect 38500 32620 41524 32676
rect 43652 32620 61516 32676
rect 61572 32620 61582 32676
rect 72828 32620 82236 32676
rect 82292 32620 82302 32676
rect 90066 32620 90076 32676
rect 90132 32620 91644 32676
rect 91700 32620 116844 32676
rect 116900 32620 116910 32676
rect 43652 32564 43708 32620
rect 38994 32508 39004 32564
rect 39060 32508 40796 32564
rect 40852 32508 43708 32564
rect 48514 32508 48524 32564
rect 48580 32508 58828 32564
rect 58884 32508 91980 32564
rect 92036 32508 92046 32564
rect 95218 32508 95228 32564
rect 95284 32508 115612 32564
rect 115668 32508 115678 32564
rect 78932 32396 91756 32452
rect 91812 32396 93548 32452
rect 93604 32396 93614 32452
rect 118738 32396 118748 32452
rect 118804 32396 118972 32452
rect 119028 32396 141820 32452
rect 141876 32396 141886 32452
rect 78932 32340 78988 32396
rect 31378 32284 31388 32340
rect 31444 32284 39564 32340
rect 39620 32284 39630 32340
rect 54236 32284 78988 32340
rect 85652 32284 105756 32340
rect 105812 32284 113596 32340
rect 113652 32284 114044 32340
rect 114100 32284 114110 32340
rect 19612 32116 19622 32172
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19886 32116 19896 32172
rect 54236 32116 54292 32284
rect 85652 32228 85708 32284
rect 61842 32172 61852 32228
rect 61908 32172 85708 32228
rect 56432 32116 56442 32172
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56706 32116 56716 32172
rect 93252 32116 93262 32172
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93526 32116 93536 32172
rect 130072 32116 130082 32172
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130346 32116 130356 32172
rect 46946 32060 46956 32116
rect 47012 32060 54236 32116
rect 54292 32060 54302 32116
rect 34850 31948 34860 32004
rect 34916 31948 64428 32004
rect 64484 31948 64494 32004
rect 66658 31948 66668 32004
rect 66724 31948 67508 32004
rect 70802 31948 70812 32004
rect 70868 31948 105756 32004
rect 105812 31948 107996 32004
rect 108052 31948 108062 32004
rect 7186 31836 7196 31892
rect 7252 31836 31948 31892
rect 40114 31836 40124 31892
rect 40180 31836 45052 31892
rect 45108 31836 45118 31892
rect 63298 31836 63308 31892
rect 63364 31836 64876 31892
rect 64932 31836 64942 31892
rect 31892 31780 31948 31836
rect 67452 31780 67508 31948
rect 71922 31836 71932 31892
rect 71988 31836 123564 31892
rect 123620 31836 123630 31892
rect 31892 31724 45388 31780
rect 45444 31724 45454 31780
rect 51874 31724 51884 31780
rect 51940 31724 52556 31780
rect 52612 31724 62972 31780
rect 63028 31724 63038 31780
rect 67452 31724 119196 31780
rect 119252 31724 119262 31780
rect 58930 31612 58940 31668
rect 58996 31612 93996 31668
rect 94052 31612 94062 31668
rect 94882 31612 94892 31668
rect 94948 31612 144844 31668
rect 144900 31612 144910 31668
rect 105746 31500 105756 31556
rect 105812 31500 107548 31556
rect 107604 31500 107614 31556
rect 38022 31332 38032 31388
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38296 31332 38306 31388
rect 74842 31332 74852 31388
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 75116 31332 75126 31388
rect 111662 31332 111672 31388
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111936 31332 111946 31388
rect 148482 31332 148492 31388
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148756 31332 148766 31388
rect 77186 31276 77196 31332
rect 77252 31276 102732 31332
rect 102788 31276 102798 31332
rect 44594 31164 44604 31220
rect 44660 31164 82012 31220
rect 82068 31164 82078 31220
rect 31938 31052 31948 31108
rect 32004 31052 60396 31108
rect 60452 31052 60462 31108
rect 131618 31052 131628 31108
rect 131684 31052 147980 31108
rect 148036 31052 148046 31108
rect 60722 30940 60732 30996
rect 60788 30940 99036 30996
rect 99092 30940 99102 30996
rect 60834 30828 60844 30884
rect 60900 30828 87724 30884
rect 87780 30828 87790 30884
rect 19612 30548 19622 30604
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19886 30548 19896 30604
rect 56432 30548 56442 30604
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56706 30548 56716 30604
rect 93252 30548 93262 30604
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93526 30548 93536 30604
rect 130072 30548 130082 30604
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130346 30548 130356 30604
rect 60386 30268 60396 30324
rect 60452 30268 61740 30324
rect 61796 30268 61806 30324
rect 59042 30156 59052 30212
rect 59108 30156 127596 30212
rect 127652 30156 127662 30212
rect 69458 30044 69468 30100
rect 69524 30044 104300 30100
rect 104356 30044 104366 30100
rect 22194 29932 22204 29988
rect 22260 29932 81452 29988
rect 81508 29932 81518 29988
rect 38022 29764 38032 29820
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38296 29764 38306 29820
rect 74842 29764 74852 29820
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 75116 29764 75126 29820
rect 111662 29764 111672 29820
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111936 29764 111946 29820
rect 148482 29764 148492 29820
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148756 29764 148766 29820
rect 18386 29596 18396 29652
rect 18452 29596 79100 29652
rect 79156 29596 79166 29652
rect 64978 29484 64988 29540
rect 65044 29484 112476 29540
rect 112532 29484 112542 29540
rect 40898 29260 40908 29316
rect 40964 29260 92204 29316
rect 92260 29260 92270 29316
rect 19612 28980 19622 29036
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19886 28980 19896 29036
rect 56432 28980 56442 29036
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56706 28980 56716 29036
rect 93252 28980 93262 29036
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93526 28980 93536 29036
rect 130072 28980 130082 29036
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130346 28980 130356 29036
rect 104962 28588 104972 28644
rect 105028 28588 105756 28644
rect 105812 28588 105822 28644
rect 72370 28476 72380 28532
rect 72436 28476 142380 28532
rect 142436 28476 142446 28532
rect 71474 28364 71484 28420
rect 71540 28364 133084 28420
rect 133140 28364 133150 28420
rect 38022 28196 38032 28252
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38296 28196 38306 28252
rect 74842 28196 74852 28252
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 75116 28196 75126 28252
rect 111662 28196 111672 28252
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111936 28196 111946 28252
rect 148482 28196 148492 28252
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148756 28196 148766 28252
rect 47170 28028 47180 28084
rect 47236 28028 88956 28084
rect 89012 28028 89022 28084
rect 51650 27916 51660 27972
rect 51716 27916 85148 27972
rect 85204 27916 85214 27972
rect 39106 27804 39116 27860
rect 39172 27804 79772 27860
rect 79828 27804 79838 27860
rect 37650 27692 37660 27748
rect 37716 27692 42812 27748
rect 42868 27692 64316 27748
rect 64372 27692 64382 27748
rect 92642 27692 92652 27748
rect 92708 27692 126812 27748
rect 126868 27692 126878 27748
rect 24210 27580 24220 27636
rect 24276 27580 79660 27636
rect 79716 27580 79726 27636
rect 19612 27412 19622 27468
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19886 27412 19896 27468
rect 56432 27412 56442 27468
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56706 27412 56716 27468
rect 93252 27412 93262 27468
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93526 27412 93536 27468
rect 130072 27412 130082 27468
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130346 27412 130356 27468
rect 36530 27244 36540 27300
rect 36596 27244 87500 27300
rect 87556 27244 87566 27300
rect 42466 27132 42476 27188
rect 42532 27132 89740 27188
rect 89796 27132 89806 27188
rect 75506 26908 75516 26964
rect 75572 26908 76636 26964
rect 76692 26908 76702 26964
rect 59714 26796 59724 26852
rect 59780 26796 137004 26852
rect 137060 26796 137070 26852
rect 38022 26628 38032 26684
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38296 26628 38306 26684
rect 74842 26628 74852 26684
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 75116 26628 75126 26684
rect 111662 26628 111672 26684
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111936 26628 111946 26684
rect 148482 26628 148492 26684
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148756 26628 148766 26684
rect 28466 26460 28476 26516
rect 28532 26460 87052 26516
rect 87108 26460 87118 26516
rect 47282 26348 47292 26404
rect 47348 26348 99708 26404
rect 99764 26348 99774 26404
rect 57922 26236 57932 26292
rect 57988 26236 94220 26292
rect 94276 26236 94286 26292
rect 98242 26236 98252 26292
rect 98308 26236 124796 26292
rect 124852 26236 124862 26292
rect 26114 26124 26124 26180
rect 26180 26124 85484 26180
rect 85540 26124 85550 26180
rect 106642 26124 106652 26180
rect 106708 26124 117628 26180
rect 117684 26124 117694 26180
rect 120082 26124 120092 26180
rect 120148 26124 125132 26180
rect 125188 26124 133196 26180
rect 133252 26124 133262 26180
rect 18498 26012 18508 26068
rect 18564 26012 20076 26068
rect 20132 26012 20142 26068
rect 120978 26012 120988 26068
rect 121044 26012 122444 26068
rect 122500 26012 122510 26068
rect 19612 25844 19622 25900
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19886 25844 19896 25900
rect 56432 25844 56442 25900
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56706 25844 56716 25900
rect 93252 25844 93262 25900
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93526 25844 93536 25900
rect 130072 25844 130082 25900
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130346 25844 130356 25900
rect 55682 25676 55692 25732
rect 55748 25676 126028 25732
rect 126084 25676 126094 25732
rect 58818 25116 58828 25172
rect 58884 25116 62636 25172
rect 62692 25116 62702 25172
rect 38022 25060 38032 25116
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38296 25060 38306 25116
rect 74842 25060 74852 25116
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 75116 25060 75126 25116
rect 111662 25060 111672 25116
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111936 25060 111946 25116
rect 148482 25060 148492 25116
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148756 25060 148766 25116
rect 31826 24892 31836 24948
rect 31892 24892 89516 24948
rect 89572 24892 89582 24948
rect 42018 24780 42028 24836
rect 42084 24780 92876 24836
rect 92932 24780 92942 24836
rect 30146 24668 30156 24724
rect 30212 24668 77980 24724
rect 78036 24668 78046 24724
rect 52098 24556 52108 24612
rect 52164 24556 119308 24612
rect 119364 24556 119374 24612
rect 89618 24444 89628 24500
rect 89684 24444 108556 24500
rect 108612 24444 108622 24500
rect 62178 24332 62188 24388
rect 62244 24332 80668 24388
rect 80724 24332 80734 24388
rect 101826 24332 101836 24388
rect 101892 24332 107548 24388
rect 107604 24332 107614 24388
rect 19612 24276 19622 24332
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19886 24276 19896 24332
rect 56432 24276 56442 24332
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56706 24276 56716 24332
rect 93252 24276 93262 24332
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93526 24276 93536 24332
rect 130072 24276 130082 24332
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130346 24276 130356 24332
rect 61618 24108 61628 24164
rect 61684 24108 135996 24164
rect 136052 24108 136062 24164
rect 38022 23492 38032 23548
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38296 23492 38306 23548
rect 74842 23492 74852 23548
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 75116 23492 75126 23548
rect 111662 23492 111672 23548
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111936 23492 111946 23548
rect 148482 23492 148492 23548
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148756 23492 148766 23548
rect 49186 23436 49196 23492
rect 49252 23436 52892 23492
rect 52948 23436 52958 23492
rect 45042 23324 45052 23380
rect 45108 23324 98588 23380
rect 98644 23324 98654 23380
rect 60386 23212 60396 23268
rect 60452 23212 105420 23268
rect 105476 23212 105486 23268
rect 58594 23100 58604 23156
rect 58660 23100 89404 23156
rect 89460 23100 89470 23156
rect 45826 22988 45836 23044
rect 45892 22988 61740 23044
rect 61796 22988 61806 23044
rect 79762 22988 79772 23044
rect 79828 22988 107884 23044
rect 107940 22988 107950 23044
rect 52434 22876 52444 22932
rect 52500 22876 71708 22932
rect 71764 22876 71774 22932
rect 86482 22876 86492 22932
rect 86548 22876 117404 22932
rect 117460 22876 117470 22932
rect 19612 22708 19622 22764
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19886 22708 19896 22764
rect 56432 22708 56442 22764
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56706 22708 56716 22764
rect 93252 22708 93262 22764
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93526 22708 93536 22764
rect 130072 22708 130082 22764
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130346 22708 130356 22764
rect 102386 22652 102396 22708
rect 102452 22652 113260 22708
rect 113316 22652 113326 22708
rect 54338 22540 54348 22596
rect 54404 22540 121772 22596
rect 121828 22540 121838 22596
rect 38022 21924 38032 21980
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38296 21924 38306 21980
rect 74842 21924 74852 21980
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 75116 21924 75126 21980
rect 111662 21924 111672 21980
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111936 21924 111946 21980
rect 148482 21924 148492 21980
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148756 21924 148766 21980
rect 133634 21756 133644 21812
rect 133700 21756 134428 21812
rect 134484 21756 134494 21812
rect 54898 21308 54908 21364
rect 54964 21308 84924 21364
rect 84980 21308 84990 21364
rect 19612 21140 19622 21196
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19886 21140 19896 21196
rect 56432 21140 56442 21196
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56706 21140 56716 21196
rect 93252 21140 93262 21196
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93526 21140 93536 21196
rect 130072 21140 130082 21196
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130346 21140 130356 21196
rect 83122 20972 83132 21028
rect 83188 20972 115276 21028
rect 115332 20972 115342 21028
rect 38022 20356 38032 20412
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38296 20356 38306 20412
rect 74842 20356 74852 20412
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 75116 20356 75126 20412
rect 111662 20356 111672 20412
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111936 20356 111946 20412
rect 148482 20356 148492 20412
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148756 20356 148766 20412
rect 45714 20076 45724 20132
rect 45780 20076 92988 20132
rect 93044 20076 93054 20132
rect 19612 19572 19622 19628
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19886 19572 19896 19628
rect 56432 19572 56442 19628
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56706 19572 56716 19628
rect 93252 19572 93262 19628
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93526 19572 93536 19628
rect 130072 19572 130082 19628
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130346 19572 130356 19628
rect 38022 18788 38032 18844
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38296 18788 38306 18844
rect 74842 18788 74852 18844
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 75116 18788 75126 18844
rect 111662 18788 111672 18844
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111936 18788 111946 18844
rect 148482 18788 148492 18844
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148756 18788 148766 18844
rect 19612 18004 19622 18060
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19886 18004 19896 18060
rect 56432 18004 56442 18060
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56706 18004 56716 18060
rect 93252 18004 93262 18060
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93526 18004 93536 18060
rect 130072 18004 130082 18060
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130346 18004 130356 18060
rect 17938 17612 17948 17668
rect 18004 17612 51324 17668
rect 51380 17612 51390 17668
rect 57026 17612 57036 17668
rect 57092 17612 92428 17668
rect 92484 17612 92494 17668
rect 38022 17220 38032 17276
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38296 17220 38306 17276
rect 74842 17220 74852 17276
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 75116 17220 75126 17276
rect 111662 17220 111672 17276
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111936 17220 111946 17276
rect 148482 17220 148492 17276
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148756 17220 148766 17276
rect 48962 16828 48972 16884
rect 49028 16828 51436 16884
rect 51492 16828 51502 16884
rect 19612 16436 19622 16492
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19886 16436 19896 16492
rect 56432 16436 56442 16492
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56706 16436 56716 16492
rect 93252 16436 93262 16492
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93526 16436 93536 16492
rect 130072 16436 130082 16492
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130346 16436 130356 16492
rect 35410 16044 35420 16100
rect 35476 16044 45276 16100
rect 45332 16044 45342 16100
rect 84914 15932 84924 15988
rect 84980 15932 88620 15988
rect 88676 15932 122108 15988
rect 122164 15932 122174 15988
rect 38022 15652 38032 15708
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38296 15652 38306 15708
rect 74842 15652 74852 15708
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 75116 15652 75126 15708
rect 111662 15652 111672 15708
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111936 15652 111946 15708
rect 148482 15652 148492 15708
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148756 15652 148766 15708
rect 38434 15036 38444 15092
rect 38500 15036 43932 15092
rect 43988 15036 43998 15092
rect 19612 14868 19622 14924
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19886 14868 19896 14924
rect 56432 14868 56442 14924
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56706 14868 56716 14924
rect 93252 14868 93262 14924
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93526 14868 93536 14924
rect 130072 14868 130082 14924
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130346 14868 130356 14924
rect 46498 14364 46508 14420
rect 46564 14364 58044 14420
rect 58100 14364 58110 14420
rect 57810 14252 57820 14308
rect 57876 14252 84700 14308
rect 84756 14252 86492 14308
rect 86548 14252 86558 14308
rect 38022 14084 38032 14140
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38296 14084 38306 14140
rect 74842 14084 74852 14140
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 75116 14084 75126 14140
rect 111662 14084 111672 14140
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111936 14084 111946 14140
rect 148482 14084 148492 14140
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148756 14084 148766 14140
rect 42130 13356 42140 13412
rect 42196 13356 46732 13412
rect 46788 13356 46798 13412
rect 113922 13356 113932 13412
rect 113988 13356 115724 13412
rect 115780 13356 115790 13412
rect 19612 13300 19622 13356
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19886 13300 19896 13356
rect 56432 13300 56442 13356
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56706 13300 56716 13356
rect 93252 13300 93262 13356
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93526 13300 93536 13356
rect 130072 13300 130082 13356
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130346 13300 130356 13356
rect 53666 12796 53676 12852
rect 53732 12796 75852 12852
rect 75908 12796 76972 12852
rect 77028 12796 77038 12852
rect 30482 12684 30492 12740
rect 30548 12684 39900 12740
rect 39956 12684 39966 12740
rect 71698 12684 71708 12740
rect 71764 12684 103740 12740
rect 103796 12684 103806 12740
rect 108546 12684 108556 12740
rect 108612 12684 114268 12740
rect 114212 12628 114268 12684
rect 114212 12572 128828 12628
rect 128884 12572 128894 12628
rect 38022 12516 38032 12572
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38296 12516 38306 12572
rect 74842 12516 74852 12572
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 75116 12516 75126 12572
rect 111662 12516 111672 12572
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111936 12516 111946 12572
rect 148482 12516 148492 12572
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148756 12516 148766 12572
rect 76962 11788 76972 11844
rect 77028 11788 79772 11844
rect 79828 11788 79838 11844
rect 19612 11732 19622 11788
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19886 11732 19896 11788
rect 56432 11732 56442 11788
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56706 11732 56716 11788
rect 93252 11732 93262 11788
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93526 11732 93536 11788
rect 130072 11732 130082 11788
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130346 11732 130356 11788
rect 73714 11676 73724 11732
rect 73780 11676 78428 11732
rect 78484 11676 78494 11732
rect 91410 11116 91420 11172
rect 91476 11116 126364 11172
rect 126420 11116 126430 11172
rect 38022 10948 38032 11004
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38296 10948 38306 11004
rect 74842 10948 74852 11004
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 75116 10948 75126 11004
rect 111662 10948 111672 11004
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111936 10948 111946 11004
rect 148482 10948 148492 11004
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148756 10948 148766 11004
rect 22306 10892 22316 10948
rect 22372 10892 34972 10948
rect 35028 10892 35038 10948
rect 40562 10892 40572 10948
rect 40628 10892 59836 10948
rect 59892 10892 59902 10948
rect 32946 10780 32956 10836
rect 33012 10780 41244 10836
rect 41300 10780 41310 10836
rect 19612 10164 19622 10220
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19886 10164 19896 10220
rect 56432 10164 56442 10220
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56706 10164 56716 10220
rect 93252 10164 93262 10220
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93526 10164 93536 10220
rect 130072 10164 130082 10220
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130346 10164 130356 10220
rect 24994 9996 25004 10052
rect 25060 9996 29484 10052
rect 29540 9996 29550 10052
rect 119186 9996 119196 10052
rect 119252 9996 120988 10052
rect 121044 9996 121054 10052
rect 126802 9884 126812 9940
rect 126868 9884 128716 9940
rect 128772 9884 129500 9940
rect 129556 9884 129566 9940
rect 38022 9380 38032 9436
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38296 9380 38306 9436
rect 74842 9380 74852 9436
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 75116 9380 75126 9436
rect 111662 9380 111672 9436
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111936 9380 111946 9436
rect 148482 9380 148492 9436
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148756 9380 148766 9436
rect 29810 9324 29820 9380
rect 29876 9324 35644 9380
rect 35700 9324 35710 9380
rect 34514 9212 34524 9268
rect 34580 9212 47068 9268
rect 47124 9212 47134 9268
rect 65986 9212 65996 9268
rect 66052 9212 67228 9268
rect 67284 9212 67294 9268
rect 64642 9100 64652 9156
rect 64708 9100 64876 9156
rect 64932 9100 66444 9156
rect 66500 9100 66510 9156
rect 130162 9100 130172 9156
rect 130228 9100 131292 9156
rect 131348 9100 131358 9156
rect 128034 8988 128044 9044
rect 128100 8988 129164 9044
rect 129220 8988 129230 9044
rect 62850 8764 62860 8820
rect 62916 8764 65548 8820
rect 65604 8764 65614 8820
rect 110450 8652 110460 8708
rect 110516 8652 115836 8708
rect 115892 8652 115902 8708
rect 19612 8596 19622 8652
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19886 8596 19896 8652
rect 56432 8596 56442 8652
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56706 8596 56716 8652
rect 93252 8596 93262 8652
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93526 8596 93536 8652
rect 130072 8596 130082 8652
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130346 8596 130356 8652
rect 50306 8428 50316 8484
rect 50372 8428 110460 8484
rect 110516 8428 110526 8484
rect 35074 8316 35084 8372
rect 35140 8316 40572 8372
rect 40628 8316 40638 8372
rect 65762 8316 65772 8372
rect 65828 8316 67676 8372
rect 67732 8316 67742 8372
rect 80770 8316 80780 8372
rect 80836 8316 83132 8372
rect 83188 8316 83198 8372
rect 92530 8316 92540 8372
rect 92596 8316 98252 8372
rect 98308 8316 98318 8372
rect 119186 8204 119196 8260
rect 119252 8204 120540 8260
rect 120596 8204 120606 8260
rect 113586 8092 113596 8148
rect 113652 8092 115164 8148
rect 115220 8092 118300 8148
rect 118356 8092 119420 8148
rect 119476 8092 119486 8148
rect 121426 7980 121436 8036
rect 121492 7980 122444 8036
rect 122500 7980 122510 8036
rect 128930 7980 128940 8036
rect 128996 7980 132300 8036
rect 132356 7980 134764 8036
rect 134820 7980 134830 8036
rect 131282 7868 131292 7924
rect 131348 7868 132860 7924
rect 132916 7868 143836 7924
rect 143892 7868 143902 7924
rect 38022 7812 38032 7868
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38296 7812 38306 7868
rect 74842 7812 74852 7868
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 75116 7812 75126 7868
rect 111662 7812 111672 7868
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111936 7812 111946 7868
rect 148482 7812 148492 7868
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148756 7812 148766 7868
rect 125972 7756 128156 7812
rect 128212 7756 145964 7812
rect 146020 7756 146030 7812
rect 125972 7700 126028 7756
rect 18498 7644 18508 7700
rect 18564 7644 19964 7700
rect 20020 7644 20030 7700
rect 31490 7644 31500 7700
rect 31556 7644 33404 7700
rect 33460 7644 33470 7700
rect 90850 7644 90860 7700
rect 90916 7644 94332 7700
rect 94388 7644 94398 7700
rect 101714 7644 101724 7700
rect 101780 7644 126028 7700
rect 128034 7644 128044 7700
rect 128100 7644 131628 7700
rect 131684 7644 131694 7700
rect 128044 7588 128100 7644
rect 15138 7532 15148 7588
rect 15204 7532 19068 7588
rect 19124 7532 19134 7588
rect 31892 7532 50316 7588
rect 50372 7532 50382 7588
rect 81778 7532 81788 7588
rect 81844 7532 97244 7588
rect 97300 7532 97310 7588
rect 126018 7532 126028 7588
rect 126084 7532 128100 7588
rect 129714 7532 129724 7588
rect 129780 7532 133644 7588
rect 133700 7532 133710 7588
rect 31892 7476 31948 7532
rect 14914 7420 14924 7476
rect 14980 7420 31948 7476
rect 47842 7420 47852 7476
rect 47908 7420 48748 7476
rect 48804 7420 48814 7476
rect 50082 7420 50092 7476
rect 50148 7420 51548 7476
rect 51604 7420 51614 7476
rect 63858 7420 63868 7476
rect 63924 7420 65548 7476
rect 65604 7420 65614 7476
rect 76962 7420 76972 7476
rect 77028 7420 78316 7476
rect 78372 7420 78382 7476
rect 89730 7420 89740 7476
rect 89796 7420 90860 7476
rect 90916 7420 90926 7476
rect 119410 7420 119420 7476
rect 119476 7420 121436 7476
rect 121492 7420 121502 7476
rect 121986 7420 121996 7476
rect 122052 7420 123340 7476
rect 123396 7420 123406 7476
rect 127026 7420 127036 7476
rect 127092 7420 128156 7476
rect 128212 7420 130844 7476
rect 130900 7420 142492 7476
rect 142548 7420 142558 7476
rect 27122 7308 27132 7364
rect 27188 7308 29148 7364
rect 29204 7308 29214 7364
rect 37874 7308 37884 7364
rect 37940 7308 39228 7364
rect 39284 7308 39294 7364
rect 74610 7308 74620 7364
rect 74676 7308 75068 7364
rect 75124 7308 89068 7364
rect 89124 7308 91420 7364
rect 91476 7308 92876 7364
rect 92932 7308 92942 7364
rect 100258 7308 100268 7364
rect 100324 7308 117516 7364
rect 117572 7308 119644 7364
rect 119700 7308 121212 7364
rect 121268 7308 122892 7364
rect 122948 7308 122958 7364
rect 129602 7308 129612 7364
rect 129668 7308 133532 7364
rect 133588 7308 142380 7364
rect 142436 7308 142446 7364
rect 16594 7196 16604 7252
rect 16660 7196 18172 7252
rect 18228 7196 18238 7252
rect 20402 7196 20412 7252
rect 20468 7196 20748 7252
rect 20804 7196 49756 7252
rect 49812 7196 50540 7252
rect 50596 7196 51100 7252
rect 51156 7196 51166 7252
rect 65874 7196 65884 7252
rect 65940 7196 66444 7252
rect 66500 7196 67228 7252
rect 67284 7196 67294 7252
rect 74050 7196 74060 7252
rect 74116 7196 75180 7252
rect 75236 7196 76748 7252
rect 76804 7196 77868 7252
rect 77924 7196 87612 7252
rect 87668 7196 89180 7252
rect 89236 7196 89628 7252
rect 89684 7196 89694 7252
rect 125972 7196 128940 7252
rect 128996 7196 143164 7252
rect 143220 7196 143230 7252
rect 125972 7140 126028 7196
rect 105746 7084 105756 7140
rect 105812 7084 126028 7140
rect 132066 7084 132076 7140
rect 132132 7084 133084 7140
rect 133140 7084 143612 7140
rect 143668 7084 143678 7140
rect 19612 7028 19622 7084
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19886 7028 19896 7084
rect 56432 7028 56442 7084
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56706 7028 56716 7084
rect 93252 7028 93262 7084
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93526 7028 93536 7084
rect 130072 7028 130082 7084
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130346 7028 130356 7084
rect 30034 6860 30044 6916
rect 30100 6860 31612 6916
rect 31668 6860 31678 6916
rect 68114 6860 68124 6916
rect 68180 6860 69468 6916
rect 69524 6860 69534 6916
rect 90402 6860 90412 6916
rect 90468 6860 91196 6916
rect 91252 6860 91262 6916
rect 99474 6860 99484 6916
rect 99540 6860 101052 6916
rect 101108 6860 101118 6916
rect 102452 6860 116508 6916
rect 116564 6860 121324 6916
rect 121380 6860 121390 6916
rect 142258 6860 142268 6916
rect 142324 6860 143948 6916
rect 144004 6860 144014 6916
rect 102452 6804 102508 6860
rect 11666 6748 11676 6804
rect 11732 6748 18620 6804
rect 18676 6748 18686 6804
rect 19058 6748 19068 6804
rect 19124 6748 20748 6804
rect 20804 6748 20814 6804
rect 26338 6748 26348 6804
rect 26404 6748 26414 6804
rect 39106 6748 39116 6804
rect 39172 6748 40124 6804
rect 40180 6748 40190 6804
rect 67330 6748 67340 6804
rect 67396 6748 67406 6804
rect 97122 6748 97132 6804
rect 97188 6748 102508 6804
rect 114370 6748 114380 6804
rect 114436 6748 115724 6804
rect 115780 6748 115790 6804
rect 131618 6748 131628 6804
rect 131684 6748 139916 6804
rect 139972 6748 139982 6804
rect 26348 6692 26404 6748
rect 67340 6692 67396 6748
rect 18946 6636 18956 6692
rect 19012 6636 20300 6692
rect 20356 6636 20860 6692
rect 20916 6636 27860 6692
rect 48290 6636 48300 6692
rect 48356 6636 49532 6692
rect 49588 6636 49598 6692
rect 64642 6636 64652 6692
rect 64708 6636 68236 6692
rect 68292 6636 68302 6692
rect 91970 6636 91980 6692
rect 92036 6636 93100 6692
rect 93156 6636 98476 6692
rect 98532 6636 100268 6692
rect 100324 6636 100334 6692
rect 113026 6636 113036 6692
rect 113092 6636 116732 6692
rect 116788 6636 116798 6692
rect 27804 6580 27860 6636
rect 10882 6524 10892 6580
rect 10948 6524 13580 6580
rect 13636 6524 20412 6580
rect 20468 6524 20478 6580
rect 27794 6524 27804 6580
rect 27860 6524 28812 6580
rect 28868 6524 30268 6580
rect 30324 6524 30334 6580
rect 37426 6524 37436 6580
rect 37492 6524 38332 6580
rect 38388 6524 38398 6580
rect 50530 6524 50540 6580
rect 50596 6524 52108 6580
rect 52164 6524 52174 6580
rect 64082 6524 64092 6580
rect 64148 6524 66332 6580
rect 66388 6524 66398 6580
rect 67554 6524 67564 6580
rect 67620 6524 69132 6580
rect 69188 6524 69198 6580
rect 72594 6524 72604 6580
rect 72660 6524 73276 6580
rect 73332 6524 73342 6580
rect 75730 6524 75740 6580
rect 75796 6524 77644 6580
rect 77700 6524 77710 6580
rect 81106 6524 81116 6580
rect 81172 6524 81564 6580
rect 81620 6524 88172 6580
rect 88228 6524 88956 6580
rect 89012 6524 89022 6580
rect 90692 6524 91868 6580
rect 91924 6524 93660 6580
rect 93716 6524 93726 6580
rect 110338 6524 110348 6580
rect 110404 6524 111580 6580
rect 111636 6524 113484 6580
rect 113540 6524 113550 6580
rect 115042 6524 115052 6580
rect 115108 6524 115724 6580
rect 115780 6524 116284 6580
rect 116340 6524 116350 6580
rect 130946 6524 130956 6580
rect 131012 6524 131964 6580
rect 132020 6524 132030 6580
rect 141250 6524 141260 6580
rect 141316 6524 142716 6580
rect 142772 6524 142782 6580
rect 90692 6468 90748 6524
rect 7410 6412 7420 6468
rect 7476 6412 11228 6468
rect 11284 6412 12908 6468
rect 12964 6412 16156 6468
rect 16212 6412 16828 6468
rect 16884 6412 21532 6468
rect 21588 6412 21598 6468
rect 38882 6412 38892 6468
rect 38948 6412 39788 6468
rect 39844 6412 40460 6468
rect 40516 6412 48076 6468
rect 48132 6412 48142 6468
rect 50306 6412 50316 6468
rect 50372 6412 51548 6468
rect 51604 6412 60844 6468
rect 60900 6412 60910 6468
rect 65314 6412 65324 6468
rect 65380 6412 69356 6468
rect 69412 6412 69422 6468
rect 76066 6412 76076 6468
rect 76132 6412 77308 6468
rect 77364 6412 77374 6468
rect 78530 6412 78540 6468
rect 78596 6412 79324 6468
rect 79380 6412 79390 6468
rect 85586 6412 85596 6468
rect 85652 6412 90748 6468
rect 119858 6412 119868 6468
rect 119924 6412 121324 6468
rect 121380 6412 125020 6468
rect 125076 6412 125086 6468
rect 126914 6412 126924 6468
rect 126980 6412 127372 6468
rect 127428 6412 128044 6468
rect 128100 6412 129164 6468
rect 129220 6412 131852 6468
rect 131908 6412 132636 6468
rect 132692 6412 134204 6468
rect 134260 6412 134270 6468
rect 142482 6412 142492 6468
rect 142548 6412 143500 6468
rect 143556 6412 143566 6468
rect 59938 6300 59948 6356
rect 60004 6300 60396 6356
rect 60452 6300 67564 6356
rect 67620 6300 67630 6356
rect 116274 6300 116284 6356
rect 116340 6300 126476 6356
rect 126532 6300 127148 6356
rect 127204 6300 127214 6356
rect 131506 6300 131516 6356
rect 131572 6300 146524 6356
rect 146580 6300 146590 6356
rect 38022 6244 38032 6300
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38296 6244 38306 6300
rect 74842 6244 74852 6300
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 75116 6244 75126 6300
rect 111662 6244 111672 6300
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111936 6244 111946 6300
rect 148482 6244 148492 6300
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148756 6244 148766 6300
rect 65548 6188 72436 6244
rect 114146 6188 114156 6244
rect 114212 6188 132860 6244
rect 132916 6188 132926 6244
rect 65548 6132 65604 6188
rect 72380 6132 72436 6188
rect 16034 6076 16044 6132
rect 16100 6076 16716 6132
rect 16772 6076 16782 6132
rect 17826 6076 17836 6132
rect 17892 6076 18956 6132
rect 19012 6076 19022 6132
rect 19170 6076 19180 6132
rect 19236 6076 20524 6132
rect 20580 6076 20590 6132
rect 49746 6076 49756 6132
rect 49812 6076 51100 6132
rect 51156 6076 51166 6132
rect 60834 6076 60844 6132
rect 60900 6076 65548 6132
rect 65604 6076 65614 6132
rect 68674 6076 68684 6132
rect 68740 6076 72156 6132
rect 72212 6076 72222 6132
rect 72380 6076 87388 6132
rect 87444 6076 88508 6132
rect 88564 6076 90076 6132
rect 90132 6076 90412 6132
rect 90468 6076 90478 6132
rect 107202 6076 107212 6132
rect 107268 6076 107884 6132
rect 107940 6076 108892 6132
rect 108948 6076 108958 6132
rect 110450 6076 110460 6132
rect 110516 6076 111020 6132
rect 111076 6076 126028 6132
rect 132066 6076 132076 6132
rect 132132 6076 132972 6132
rect 133028 6076 133038 6132
rect 139346 6076 139356 6132
rect 139412 6076 140252 6132
rect 140308 6076 140318 6132
rect 142594 6076 142604 6132
rect 142660 6076 143724 6132
rect 143780 6076 143790 6132
rect 145282 6076 145292 6132
rect 145348 6076 147980 6132
rect 148036 6076 148046 6132
rect 18722 5964 18732 6020
rect 18788 5964 21308 6020
rect 21364 5964 21980 6020
rect 22036 5964 22046 6020
rect 36754 5964 36764 6020
rect 36820 5964 37436 6020
rect 37492 5964 37502 6020
rect 39666 5964 39676 6020
rect 39732 5964 40460 6020
rect 40516 5964 40526 6020
rect 46946 5964 46956 6020
rect 47012 5964 47516 6020
rect 47572 5964 47582 6020
rect 66658 5964 66668 6020
rect 66724 5964 67340 6020
rect 67396 5964 67406 6020
rect 70130 5964 70140 6020
rect 70196 5964 71148 6020
rect 71204 5964 71214 6020
rect 72930 5964 72940 6020
rect 72996 5964 74732 6020
rect 74788 5964 74798 6020
rect 91858 5964 91868 6020
rect 91924 5964 95564 6020
rect 95620 5964 95630 6020
rect 112018 5964 112028 6020
rect 112084 5964 114044 6020
rect 114100 5964 114110 6020
rect 114370 5964 114380 6020
rect 114436 5964 115612 6020
rect 115668 5964 115678 6020
rect 125972 5908 126028 6076
rect 132178 5964 132188 6020
rect 132244 5964 133084 6020
rect 133140 5964 134092 6020
rect 134148 5964 134158 6020
rect 137890 5964 137900 6020
rect 137956 5964 138684 6020
rect 138740 5964 138750 6020
rect 143378 5964 143388 6020
rect 143444 5964 144844 6020
rect 144900 5964 144910 6020
rect 15810 5852 15820 5908
rect 15876 5852 18396 5908
rect 18452 5852 18462 5908
rect 28018 5852 28028 5908
rect 28084 5852 31836 5908
rect 31892 5852 41020 5908
rect 41076 5852 41468 5908
rect 41524 5852 43708 5908
rect 48738 5852 48748 5908
rect 48804 5852 49084 5908
rect 49140 5852 49420 5908
rect 49476 5852 49486 5908
rect 52882 5852 52892 5908
rect 52948 5852 53340 5908
rect 53396 5852 55468 5908
rect 66098 5852 66108 5908
rect 66164 5852 67900 5908
rect 67956 5852 67966 5908
rect 69122 5852 69132 5908
rect 69188 5852 70700 5908
rect 70756 5852 70766 5908
rect 90962 5852 90972 5908
rect 91028 5852 91980 5908
rect 92036 5852 92046 5908
rect 109554 5852 109564 5908
rect 109620 5852 110348 5908
rect 110404 5852 110414 5908
rect 119634 5852 119644 5908
rect 119700 5852 121772 5908
rect 121828 5852 121838 5908
rect 125972 5852 140812 5908
rect 140868 5852 141372 5908
rect 141428 5852 142268 5908
rect 142324 5852 142334 5908
rect 43652 5796 43708 5852
rect 55412 5796 55468 5852
rect 20626 5740 20636 5796
rect 20692 5740 21196 5796
rect 21252 5740 21262 5796
rect 24546 5740 24556 5796
rect 24612 5740 25788 5796
rect 25844 5740 25854 5796
rect 26898 5740 26908 5796
rect 26964 5740 27916 5796
rect 27972 5740 27982 5796
rect 40226 5740 40236 5796
rect 40292 5740 40908 5796
rect 40964 5740 40974 5796
rect 43652 5740 52556 5796
rect 52612 5740 52622 5796
rect 55412 5740 64876 5796
rect 64932 5740 64942 5796
rect 67106 5740 67116 5796
rect 67172 5740 68684 5796
rect 68740 5740 68750 5796
rect 108210 5740 108220 5796
rect 108276 5740 116172 5796
rect 116228 5740 119980 5796
rect 120036 5740 120046 5796
rect 134306 5740 134316 5796
rect 134372 5740 134988 5796
rect 135044 5740 141260 5796
rect 141316 5740 141326 5796
rect 141922 5740 141932 5796
rect 141988 5740 142492 5796
rect 142548 5740 142558 5796
rect 141932 5684 141988 5740
rect 36754 5628 36764 5684
rect 36820 5628 37548 5684
rect 37604 5628 37614 5684
rect 38210 5628 38220 5684
rect 38276 5628 40348 5684
rect 40404 5628 40414 5684
rect 66658 5628 66668 5684
rect 66724 5628 67788 5684
rect 67844 5628 67854 5684
rect 70466 5628 70476 5684
rect 70532 5628 76300 5684
rect 76356 5628 76366 5684
rect 111010 5628 111020 5684
rect 111076 5628 113932 5684
rect 113988 5628 113998 5684
rect 131842 5628 131852 5684
rect 131908 5628 133980 5684
rect 134036 5628 134046 5684
rect 137330 5628 137340 5684
rect 137396 5628 139692 5684
rect 139748 5628 139758 5684
rect 141362 5628 141372 5684
rect 141428 5628 141988 5684
rect 66770 5516 66780 5572
rect 66836 5516 68460 5572
rect 68516 5516 68526 5572
rect 110338 5516 110348 5572
rect 110404 5516 111132 5572
rect 111188 5516 126028 5572
rect 19612 5460 19622 5516
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19886 5460 19896 5516
rect 56432 5460 56442 5516
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56706 5460 56716 5516
rect 93252 5460 93262 5516
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93526 5460 93536 5516
rect 44594 5404 44604 5460
rect 44660 5404 48412 5460
rect 48468 5404 48860 5460
rect 48916 5404 48926 5460
rect 125972 5348 126028 5516
rect 130072 5460 130082 5516
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130346 5460 130356 5516
rect 132850 5404 132860 5460
rect 132916 5404 138908 5460
rect 138964 5404 139692 5460
rect 139748 5404 139758 5460
rect 27906 5292 27916 5348
rect 27972 5292 28700 5348
rect 28756 5292 28766 5348
rect 30930 5292 30940 5348
rect 30996 5292 31948 5348
rect 32004 5292 32014 5348
rect 48636 5292 53564 5348
rect 53620 5292 54124 5348
rect 54180 5292 54190 5348
rect 72370 5292 72380 5348
rect 72436 5292 72940 5348
rect 72996 5292 73006 5348
rect 93650 5292 93660 5348
rect 93716 5292 98700 5348
rect 98756 5292 98766 5348
rect 102452 5292 115948 5348
rect 116004 5292 116172 5348
rect 116228 5292 119868 5348
rect 119924 5292 120988 5348
rect 121044 5292 121054 5348
rect 125972 5292 128492 5348
rect 128548 5292 137900 5348
rect 137956 5292 137966 5348
rect 12674 5180 12684 5236
rect 12740 5180 13580 5236
rect 13636 5180 13646 5236
rect 21186 5180 21196 5236
rect 21252 5180 21756 5236
rect 21812 5180 22204 5236
rect 22260 5180 28252 5236
rect 28308 5180 28318 5236
rect 40898 5180 40908 5236
rect 40964 5180 41692 5236
rect 41748 5180 42308 5236
rect 42252 5124 42308 5180
rect 48636 5124 48692 5292
rect 102452 5236 102508 5292
rect 52546 5180 52556 5236
rect 52612 5180 54460 5236
rect 54516 5180 60620 5236
rect 60676 5180 62300 5236
rect 62356 5180 67004 5236
rect 67060 5180 67070 5236
rect 76300 5180 77308 5236
rect 77364 5180 77374 5236
rect 88386 5180 88396 5236
rect 88452 5180 89404 5236
rect 89460 5180 89470 5236
rect 90738 5180 90748 5236
rect 90804 5180 91644 5236
rect 91700 5180 92204 5236
rect 92260 5180 93100 5236
rect 93156 5180 93166 5236
rect 94546 5180 94556 5236
rect 94612 5180 97804 5236
rect 97860 5180 98364 5236
rect 98420 5180 101948 5236
rect 102004 5180 102508 5236
rect 102564 5180 102574 5236
rect 107538 5180 107548 5236
rect 107604 5180 108220 5236
rect 108276 5180 108286 5236
rect 115042 5180 115052 5236
rect 115108 5180 116732 5236
rect 116788 5180 121100 5236
rect 121156 5180 121166 5236
rect 136210 5180 136220 5236
rect 136276 5180 138012 5236
rect 138068 5180 138078 5236
rect 138338 5180 138348 5236
rect 138404 5180 140140 5236
rect 140196 5180 140206 5236
rect 144498 5180 144508 5236
rect 144564 5180 145852 5236
rect 145908 5180 147868 5236
rect 147924 5180 147934 5236
rect 76300 5124 76356 5180
rect 107548 5124 107604 5180
rect 10210 5068 10220 5124
rect 10276 5068 11676 5124
rect 11732 5068 11742 5124
rect 21522 5068 21532 5124
rect 21588 5068 25116 5124
rect 25172 5068 29484 5124
rect 29540 5068 35532 5124
rect 35588 5068 35598 5124
rect 38546 5068 38556 5124
rect 38612 5068 41580 5124
rect 41636 5068 41646 5124
rect 42242 5068 42252 5124
rect 42308 5068 48076 5124
rect 48132 5068 48636 5124
rect 48692 5068 48702 5124
rect 49858 5068 49868 5124
rect 49924 5068 53452 5124
rect 53508 5068 53518 5124
rect 54114 5068 54124 5124
rect 54180 5068 57820 5124
rect 57876 5068 57886 5124
rect 61730 5068 61740 5124
rect 61796 5068 62524 5124
rect 62580 5068 62590 5124
rect 67554 5068 67564 5124
rect 67620 5068 69468 5124
rect 69524 5068 69534 5124
rect 72482 5068 72492 5124
rect 72548 5068 75628 5124
rect 75684 5068 76300 5124
rect 76356 5068 76366 5124
rect 76626 5068 76636 5124
rect 76692 5068 80444 5124
rect 80500 5068 84476 5124
rect 84532 5068 85484 5124
rect 85540 5068 94892 5124
rect 94948 5068 95228 5124
rect 95284 5068 107604 5124
rect 107874 5068 107884 5124
rect 107940 5068 109228 5124
rect 109284 5068 109294 5124
rect 117170 5068 117180 5124
rect 117236 5068 126924 5124
rect 126980 5068 126990 5124
rect 130946 5068 130956 5124
rect 131012 5068 131964 5124
rect 132020 5068 132030 5124
rect 134194 5068 134204 5124
rect 134260 5068 136332 5124
rect 136388 5068 136398 5124
rect 11778 4956 11788 5012
rect 11844 4956 12236 5012
rect 12292 4956 12460 5012
rect 12516 4956 15820 5012
rect 15876 4956 16492 5012
rect 16548 4956 16558 5012
rect 44706 4956 44716 5012
rect 44772 4956 45276 5012
rect 45332 4956 45612 5012
rect 45668 4956 45678 5012
rect 52994 4956 53004 5012
rect 53060 4956 55692 5012
rect 55748 4956 55758 5012
rect 62178 4956 62188 5012
rect 62244 4956 63196 5012
rect 63252 4956 63262 5012
rect 67172 4956 71484 5012
rect 71540 4956 71932 5012
rect 71988 4956 82068 5012
rect 82226 4956 82236 5012
rect 82292 4956 86268 5012
rect 86324 4956 86334 5012
rect 90692 4956 91084 5012
rect 91140 4956 92428 5012
rect 92484 4956 93660 5012
rect 93716 4956 94220 5012
rect 94276 4956 94286 5012
rect 109666 4956 109676 5012
rect 109732 4956 110684 5012
rect 110740 4956 110750 5012
rect 133298 4956 133308 5012
rect 133364 4956 134540 5012
rect 134596 4956 135212 5012
rect 135268 4956 135278 5012
rect 139122 4956 139132 5012
rect 139188 4956 142716 5012
rect 142772 4956 145180 5012
rect 145236 4956 145246 5012
rect 67172 4900 67228 4956
rect 82012 4900 82068 4956
rect 90692 4900 90748 4956
rect 11106 4844 11116 4900
rect 11172 4844 17948 4900
rect 18004 4844 18014 4900
rect 20290 4844 20300 4900
rect 20356 4844 21644 4900
rect 21700 4844 21710 4900
rect 26002 4844 26012 4900
rect 26068 4844 31388 4900
rect 31444 4844 31454 4900
rect 56802 4844 56812 4900
rect 56868 4844 57260 4900
rect 57316 4844 58156 4900
rect 58212 4844 67228 4900
rect 69346 4844 69356 4900
rect 69412 4844 71148 4900
rect 71204 4844 71214 4900
rect 73714 4844 73724 4900
rect 73780 4844 80220 4900
rect 80276 4844 80286 4900
rect 82012 4844 90748 4900
rect 111346 4844 111356 4900
rect 111412 4844 113596 4900
rect 113652 4844 113662 4900
rect 115826 4844 115836 4900
rect 115892 4844 117180 4900
rect 117236 4844 117246 4900
rect 128594 4844 128604 4900
rect 128660 4844 137004 4900
rect 137060 4844 137070 4900
rect 139010 4844 139020 4900
rect 139076 4844 141708 4900
rect 141764 4844 142604 4900
rect 142660 4844 142670 4900
rect 143154 4844 143164 4900
rect 143220 4844 143500 4900
rect 143556 4844 145068 4900
rect 145124 4844 145134 4900
rect 38022 4676 38032 4732
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38296 4676 38306 4732
rect 74842 4676 74852 4732
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 75116 4676 75126 4732
rect 111662 4676 111672 4732
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111936 4676 111946 4732
rect 148482 4676 148492 4732
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148756 4676 148766 4732
rect 80434 4620 80444 4676
rect 80500 4620 81228 4676
rect 81284 4620 81676 4676
rect 81732 4620 89516 4676
rect 89572 4620 90748 4676
rect 90804 4620 90814 4676
rect 8306 4508 8316 4564
rect 8372 4508 10108 4564
rect 10164 4508 10174 4564
rect 10322 4508 10332 4564
rect 10388 4508 12012 4564
rect 12068 4508 12078 4564
rect 38434 4508 38444 4564
rect 38500 4508 39116 4564
rect 39172 4508 39564 4564
rect 39620 4508 39630 4564
rect 55010 4508 55020 4564
rect 55076 4508 56476 4564
rect 56532 4508 65884 4564
rect 65940 4508 65950 4564
rect 100034 4508 100044 4564
rect 100100 4508 100110 4564
rect 102050 4508 102060 4564
rect 102116 4508 102508 4564
rect 102564 4508 102574 4564
rect 119970 4508 119980 4564
rect 120036 4508 124236 4564
rect 124292 4508 124684 4564
rect 124740 4508 127372 4564
rect 127428 4508 127438 4564
rect 132178 4508 132188 4564
rect 132244 4508 133756 4564
rect 133812 4508 134876 4564
rect 134932 4508 134942 4564
rect 145954 4508 145964 4564
rect 146020 4508 146748 4564
rect 146804 4508 146814 4564
rect 100044 4452 100100 4508
rect 6850 4396 6860 4452
rect 6916 4396 7420 4452
rect 7476 4396 7486 4452
rect 9762 4396 9772 4452
rect 9828 4396 11004 4452
rect 11060 4396 11070 4452
rect 20514 4396 20524 4452
rect 20580 4396 21084 4452
rect 21140 4396 21150 4452
rect 27458 4396 27468 4452
rect 27524 4396 28924 4452
rect 28980 4396 28990 4452
rect 31266 4396 31276 4452
rect 31332 4396 32732 4452
rect 32788 4396 33516 4452
rect 33572 4396 33582 4452
rect 56802 4396 56812 4452
rect 56868 4396 57596 4452
rect 57652 4396 57662 4452
rect 86818 4396 86828 4452
rect 86884 4396 88508 4452
rect 88564 4396 101612 4452
rect 101668 4396 103180 4452
rect 103236 4396 103246 4452
rect 132626 4396 132636 4452
rect 132692 4396 137340 4452
rect 137396 4396 137406 4452
rect 137732 4396 141484 4452
rect 141540 4396 141550 4452
rect 145170 4396 145180 4452
rect 145236 4396 145628 4452
rect 145684 4396 145694 4452
rect 137732 4340 137788 4396
rect 40226 4284 40236 4340
rect 40292 4284 45276 4340
rect 45332 4284 45342 4340
rect 66658 4284 66668 4340
rect 66724 4284 68572 4340
rect 68628 4284 69244 4340
rect 69300 4284 72492 4340
rect 72548 4284 72558 4340
rect 86258 4284 86268 4340
rect 86324 4284 89180 4340
rect 89236 4284 99036 4340
rect 99092 4284 99484 4340
rect 99540 4284 112028 4340
rect 112084 4284 113036 4340
rect 113092 4284 113102 4340
rect 125346 4284 125356 4340
rect 125412 4284 128604 4340
rect 128660 4284 128670 4340
rect 129602 4284 129612 4340
rect 129668 4284 136892 4340
rect 136948 4284 137788 4340
rect 6626 4172 6636 4228
rect 6692 4172 8764 4228
rect 8820 4172 10220 4228
rect 10276 4172 10286 4228
rect 27570 4172 27580 4228
rect 27636 4172 29820 4228
rect 29876 4172 29886 4228
rect 30706 4172 30716 4228
rect 30772 4172 32060 4228
rect 32116 4172 32126 4228
rect 39330 4172 39340 4228
rect 39396 4172 40348 4228
rect 40404 4172 40414 4228
rect 45042 4172 45052 4228
rect 45108 4172 50764 4228
rect 50820 4172 50830 4228
rect 91746 4172 91756 4228
rect 91812 4172 93436 4228
rect 93492 4172 93502 4228
rect 110674 4172 110684 4228
rect 110740 4172 111692 4228
rect 111748 4172 114268 4228
rect 115938 4172 115948 4228
rect 116004 4172 117292 4228
rect 117348 4172 117358 4228
rect 132066 4172 132076 4228
rect 132132 4172 133196 4228
rect 133252 4172 133262 4228
rect 145618 4172 145628 4228
rect 145684 4172 147196 4228
rect 147252 4172 147262 4228
rect 30716 4116 30772 4172
rect 114212 4116 114268 4172
rect 28242 4060 28252 4116
rect 28308 4060 29260 4116
rect 29316 4060 30772 4116
rect 78932 4060 108332 4116
rect 108388 4060 112588 4116
rect 112644 4060 112654 4116
rect 114212 4060 118188 4116
rect 118244 4060 120428 4116
rect 120484 4060 120494 4116
rect 125972 4060 132468 4116
rect 132626 4060 132636 4116
rect 132692 4060 134316 4116
rect 134372 4060 134382 4116
rect 78932 4004 78988 4060
rect 5842 3948 5852 4004
rect 5908 3948 6412 4004
rect 6468 3948 13916 4004
rect 13972 3948 14364 4004
rect 14420 3948 16604 4004
rect 16660 3948 16670 4004
rect 57026 3948 57036 4004
rect 57092 3948 58828 4004
rect 58884 3948 59836 4004
rect 59892 3948 78988 4004
rect 19612 3892 19622 3948
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19886 3892 19896 3948
rect 56432 3892 56442 3948
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56706 3892 56716 3948
rect 93252 3892 93262 3948
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93526 3892 93536 3948
rect 61954 3836 61964 3892
rect 62020 3836 67676 3892
rect 67732 3836 81788 3892
rect 81844 3836 81854 3892
rect 94546 3836 94556 3892
rect 94612 3836 95900 3892
rect 95956 3836 120652 3892
rect 120708 3836 120718 3892
rect 125972 3780 126028 4060
rect 132412 4004 132468 4060
rect 132412 3948 133308 4004
rect 133364 3948 133374 4004
rect 130072 3892 130082 3948
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130346 3892 130356 3948
rect 16482 3724 16492 3780
rect 16548 3724 29484 3780
rect 29540 3724 30044 3780
rect 30100 3724 30110 3780
rect 39666 3724 39676 3780
rect 39732 3724 40572 3780
rect 40628 3724 40638 3780
rect 77074 3724 77084 3780
rect 77140 3724 79212 3780
rect 79268 3724 79278 3780
rect 112578 3724 112588 3780
rect 112644 3724 126028 3780
rect 127810 3724 127820 3780
rect 127876 3724 131516 3780
rect 131572 3724 131582 3780
rect 132290 3724 132300 3780
rect 132356 3724 133420 3780
rect 133476 3724 133486 3780
rect 6402 3612 6412 3668
rect 6468 3612 11340 3668
rect 11396 3612 11406 3668
rect 23314 3612 23324 3668
rect 23380 3612 25004 3668
rect 25060 3612 25070 3668
rect 31154 3612 31164 3668
rect 31220 3612 32956 3668
rect 33012 3612 33022 3668
rect 33394 3612 33404 3668
rect 33460 3612 34860 3668
rect 34916 3612 34926 3668
rect 35522 3612 35532 3668
rect 35588 3612 40236 3668
rect 40292 3612 40302 3668
rect 46722 3612 46732 3668
rect 46788 3612 47516 3668
rect 47572 3612 47582 3668
rect 58034 3612 58044 3668
rect 58100 3612 59612 3668
rect 59668 3612 59678 3668
rect 64642 3612 64652 3668
rect 64708 3612 68572 3668
rect 68628 3612 69356 3668
rect 69412 3612 69422 3668
rect 79314 3612 79324 3668
rect 79380 3612 80332 3668
rect 80388 3612 80398 3668
rect 98802 3612 98812 3668
rect 98868 3612 101836 3668
rect 101892 3612 101902 3668
rect 102834 3612 102844 3668
rect 102900 3612 104972 3668
rect 105028 3612 105038 3668
rect 108770 3612 108780 3668
rect 108836 3612 110572 3668
rect 110628 3612 110638 3668
rect 114594 3612 114604 3668
rect 114660 3612 119980 3668
rect 120036 3612 120046 3668
rect 131618 3612 131628 3668
rect 131684 3612 132188 3668
rect 132244 3612 132254 3668
rect 137330 3612 137340 3668
rect 137396 3612 139020 3668
rect 139076 3612 139086 3668
rect 140130 3612 140140 3668
rect 140196 3612 141036 3668
rect 141092 3612 141102 3668
rect 144162 3612 144172 3668
rect 144228 3612 147532 3668
rect 147588 3612 147598 3668
rect 6290 3500 6300 3556
rect 6356 3500 10164 3556
rect 11106 3500 11116 3556
rect 11172 3500 11900 3556
rect 11956 3500 12348 3556
rect 12404 3500 12414 3556
rect 16268 3500 19404 3556
rect 19460 3500 19470 3556
rect 30034 3500 30044 3556
rect 30100 3500 59388 3556
rect 59444 3500 59454 3556
rect 60834 3500 60844 3556
rect 60900 3500 64876 3556
rect 64932 3500 65212 3556
rect 65268 3500 65278 3556
rect 72594 3500 72604 3556
rect 72660 3500 76972 3556
rect 77028 3500 77308 3556
rect 77364 3500 77374 3556
rect 111794 3500 111804 3556
rect 111860 3500 112364 3556
rect 112420 3500 115668 3556
rect 117282 3500 117292 3556
rect 117348 3500 118524 3556
rect 118580 3500 123228 3556
rect 123284 3500 123294 3556
rect 129378 3500 129388 3556
rect 129444 3500 130284 3556
rect 130340 3500 135660 3556
rect 135716 3500 135726 3556
rect 144050 3500 144060 3556
rect 144116 3500 145068 3556
rect 145124 3500 145134 3556
rect 10108 3444 10164 3500
rect 16268 3444 16324 3500
rect 115612 3444 115668 3500
rect 6850 3388 6860 3444
rect 6916 3388 9884 3444
rect 9940 3388 9950 3444
rect 10098 3388 10108 3444
rect 10164 3388 14476 3444
rect 14532 3388 14542 3444
rect 15138 3388 15148 3444
rect 15204 3388 16268 3444
rect 16324 3388 16334 3444
rect 16482 3388 16492 3444
rect 16548 3388 17612 3444
rect 17668 3388 17678 3444
rect 20514 3388 20524 3444
rect 20580 3388 22204 3444
rect 22260 3388 22270 3444
rect 23202 3388 23212 3444
rect 23268 3388 24108 3444
rect 24164 3388 25228 3444
rect 25284 3388 25294 3444
rect 26562 3388 26572 3444
rect 26628 3388 27244 3444
rect 27300 3388 27310 3444
rect 36194 3388 36204 3444
rect 36260 3388 36876 3444
rect 36932 3388 36942 3444
rect 37762 3388 37772 3444
rect 37828 3388 38332 3444
rect 38388 3388 38398 3444
rect 40674 3388 40684 3444
rect 40740 3388 41244 3444
rect 41300 3388 41692 3444
rect 41748 3388 41758 3444
rect 45266 3388 45276 3444
rect 45332 3388 48860 3444
rect 48916 3388 62188 3444
rect 62244 3388 62254 3444
rect 73826 3388 73836 3444
rect 73892 3388 75628 3444
rect 75684 3388 75694 3444
rect 80994 3388 81004 3444
rect 81060 3388 82908 3444
rect 82964 3388 84028 3444
rect 84084 3388 84094 3444
rect 85026 3388 85036 3444
rect 85092 3388 86828 3444
rect 86884 3388 87948 3444
rect 88004 3388 88014 3444
rect 89058 3388 89068 3444
rect 89124 3388 91084 3444
rect 91140 3388 91868 3444
rect 91924 3388 91934 3444
rect 93090 3388 93100 3444
rect 93156 3388 94668 3444
rect 94724 3388 96236 3444
rect 96292 3388 96302 3444
rect 113250 3388 113260 3444
rect 113316 3388 114604 3444
rect 114660 3388 114670 3444
rect 115602 3388 115612 3444
rect 115668 3388 116284 3444
rect 116340 3388 119420 3444
rect 119476 3388 119486 3444
rect 120082 3388 120092 3444
rect 120148 3388 121772 3444
rect 121828 3388 121838 3444
rect 122098 3388 122108 3444
rect 122164 3388 123676 3444
rect 123732 3388 123742 3444
rect 124002 3388 124012 3444
rect 124068 3388 125692 3444
rect 125748 3388 125758 3444
rect 126018 3388 126028 3444
rect 126084 3388 126364 3444
rect 126420 3388 127148 3444
rect 127204 3388 127214 3444
rect 133298 3388 133308 3444
rect 133364 3388 138012 3444
rect 138068 3388 138078 3444
rect 9884 3332 9940 3388
rect 9884 3276 10332 3332
rect 10388 3276 10398 3332
rect 20132 3276 55916 3332
rect 55972 3276 56700 3332
rect 56756 3276 56766 3332
rect 20132 3220 20188 3276
rect 8866 3164 8876 3220
rect 8932 3164 20188 3220
rect 38022 3108 38032 3164
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38296 3108 38306 3164
rect 74842 3108 74852 3164
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 75116 3108 75126 3164
rect 111662 3108 111672 3164
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111936 3108 111946 3164
rect 148482 3108 148492 3164
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148756 3108 148766 3164
rect 5730 2492 5740 2548
rect 5796 2492 70588 2548
rect 70644 2492 70654 2548
<< via3 >>
rect 19622 36820 19678 36876
rect 19726 36820 19782 36876
rect 19830 36820 19886 36876
rect 56442 36820 56498 36876
rect 56546 36820 56602 36876
rect 56650 36820 56706 36876
rect 93262 36820 93318 36876
rect 93366 36820 93422 36876
rect 93470 36820 93526 36876
rect 130082 36820 130138 36876
rect 130186 36820 130242 36876
rect 130290 36820 130346 36876
rect 75628 36316 75684 36372
rect 38032 36036 38088 36092
rect 38136 36036 38192 36092
rect 38240 36036 38296 36092
rect 74852 36036 74908 36092
rect 74956 36036 75012 36092
rect 75060 36036 75116 36092
rect 111672 36036 111728 36092
rect 111776 36036 111832 36092
rect 111880 36036 111936 36092
rect 148492 36036 148548 36092
rect 148596 36036 148652 36092
rect 148700 36036 148756 36092
rect 91420 35980 91476 36036
rect 82236 35868 82292 35924
rect 91532 35756 91588 35812
rect 77084 35532 77140 35588
rect 19622 35252 19678 35308
rect 19726 35252 19782 35308
rect 19830 35252 19886 35308
rect 56442 35252 56498 35308
rect 56546 35252 56602 35308
rect 56650 35252 56706 35308
rect 93262 35252 93318 35308
rect 93366 35252 93422 35308
rect 93470 35252 93526 35308
rect 130082 35252 130138 35308
rect 130186 35252 130242 35308
rect 130290 35252 130346 35308
rect 75628 35084 75684 35140
rect 38032 34468 38088 34524
rect 38136 34468 38192 34524
rect 38240 34468 38296 34524
rect 115052 34972 115108 35028
rect 115052 34636 115108 34692
rect 74852 34468 74908 34524
rect 74956 34468 75012 34524
rect 75060 34468 75116 34524
rect 111672 34468 111728 34524
rect 111776 34468 111832 34524
rect 111880 34468 111936 34524
rect 82236 34412 82292 34468
rect 77084 34300 77140 34356
rect 148492 34468 148548 34524
rect 148596 34468 148652 34524
rect 148700 34468 148756 34524
rect 43596 33852 43652 33908
rect 19622 33684 19678 33740
rect 19726 33684 19782 33740
rect 19830 33684 19886 33740
rect 56442 33684 56498 33740
rect 56546 33684 56602 33740
rect 56650 33684 56706 33740
rect 93262 33684 93318 33740
rect 93366 33684 93422 33740
rect 93470 33684 93526 33740
rect 130082 33684 130138 33740
rect 130186 33684 130242 33740
rect 130290 33684 130346 33740
rect 43596 33628 43652 33684
rect 38032 32900 38088 32956
rect 38136 32900 38192 32956
rect 38240 32900 38296 32956
rect 58828 32844 58884 32900
rect 74852 32900 74908 32956
rect 74956 32900 75012 32956
rect 75060 32900 75116 32956
rect 111672 32900 111728 32956
rect 111776 32900 111832 32956
rect 111880 32900 111936 32956
rect 148492 32900 148548 32956
rect 148596 32900 148652 32956
rect 148700 32900 148756 32956
rect 19622 32116 19678 32172
rect 19726 32116 19782 32172
rect 19830 32116 19886 32172
rect 56442 32116 56498 32172
rect 56546 32116 56602 32172
rect 56650 32116 56706 32172
rect 93262 32116 93318 32172
rect 93366 32116 93422 32172
rect 93470 32116 93526 32172
rect 130082 32116 130138 32172
rect 130186 32116 130242 32172
rect 130290 32116 130346 32172
rect 105756 31948 105812 32004
rect 105756 31500 105812 31556
rect 38032 31332 38088 31388
rect 38136 31332 38192 31388
rect 38240 31332 38296 31388
rect 74852 31332 74908 31388
rect 74956 31332 75012 31388
rect 75060 31332 75116 31388
rect 111672 31332 111728 31388
rect 111776 31332 111832 31388
rect 111880 31332 111936 31388
rect 148492 31332 148548 31388
rect 148596 31332 148652 31388
rect 148700 31332 148756 31388
rect 19622 30548 19678 30604
rect 19726 30548 19782 30604
rect 19830 30548 19886 30604
rect 56442 30548 56498 30604
rect 56546 30548 56602 30604
rect 56650 30548 56706 30604
rect 93262 30548 93318 30604
rect 93366 30548 93422 30604
rect 93470 30548 93526 30604
rect 130082 30548 130138 30604
rect 130186 30548 130242 30604
rect 130290 30548 130346 30604
rect 38032 29764 38088 29820
rect 38136 29764 38192 29820
rect 38240 29764 38296 29820
rect 74852 29764 74908 29820
rect 74956 29764 75012 29820
rect 75060 29764 75116 29820
rect 111672 29764 111728 29820
rect 111776 29764 111832 29820
rect 111880 29764 111936 29820
rect 148492 29764 148548 29820
rect 148596 29764 148652 29820
rect 148700 29764 148756 29820
rect 19622 28980 19678 29036
rect 19726 28980 19782 29036
rect 19830 28980 19886 29036
rect 56442 28980 56498 29036
rect 56546 28980 56602 29036
rect 56650 28980 56706 29036
rect 93262 28980 93318 29036
rect 93366 28980 93422 29036
rect 93470 28980 93526 29036
rect 130082 28980 130138 29036
rect 130186 28980 130242 29036
rect 130290 28980 130346 29036
rect 38032 28196 38088 28252
rect 38136 28196 38192 28252
rect 38240 28196 38296 28252
rect 74852 28196 74908 28252
rect 74956 28196 75012 28252
rect 75060 28196 75116 28252
rect 111672 28196 111728 28252
rect 111776 28196 111832 28252
rect 111880 28196 111936 28252
rect 148492 28196 148548 28252
rect 148596 28196 148652 28252
rect 148700 28196 148756 28252
rect 19622 27412 19678 27468
rect 19726 27412 19782 27468
rect 19830 27412 19886 27468
rect 56442 27412 56498 27468
rect 56546 27412 56602 27468
rect 56650 27412 56706 27468
rect 93262 27412 93318 27468
rect 93366 27412 93422 27468
rect 93470 27412 93526 27468
rect 130082 27412 130138 27468
rect 130186 27412 130242 27468
rect 130290 27412 130346 27468
rect 38032 26628 38088 26684
rect 38136 26628 38192 26684
rect 38240 26628 38296 26684
rect 74852 26628 74908 26684
rect 74956 26628 75012 26684
rect 75060 26628 75116 26684
rect 111672 26628 111728 26684
rect 111776 26628 111832 26684
rect 111880 26628 111936 26684
rect 148492 26628 148548 26684
rect 148596 26628 148652 26684
rect 148700 26628 148756 26684
rect 19622 25844 19678 25900
rect 19726 25844 19782 25900
rect 19830 25844 19886 25900
rect 56442 25844 56498 25900
rect 56546 25844 56602 25900
rect 56650 25844 56706 25900
rect 93262 25844 93318 25900
rect 93366 25844 93422 25900
rect 93470 25844 93526 25900
rect 130082 25844 130138 25900
rect 130186 25844 130242 25900
rect 130290 25844 130346 25900
rect 58828 25116 58884 25172
rect 38032 25060 38088 25116
rect 38136 25060 38192 25116
rect 38240 25060 38296 25116
rect 74852 25060 74908 25116
rect 74956 25060 75012 25116
rect 75060 25060 75116 25116
rect 111672 25060 111728 25116
rect 111776 25060 111832 25116
rect 111880 25060 111936 25116
rect 148492 25060 148548 25116
rect 148596 25060 148652 25116
rect 148700 25060 148756 25116
rect 19622 24276 19678 24332
rect 19726 24276 19782 24332
rect 19830 24276 19886 24332
rect 56442 24276 56498 24332
rect 56546 24276 56602 24332
rect 56650 24276 56706 24332
rect 93262 24276 93318 24332
rect 93366 24276 93422 24332
rect 93470 24276 93526 24332
rect 130082 24276 130138 24332
rect 130186 24276 130242 24332
rect 130290 24276 130346 24332
rect 38032 23492 38088 23548
rect 38136 23492 38192 23548
rect 38240 23492 38296 23548
rect 74852 23492 74908 23548
rect 74956 23492 75012 23548
rect 75060 23492 75116 23548
rect 111672 23492 111728 23548
rect 111776 23492 111832 23548
rect 111880 23492 111936 23548
rect 148492 23492 148548 23548
rect 148596 23492 148652 23548
rect 148700 23492 148756 23548
rect 19622 22708 19678 22764
rect 19726 22708 19782 22764
rect 19830 22708 19886 22764
rect 56442 22708 56498 22764
rect 56546 22708 56602 22764
rect 56650 22708 56706 22764
rect 93262 22708 93318 22764
rect 93366 22708 93422 22764
rect 93470 22708 93526 22764
rect 130082 22708 130138 22764
rect 130186 22708 130242 22764
rect 130290 22708 130346 22764
rect 38032 21924 38088 21980
rect 38136 21924 38192 21980
rect 38240 21924 38296 21980
rect 74852 21924 74908 21980
rect 74956 21924 75012 21980
rect 75060 21924 75116 21980
rect 111672 21924 111728 21980
rect 111776 21924 111832 21980
rect 111880 21924 111936 21980
rect 148492 21924 148548 21980
rect 148596 21924 148652 21980
rect 148700 21924 148756 21980
rect 19622 21140 19678 21196
rect 19726 21140 19782 21196
rect 19830 21140 19886 21196
rect 56442 21140 56498 21196
rect 56546 21140 56602 21196
rect 56650 21140 56706 21196
rect 93262 21140 93318 21196
rect 93366 21140 93422 21196
rect 93470 21140 93526 21196
rect 130082 21140 130138 21196
rect 130186 21140 130242 21196
rect 130290 21140 130346 21196
rect 38032 20356 38088 20412
rect 38136 20356 38192 20412
rect 38240 20356 38296 20412
rect 74852 20356 74908 20412
rect 74956 20356 75012 20412
rect 75060 20356 75116 20412
rect 111672 20356 111728 20412
rect 111776 20356 111832 20412
rect 111880 20356 111936 20412
rect 148492 20356 148548 20412
rect 148596 20356 148652 20412
rect 148700 20356 148756 20412
rect 19622 19572 19678 19628
rect 19726 19572 19782 19628
rect 19830 19572 19886 19628
rect 56442 19572 56498 19628
rect 56546 19572 56602 19628
rect 56650 19572 56706 19628
rect 93262 19572 93318 19628
rect 93366 19572 93422 19628
rect 93470 19572 93526 19628
rect 130082 19572 130138 19628
rect 130186 19572 130242 19628
rect 130290 19572 130346 19628
rect 38032 18788 38088 18844
rect 38136 18788 38192 18844
rect 38240 18788 38296 18844
rect 74852 18788 74908 18844
rect 74956 18788 75012 18844
rect 75060 18788 75116 18844
rect 111672 18788 111728 18844
rect 111776 18788 111832 18844
rect 111880 18788 111936 18844
rect 148492 18788 148548 18844
rect 148596 18788 148652 18844
rect 148700 18788 148756 18844
rect 19622 18004 19678 18060
rect 19726 18004 19782 18060
rect 19830 18004 19886 18060
rect 56442 18004 56498 18060
rect 56546 18004 56602 18060
rect 56650 18004 56706 18060
rect 93262 18004 93318 18060
rect 93366 18004 93422 18060
rect 93470 18004 93526 18060
rect 130082 18004 130138 18060
rect 130186 18004 130242 18060
rect 130290 18004 130346 18060
rect 38032 17220 38088 17276
rect 38136 17220 38192 17276
rect 38240 17220 38296 17276
rect 74852 17220 74908 17276
rect 74956 17220 75012 17276
rect 75060 17220 75116 17276
rect 111672 17220 111728 17276
rect 111776 17220 111832 17276
rect 111880 17220 111936 17276
rect 148492 17220 148548 17276
rect 148596 17220 148652 17276
rect 148700 17220 148756 17276
rect 19622 16436 19678 16492
rect 19726 16436 19782 16492
rect 19830 16436 19886 16492
rect 56442 16436 56498 16492
rect 56546 16436 56602 16492
rect 56650 16436 56706 16492
rect 93262 16436 93318 16492
rect 93366 16436 93422 16492
rect 93470 16436 93526 16492
rect 130082 16436 130138 16492
rect 130186 16436 130242 16492
rect 130290 16436 130346 16492
rect 38032 15652 38088 15708
rect 38136 15652 38192 15708
rect 38240 15652 38296 15708
rect 74852 15652 74908 15708
rect 74956 15652 75012 15708
rect 75060 15652 75116 15708
rect 111672 15652 111728 15708
rect 111776 15652 111832 15708
rect 111880 15652 111936 15708
rect 148492 15652 148548 15708
rect 148596 15652 148652 15708
rect 148700 15652 148756 15708
rect 19622 14868 19678 14924
rect 19726 14868 19782 14924
rect 19830 14868 19886 14924
rect 56442 14868 56498 14924
rect 56546 14868 56602 14924
rect 56650 14868 56706 14924
rect 93262 14868 93318 14924
rect 93366 14868 93422 14924
rect 93470 14868 93526 14924
rect 130082 14868 130138 14924
rect 130186 14868 130242 14924
rect 130290 14868 130346 14924
rect 38032 14084 38088 14140
rect 38136 14084 38192 14140
rect 38240 14084 38296 14140
rect 74852 14084 74908 14140
rect 74956 14084 75012 14140
rect 75060 14084 75116 14140
rect 111672 14084 111728 14140
rect 111776 14084 111832 14140
rect 111880 14084 111936 14140
rect 148492 14084 148548 14140
rect 148596 14084 148652 14140
rect 148700 14084 148756 14140
rect 19622 13300 19678 13356
rect 19726 13300 19782 13356
rect 19830 13300 19886 13356
rect 56442 13300 56498 13356
rect 56546 13300 56602 13356
rect 56650 13300 56706 13356
rect 93262 13300 93318 13356
rect 93366 13300 93422 13356
rect 93470 13300 93526 13356
rect 130082 13300 130138 13356
rect 130186 13300 130242 13356
rect 130290 13300 130346 13356
rect 38032 12516 38088 12572
rect 38136 12516 38192 12572
rect 38240 12516 38296 12572
rect 74852 12516 74908 12572
rect 74956 12516 75012 12572
rect 75060 12516 75116 12572
rect 111672 12516 111728 12572
rect 111776 12516 111832 12572
rect 111880 12516 111936 12572
rect 148492 12516 148548 12572
rect 148596 12516 148652 12572
rect 148700 12516 148756 12572
rect 19622 11732 19678 11788
rect 19726 11732 19782 11788
rect 19830 11732 19886 11788
rect 56442 11732 56498 11788
rect 56546 11732 56602 11788
rect 56650 11732 56706 11788
rect 93262 11732 93318 11788
rect 93366 11732 93422 11788
rect 93470 11732 93526 11788
rect 130082 11732 130138 11788
rect 130186 11732 130242 11788
rect 130290 11732 130346 11788
rect 38032 10948 38088 11004
rect 38136 10948 38192 11004
rect 38240 10948 38296 11004
rect 74852 10948 74908 11004
rect 74956 10948 75012 11004
rect 75060 10948 75116 11004
rect 111672 10948 111728 11004
rect 111776 10948 111832 11004
rect 111880 10948 111936 11004
rect 148492 10948 148548 11004
rect 148596 10948 148652 11004
rect 148700 10948 148756 11004
rect 19622 10164 19678 10220
rect 19726 10164 19782 10220
rect 19830 10164 19886 10220
rect 56442 10164 56498 10220
rect 56546 10164 56602 10220
rect 56650 10164 56706 10220
rect 93262 10164 93318 10220
rect 93366 10164 93422 10220
rect 93470 10164 93526 10220
rect 130082 10164 130138 10220
rect 130186 10164 130242 10220
rect 130290 10164 130346 10220
rect 38032 9380 38088 9436
rect 38136 9380 38192 9436
rect 38240 9380 38296 9436
rect 74852 9380 74908 9436
rect 74956 9380 75012 9436
rect 75060 9380 75116 9436
rect 111672 9380 111728 9436
rect 111776 9380 111832 9436
rect 111880 9380 111936 9436
rect 148492 9380 148548 9436
rect 148596 9380 148652 9436
rect 148700 9380 148756 9436
rect 19622 8596 19678 8652
rect 19726 8596 19782 8652
rect 19830 8596 19886 8652
rect 56442 8596 56498 8652
rect 56546 8596 56602 8652
rect 56650 8596 56706 8652
rect 93262 8596 93318 8652
rect 93366 8596 93422 8652
rect 93470 8596 93526 8652
rect 130082 8596 130138 8652
rect 130186 8596 130242 8652
rect 130290 8596 130346 8652
rect 38032 7812 38088 7868
rect 38136 7812 38192 7868
rect 38240 7812 38296 7868
rect 74852 7812 74908 7868
rect 74956 7812 75012 7868
rect 75060 7812 75116 7868
rect 111672 7812 111728 7868
rect 111776 7812 111832 7868
rect 111880 7812 111936 7868
rect 148492 7812 148548 7868
rect 148596 7812 148652 7868
rect 148700 7812 148756 7868
rect 19622 7028 19678 7084
rect 19726 7028 19782 7084
rect 19830 7028 19886 7084
rect 56442 7028 56498 7084
rect 56546 7028 56602 7084
rect 56650 7028 56706 7084
rect 93262 7028 93318 7084
rect 93366 7028 93422 7084
rect 93470 7028 93526 7084
rect 130082 7028 130138 7084
rect 130186 7028 130242 7084
rect 130290 7028 130346 7084
rect 38032 6244 38088 6300
rect 38136 6244 38192 6300
rect 38240 6244 38296 6300
rect 74852 6244 74908 6300
rect 74956 6244 75012 6300
rect 75060 6244 75116 6300
rect 111672 6244 111728 6300
rect 111776 6244 111832 6300
rect 111880 6244 111936 6300
rect 148492 6244 148548 6300
rect 148596 6244 148652 6300
rect 148700 6244 148756 6300
rect 19622 5460 19678 5516
rect 19726 5460 19782 5516
rect 19830 5460 19886 5516
rect 56442 5460 56498 5516
rect 56546 5460 56602 5516
rect 56650 5460 56706 5516
rect 93262 5460 93318 5516
rect 93366 5460 93422 5516
rect 93470 5460 93526 5516
rect 130082 5460 130138 5516
rect 130186 5460 130242 5516
rect 130290 5460 130346 5516
rect 38032 4676 38088 4732
rect 38136 4676 38192 4732
rect 38240 4676 38296 4732
rect 74852 4676 74908 4732
rect 74956 4676 75012 4732
rect 75060 4676 75116 4732
rect 111672 4676 111728 4732
rect 111776 4676 111832 4732
rect 111880 4676 111936 4732
rect 148492 4676 148548 4732
rect 148596 4676 148652 4732
rect 148700 4676 148756 4732
rect 19622 3892 19678 3948
rect 19726 3892 19782 3948
rect 19830 3892 19886 3948
rect 56442 3892 56498 3948
rect 56546 3892 56602 3948
rect 56650 3892 56706 3948
rect 93262 3892 93318 3948
rect 93366 3892 93422 3948
rect 93470 3892 93526 3948
rect 130082 3892 130138 3948
rect 130186 3892 130242 3948
rect 130290 3892 130346 3948
rect 38032 3108 38088 3164
rect 38136 3108 38192 3164
rect 38240 3108 38296 3164
rect 74852 3108 74908 3164
rect 74956 3108 75012 3164
rect 75060 3108 75116 3164
rect 111672 3108 111728 3164
rect 111776 3108 111832 3164
rect 111880 3108 111936 3164
rect 148492 3108 148548 3164
rect 148596 3108 148652 3164
rect 148700 3108 148756 3164
<< metal4 >>
rect 19594 36876 19914 36908
rect 19594 36820 19622 36876
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19886 36820 19914 36876
rect 19594 35308 19914 36820
rect 19594 35252 19622 35308
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19886 35252 19914 35308
rect 19594 33740 19914 35252
rect 19594 33684 19622 33740
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19886 33684 19914 33740
rect 19594 32172 19914 33684
rect 19594 32116 19622 32172
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19886 32116 19914 32172
rect 19594 30604 19914 32116
rect 19594 30548 19622 30604
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19886 30548 19914 30604
rect 19594 29036 19914 30548
rect 19594 28980 19622 29036
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19886 28980 19914 29036
rect 19594 27468 19914 28980
rect 19594 27412 19622 27468
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19886 27412 19914 27468
rect 19594 25900 19914 27412
rect 19594 25844 19622 25900
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19886 25844 19914 25900
rect 19594 24332 19914 25844
rect 19594 24276 19622 24332
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19886 24276 19914 24332
rect 19594 22764 19914 24276
rect 19594 22708 19622 22764
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19886 22708 19914 22764
rect 19594 21196 19914 22708
rect 19594 21140 19622 21196
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19886 21140 19914 21196
rect 19594 19628 19914 21140
rect 19594 19572 19622 19628
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19886 19572 19914 19628
rect 19594 18060 19914 19572
rect 19594 18004 19622 18060
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19886 18004 19914 18060
rect 19594 16492 19914 18004
rect 19594 16436 19622 16492
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19886 16436 19914 16492
rect 19594 14924 19914 16436
rect 19594 14868 19622 14924
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19886 14868 19914 14924
rect 19594 13356 19914 14868
rect 19594 13300 19622 13356
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19886 13300 19914 13356
rect 19594 11788 19914 13300
rect 19594 11732 19622 11788
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19886 11732 19914 11788
rect 19594 10220 19914 11732
rect 19594 10164 19622 10220
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19886 10164 19914 10220
rect 19594 8652 19914 10164
rect 19594 8596 19622 8652
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19886 8596 19914 8652
rect 19594 7084 19914 8596
rect 19594 7028 19622 7084
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19886 7028 19914 7084
rect 19594 5516 19914 7028
rect 19594 5460 19622 5516
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19886 5460 19914 5516
rect 19594 3948 19914 5460
rect 19594 3892 19622 3948
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19886 3892 19914 3948
rect 19594 3076 19914 3892
rect 38004 36092 38324 36908
rect 38004 36036 38032 36092
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38296 36036 38324 36092
rect 38004 34524 38324 36036
rect 38004 34468 38032 34524
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38296 34468 38324 34524
rect 38004 32956 38324 34468
rect 56414 36876 56734 36908
rect 56414 36820 56442 36876
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56706 36820 56734 36876
rect 56414 35308 56734 36820
rect 56414 35252 56442 35308
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56706 35252 56734 35308
rect 43596 33908 43652 33918
rect 43596 33684 43652 33852
rect 43596 33618 43652 33628
rect 56414 33740 56734 35252
rect 56414 33684 56442 33740
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56706 33684 56734 33740
rect 38004 32900 38032 32956
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38296 32900 38324 32956
rect 38004 31388 38324 32900
rect 38004 31332 38032 31388
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38296 31332 38324 31388
rect 38004 29820 38324 31332
rect 38004 29764 38032 29820
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38296 29764 38324 29820
rect 38004 28252 38324 29764
rect 38004 28196 38032 28252
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38296 28196 38324 28252
rect 38004 26684 38324 28196
rect 38004 26628 38032 26684
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38296 26628 38324 26684
rect 38004 25116 38324 26628
rect 38004 25060 38032 25116
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38296 25060 38324 25116
rect 38004 23548 38324 25060
rect 38004 23492 38032 23548
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38296 23492 38324 23548
rect 38004 21980 38324 23492
rect 38004 21924 38032 21980
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38296 21924 38324 21980
rect 38004 20412 38324 21924
rect 38004 20356 38032 20412
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38296 20356 38324 20412
rect 38004 18844 38324 20356
rect 38004 18788 38032 18844
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38296 18788 38324 18844
rect 38004 17276 38324 18788
rect 38004 17220 38032 17276
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38296 17220 38324 17276
rect 38004 15708 38324 17220
rect 38004 15652 38032 15708
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38296 15652 38324 15708
rect 38004 14140 38324 15652
rect 38004 14084 38032 14140
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38296 14084 38324 14140
rect 38004 12572 38324 14084
rect 38004 12516 38032 12572
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38296 12516 38324 12572
rect 38004 11004 38324 12516
rect 38004 10948 38032 11004
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38296 10948 38324 11004
rect 38004 9436 38324 10948
rect 38004 9380 38032 9436
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38296 9380 38324 9436
rect 38004 7868 38324 9380
rect 38004 7812 38032 7868
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38296 7812 38324 7868
rect 38004 6300 38324 7812
rect 38004 6244 38032 6300
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38296 6244 38324 6300
rect 38004 4732 38324 6244
rect 38004 4676 38032 4732
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38296 4676 38324 4732
rect 38004 3164 38324 4676
rect 38004 3108 38032 3164
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38296 3108 38324 3164
rect 38004 3076 38324 3108
rect 56414 32172 56734 33684
rect 74824 36092 75144 36908
rect 93234 36876 93554 36908
rect 93234 36820 93262 36876
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93526 36820 93554 36876
rect 74824 36036 74852 36092
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 75116 36036 75144 36092
rect 74824 34524 75144 36036
rect 75628 36372 75684 36382
rect 75628 35140 75684 36316
rect 91420 36036 91476 36046
rect 91476 35980 91588 36036
rect 91420 35970 91476 35980
rect 82236 35924 82292 35934
rect 75628 35074 75684 35084
rect 77084 35588 77140 35598
rect 74824 34468 74852 34524
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 75116 34468 75144 34524
rect 74824 32956 75144 34468
rect 77084 34356 77140 35532
rect 82236 34468 82292 35868
rect 91532 35812 91588 35980
rect 91532 35746 91588 35756
rect 82236 34402 82292 34412
rect 93234 35308 93554 36820
rect 93234 35252 93262 35308
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93526 35252 93554 35308
rect 77084 34290 77140 34300
rect 56414 32116 56442 32172
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56706 32116 56734 32172
rect 56414 30604 56734 32116
rect 56414 30548 56442 30604
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56706 30548 56734 30604
rect 56414 29036 56734 30548
rect 56414 28980 56442 29036
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56706 28980 56734 29036
rect 56414 27468 56734 28980
rect 56414 27412 56442 27468
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56706 27412 56734 27468
rect 56414 25900 56734 27412
rect 56414 25844 56442 25900
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56706 25844 56734 25900
rect 56414 24332 56734 25844
rect 58828 32900 58884 32910
rect 58828 25172 58884 32844
rect 58828 25106 58884 25116
rect 74824 32900 74852 32956
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 75116 32900 75144 32956
rect 74824 31388 75144 32900
rect 74824 31332 74852 31388
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 75116 31332 75144 31388
rect 74824 29820 75144 31332
rect 74824 29764 74852 29820
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 75116 29764 75144 29820
rect 74824 28252 75144 29764
rect 74824 28196 74852 28252
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 75116 28196 75144 28252
rect 74824 26684 75144 28196
rect 74824 26628 74852 26684
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 75116 26628 75144 26684
rect 74824 25116 75144 26628
rect 56414 24276 56442 24332
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56706 24276 56734 24332
rect 56414 22764 56734 24276
rect 56414 22708 56442 22764
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56706 22708 56734 22764
rect 56414 21196 56734 22708
rect 56414 21140 56442 21196
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56706 21140 56734 21196
rect 56414 19628 56734 21140
rect 56414 19572 56442 19628
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56706 19572 56734 19628
rect 56414 18060 56734 19572
rect 56414 18004 56442 18060
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56706 18004 56734 18060
rect 56414 16492 56734 18004
rect 56414 16436 56442 16492
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56706 16436 56734 16492
rect 56414 14924 56734 16436
rect 56414 14868 56442 14924
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56706 14868 56734 14924
rect 56414 13356 56734 14868
rect 56414 13300 56442 13356
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56706 13300 56734 13356
rect 56414 11788 56734 13300
rect 56414 11732 56442 11788
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56706 11732 56734 11788
rect 56414 10220 56734 11732
rect 56414 10164 56442 10220
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56706 10164 56734 10220
rect 56414 8652 56734 10164
rect 56414 8596 56442 8652
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56706 8596 56734 8652
rect 56414 7084 56734 8596
rect 56414 7028 56442 7084
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56706 7028 56734 7084
rect 56414 5516 56734 7028
rect 56414 5460 56442 5516
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56706 5460 56734 5516
rect 56414 3948 56734 5460
rect 56414 3892 56442 3948
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56706 3892 56734 3948
rect 56414 3076 56734 3892
rect 74824 25060 74852 25116
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 75116 25060 75144 25116
rect 74824 23548 75144 25060
rect 74824 23492 74852 23548
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 75116 23492 75144 23548
rect 74824 21980 75144 23492
rect 74824 21924 74852 21980
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 75116 21924 75144 21980
rect 74824 20412 75144 21924
rect 74824 20356 74852 20412
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 75116 20356 75144 20412
rect 74824 18844 75144 20356
rect 74824 18788 74852 18844
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 75116 18788 75144 18844
rect 74824 17276 75144 18788
rect 74824 17220 74852 17276
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 75116 17220 75144 17276
rect 74824 15708 75144 17220
rect 74824 15652 74852 15708
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 75116 15652 75144 15708
rect 74824 14140 75144 15652
rect 74824 14084 74852 14140
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 75116 14084 75144 14140
rect 74824 12572 75144 14084
rect 74824 12516 74852 12572
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 75116 12516 75144 12572
rect 74824 11004 75144 12516
rect 74824 10948 74852 11004
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 75116 10948 75144 11004
rect 74824 9436 75144 10948
rect 74824 9380 74852 9436
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 75116 9380 75144 9436
rect 74824 7868 75144 9380
rect 74824 7812 74852 7868
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 75116 7812 75144 7868
rect 74824 6300 75144 7812
rect 74824 6244 74852 6300
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 75116 6244 75144 6300
rect 74824 4732 75144 6244
rect 74824 4676 74852 4732
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 75116 4676 75144 4732
rect 74824 3164 75144 4676
rect 74824 3108 74852 3164
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 75116 3108 75144 3164
rect 74824 3076 75144 3108
rect 93234 33740 93554 35252
rect 93234 33684 93262 33740
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93526 33684 93554 33740
rect 93234 32172 93554 33684
rect 93234 32116 93262 32172
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93526 32116 93554 32172
rect 93234 30604 93554 32116
rect 111644 36092 111964 36908
rect 111644 36036 111672 36092
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111936 36036 111964 36092
rect 111644 34524 111964 36036
rect 130054 36876 130374 36908
rect 130054 36820 130082 36876
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130346 36820 130374 36876
rect 130054 35308 130374 36820
rect 130054 35252 130082 35308
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130346 35252 130374 35308
rect 115052 35028 115108 35038
rect 115052 34692 115108 34972
rect 115052 34626 115108 34636
rect 111644 34468 111672 34524
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111936 34468 111964 34524
rect 111644 32956 111964 34468
rect 111644 32900 111672 32956
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111936 32900 111964 32956
rect 105756 32004 105812 32014
rect 105756 31556 105812 31948
rect 105756 31490 105812 31500
rect 93234 30548 93262 30604
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93526 30548 93554 30604
rect 93234 29036 93554 30548
rect 93234 28980 93262 29036
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93526 28980 93554 29036
rect 93234 27468 93554 28980
rect 93234 27412 93262 27468
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93526 27412 93554 27468
rect 93234 25900 93554 27412
rect 93234 25844 93262 25900
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93526 25844 93554 25900
rect 93234 24332 93554 25844
rect 93234 24276 93262 24332
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93526 24276 93554 24332
rect 93234 22764 93554 24276
rect 93234 22708 93262 22764
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93526 22708 93554 22764
rect 93234 21196 93554 22708
rect 93234 21140 93262 21196
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93526 21140 93554 21196
rect 93234 19628 93554 21140
rect 93234 19572 93262 19628
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93526 19572 93554 19628
rect 93234 18060 93554 19572
rect 93234 18004 93262 18060
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93526 18004 93554 18060
rect 93234 16492 93554 18004
rect 93234 16436 93262 16492
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93526 16436 93554 16492
rect 93234 14924 93554 16436
rect 93234 14868 93262 14924
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93526 14868 93554 14924
rect 93234 13356 93554 14868
rect 93234 13300 93262 13356
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93526 13300 93554 13356
rect 93234 11788 93554 13300
rect 93234 11732 93262 11788
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93526 11732 93554 11788
rect 93234 10220 93554 11732
rect 93234 10164 93262 10220
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93526 10164 93554 10220
rect 93234 8652 93554 10164
rect 93234 8596 93262 8652
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93526 8596 93554 8652
rect 93234 7084 93554 8596
rect 93234 7028 93262 7084
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93526 7028 93554 7084
rect 93234 5516 93554 7028
rect 93234 5460 93262 5516
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93526 5460 93554 5516
rect 93234 3948 93554 5460
rect 93234 3892 93262 3948
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93526 3892 93554 3948
rect 93234 3076 93554 3892
rect 111644 31388 111964 32900
rect 111644 31332 111672 31388
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111936 31332 111964 31388
rect 111644 29820 111964 31332
rect 111644 29764 111672 29820
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111936 29764 111964 29820
rect 111644 28252 111964 29764
rect 111644 28196 111672 28252
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111936 28196 111964 28252
rect 111644 26684 111964 28196
rect 111644 26628 111672 26684
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111936 26628 111964 26684
rect 111644 25116 111964 26628
rect 111644 25060 111672 25116
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111936 25060 111964 25116
rect 111644 23548 111964 25060
rect 111644 23492 111672 23548
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111936 23492 111964 23548
rect 111644 21980 111964 23492
rect 111644 21924 111672 21980
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111936 21924 111964 21980
rect 111644 20412 111964 21924
rect 111644 20356 111672 20412
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111936 20356 111964 20412
rect 111644 18844 111964 20356
rect 111644 18788 111672 18844
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111936 18788 111964 18844
rect 111644 17276 111964 18788
rect 111644 17220 111672 17276
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111936 17220 111964 17276
rect 111644 15708 111964 17220
rect 111644 15652 111672 15708
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111936 15652 111964 15708
rect 111644 14140 111964 15652
rect 111644 14084 111672 14140
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111936 14084 111964 14140
rect 111644 12572 111964 14084
rect 111644 12516 111672 12572
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111936 12516 111964 12572
rect 111644 11004 111964 12516
rect 111644 10948 111672 11004
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111936 10948 111964 11004
rect 111644 9436 111964 10948
rect 111644 9380 111672 9436
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111936 9380 111964 9436
rect 111644 7868 111964 9380
rect 111644 7812 111672 7868
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111936 7812 111964 7868
rect 111644 6300 111964 7812
rect 111644 6244 111672 6300
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111936 6244 111964 6300
rect 111644 4732 111964 6244
rect 111644 4676 111672 4732
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111936 4676 111964 4732
rect 111644 3164 111964 4676
rect 111644 3108 111672 3164
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111936 3108 111964 3164
rect 111644 3076 111964 3108
rect 130054 33740 130374 35252
rect 130054 33684 130082 33740
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130346 33684 130374 33740
rect 130054 32172 130374 33684
rect 130054 32116 130082 32172
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130346 32116 130374 32172
rect 130054 30604 130374 32116
rect 130054 30548 130082 30604
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130346 30548 130374 30604
rect 130054 29036 130374 30548
rect 130054 28980 130082 29036
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130346 28980 130374 29036
rect 130054 27468 130374 28980
rect 130054 27412 130082 27468
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130346 27412 130374 27468
rect 130054 25900 130374 27412
rect 130054 25844 130082 25900
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130346 25844 130374 25900
rect 130054 24332 130374 25844
rect 130054 24276 130082 24332
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130346 24276 130374 24332
rect 130054 22764 130374 24276
rect 130054 22708 130082 22764
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130346 22708 130374 22764
rect 130054 21196 130374 22708
rect 130054 21140 130082 21196
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130346 21140 130374 21196
rect 130054 19628 130374 21140
rect 130054 19572 130082 19628
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130346 19572 130374 19628
rect 130054 18060 130374 19572
rect 130054 18004 130082 18060
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130346 18004 130374 18060
rect 130054 16492 130374 18004
rect 130054 16436 130082 16492
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130346 16436 130374 16492
rect 130054 14924 130374 16436
rect 130054 14868 130082 14924
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130346 14868 130374 14924
rect 130054 13356 130374 14868
rect 130054 13300 130082 13356
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130346 13300 130374 13356
rect 130054 11788 130374 13300
rect 130054 11732 130082 11788
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130346 11732 130374 11788
rect 130054 10220 130374 11732
rect 130054 10164 130082 10220
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130346 10164 130374 10220
rect 130054 8652 130374 10164
rect 130054 8596 130082 8652
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130346 8596 130374 8652
rect 130054 7084 130374 8596
rect 130054 7028 130082 7084
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130346 7028 130374 7084
rect 130054 5516 130374 7028
rect 130054 5460 130082 5516
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130346 5460 130374 5516
rect 130054 3948 130374 5460
rect 130054 3892 130082 3948
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130346 3892 130374 3948
rect 130054 3076 130374 3892
rect 148464 36092 148784 36908
rect 148464 36036 148492 36092
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148756 36036 148784 36092
rect 148464 34524 148784 36036
rect 148464 34468 148492 34524
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148756 34468 148784 34524
rect 148464 32956 148784 34468
rect 148464 32900 148492 32956
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148756 32900 148784 32956
rect 148464 31388 148784 32900
rect 148464 31332 148492 31388
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148756 31332 148784 31388
rect 148464 29820 148784 31332
rect 148464 29764 148492 29820
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148756 29764 148784 29820
rect 148464 28252 148784 29764
rect 148464 28196 148492 28252
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148756 28196 148784 28252
rect 148464 26684 148784 28196
rect 148464 26628 148492 26684
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148756 26628 148784 26684
rect 148464 25116 148784 26628
rect 148464 25060 148492 25116
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148756 25060 148784 25116
rect 148464 23548 148784 25060
rect 148464 23492 148492 23548
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148756 23492 148784 23548
rect 148464 21980 148784 23492
rect 148464 21924 148492 21980
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148756 21924 148784 21980
rect 148464 20412 148784 21924
rect 148464 20356 148492 20412
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148756 20356 148784 20412
rect 148464 18844 148784 20356
rect 148464 18788 148492 18844
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148756 18788 148784 18844
rect 148464 17276 148784 18788
rect 148464 17220 148492 17276
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148756 17220 148784 17276
rect 148464 15708 148784 17220
rect 148464 15652 148492 15708
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148756 15652 148784 15708
rect 148464 14140 148784 15652
rect 148464 14084 148492 14140
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148756 14084 148784 14140
rect 148464 12572 148784 14084
rect 148464 12516 148492 12572
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148756 12516 148784 12572
rect 148464 11004 148784 12516
rect 148464 10948 148492 11004
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148756 10948 148784 11004
rect 148464 9436 148784 10948
rect 148464 9380 148492 9436
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148756 9380 148784 9436
rect 148464 7868 148784 9380
rect 148464 7812 148492 7868
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148756 7812 148784 7868
rect 148464 6300 148784 7812
rect 148464 6244 148492 6300
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148756 6244 148784 6300
rect 148464 4732 148784 6244
rect 148464 4676 148492 4732
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148756 4676 148784 4732
rect 148464 3164 148784 4676
rect 148464 3108 148492 3164
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148756 3108 148784 3164
rect 148464 3076 148784 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__I dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 63392 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__I0
timestamp 1669390400
transform 1 0 92736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__I1
timestamp 1669390400
transform -1 0 94864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__S
timestamp 1669390400
transform 1 0 93744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__I
timestamp 1669390400
transform 1 0 49728 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__I
timestamp 1669390400
transform 1 0 140784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I0
timestamp 1669390400
transform 1 0 131264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I1
timestamp 1669390400
transform 1 0 128688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__S
timestamp 1669390400
transform 1 0 130816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__I0
timestamp 1669390400
transform -1 0 88704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__I1
timestamp 1669390400
transform -1 0 91952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__S
timestamp 1669390400
transform 1 0 88928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I0
timestamp 1669390400
transform -1 0 126112 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I1
timestamp 1669390400
transform 1 0 126336 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__S
timestamp 1669390400
transform -1 0 127120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__I
timestamp 1669390400
transform 1 0 63168 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1669390400
transform 1 0 110656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__I0
timestamp 1669390400
transform -1 0 142464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__S
timestamp 1669390400
transform 1 0 141792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I0
timestamp 1669390400
transform 1 0 141680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I1
timestamp 1669390400
transform 1 0 144816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__S
timestamp 1669390400
transform -1 0 141456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I0
timestamp 1669390400
transform -1 0 142912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__S
timestamp 1669390400
transform 1 0 143920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I0
timestamp 1669390400
transform -1 0 141344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I1
timestamp 1669390400
transform 1 0 143920 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__S
timestamp 1669390400
transform 1 0 143472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I0
timestamp 1669390400
transform -1 0 112000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I1
timestamp 1669390400
transform -1 0 114688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__S
timestamp 1669390400
transform 1 0 110880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1669390400
transform 1 0 110432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__I0
timestamp 1669390400
transform -1 0 116368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__I1
timestamp 1669390400
transform 1 0 115696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__S
timestamp 1669390400
transform 1 0 113568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I0
timestamp 1669390400
transform 1 0 121520 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I1
timestamp 1669390400
transform -1 0 120736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__S
timestamp 1669390400
transform -1 0 118832 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__I1
timestamp 1669390400
transform 1 0 120512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__S
timestamp 1669390400
transform -1 0 118384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__I
timestamp 1669390400
transform -1 0 105504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__I0
timestamp 1669390400
transform -1 0 112560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__I1
timestamp 1669390400
transform 1 0 115024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__S
timestamp 1669390400
transform 1 0 111888 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__I1
timestamp 1669390400
transform 1 0 115584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__S
timestamp 1669390400
transform -1 0 113456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__I0
timestamp 1669390400
transform -1 0 105952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__I1
timestamp 1669390400
transform -1 0 107744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__S
timestamp 1669390400
transform -1 0 106400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I0
timestamp 1669390400
transform 1 0 110656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I1
timestamp 1669390400
transform 1 0 107856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__S
timestamp 1669390400
transform -1 0 110432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__I0
timestamp 1669390400
transform -1 0 136416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__S
timestamp 1669390400
transform 1 0 139664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__I
timestamp 1669390400
transform 1 0 140784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__I0
timestamp 1669390400
transform 1 0 139664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__I1
timestamp 1669390400
transform 1 0 140112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I0
timestamp 1669390400
transform -1 0 137088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I1
timestamp 1669390400
transform 1 0 137312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__S
timestamp 1669390400
transform 1 0 137312 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__I0
timestamp 1669390400
transform 1 0 137872 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__I1
timestamp 1669390400
transform 1 0 140224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I
timestamp 1669390400
transform 1 0 63840 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__I
timestamp 1669390400
transform 1 0 105056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__I0
timestamp 1669390400
transform 1 0 129248 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__S
timestamp 1669390400
transform 1 0 128800 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I0
timestamp 1669390400
transform 1 0 143472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I1
timestamp 1669390400
transform 1 0 145824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__I0
timestamp 1669390400
transform -1 0 130032 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__S
timestamp 1669390400
transform 1 0 129360 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__I0
timestamp 1669390400
transform 1 0 146720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__I1
timestamp 1669390400
transform 1 0 145264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__I0
timestamp 1669390400
transform -1 0 121856 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__S
timestamp 1669390400
transform 1 0 123984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__I
timestamp 1669390400
transform 1 0 51072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__I
timestamp 1669390400
transform 1 0 90048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__I0
timestamp 1669390400
transform -1 0 121184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__I1
timestamp 1669390400
transform 1 0 123312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__S
timestamp 1669390400
transform 1 0 122864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__I0
timestamp 1669390400
transform -1 0 119392 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__S
timestamp 1669390400
transform -1 0 119840 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__I0
timestamp 1669390400
transform 1 0 120960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__I1
timestamp 1669390400
transform 1 0 121408 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__S
timestamp 1669390400
transform 1 0 117488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__I
timestamp 1669390400
transform 1 0 101472 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__I0
timestamp 1669390400
transform -1 0 98336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__I1
timestamp 1669390400
transform -1 0 102144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__S
timestamp 1669390400
transform 1 0 101024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__I0
timestamp 1669390400
transform -1 0 101696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__I1
timestamp 1669390400
transform 1 0 101024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__S
timestamp 1669390400
transform 1 0 98448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__I0
timestamp 1669390400
transform -1 0 89376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__I1
timestamp 1669390400
transform -1 0 93296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__S
timestamp 1669390400
transform -1 0 90832 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__I0
timestamp 1669390400
transform -1 0 93744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__I1
timestamp 1669390400
transform 1 0 90384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__S
timestamp 1669390400
transform 1 0 93072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__I0
timestamp 1669390400
transform 1 0 91280 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__I1
timestamp 1669390400
transform -1 0 91728 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__S
timestamp 1669390400
transform -1 0 91280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__I
timestamp 1669390400
transform 1 0 87360 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__I0
timestamp 1669390400
transform 1 0 88928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__I1
timestamp 1669390400
transform 1 0 88480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__S
timestamp 1669390400
transform 1 0 89600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__I0
timestamp 1669390400
transform -1 0 93072 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__I1
timestamp 1669390400
transform -1 0 95312 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__S
timestamp 1669390400
transform 1 0 95536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__I0
timestamp 1669390400
transform -1 0 91504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__I1
timestamp 1669390400
transform 1 0 90832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__S
timestamp 1669390400
transform 1 0 89152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__I
timestamp 1669390400
transform 1 0 75040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__I0
timestamp 1669390400
transform -1 0 74816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__I1
timestamp 1669390400
transform -1 0 78288 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__S
timestamp 1669390400
transform 1 0 78960 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__I1
timestamp 1669390400
transform 1 0 75488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__S
timestamp 1669390400
transform -1 0 74144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__I0
timestamp 1669390400
transform -1 0 76608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__I1
timestamp 1669390400
transform -1 0 78736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__S
timestamp 1669390400
transform -1 0 76160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__I1
timestamp 1669390400
transform 1 0 78288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__S
timestamp 1669390400
transform 1 0 77840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__I0
timestamp 1669390400
transform -1 0 67200 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__I1
timestamp 1669390400
transform -1 0 69440 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__S
timestamp 1669390400
transform -1 0 66864 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__I
timestamp 1669390400
transform 1 0 60816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__I1
timestamp 1669390400
transform -1 0 66752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__I0
timestamp 1669390400
transform -1 0 67760 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__I1
timestamp 1669390400
transform -1 0 69888 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__S
timestamp 1669390400
transform 1 0 69440 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__I0
timestamp 1669390400
transform -1 0 69216 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__I1
timestamp 1669390400
transform 1 0 69440 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__I
timestamp 1669390400
transform -1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__I0
timestamp 1669390400
transform 1 0 65744 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__I1
timestamp 1669390400
transform -1 0 67200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__S
timestamp 1669390400
transform 1 0 62608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__I0
timestamp 1669390400
transform 1 0 67200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__I1
timestamp 1669390400
transform 1 0 67648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__I0
timestamp 1669390400
transform -1 0 64512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__I1
timestamp 1669390400
transform -1 0 65744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__S
timestamp 1669390400
transform 1 0 66192 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__I0
timestamp 1669390400
transform 1 0 64624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__I1
timestamp 1669390400
transform 1 0 67200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__I0
timestamp 1669390400
transform -1 0 47600 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__I1
timestamp 1669390400
transform -1 0 50848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__S
timestamp 1669390400
transform -1 0 50624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__I
timestamp 1669390400
transform -1 0 51632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__I1
timestamp 1669390400
transform 1 0 51520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__S
timestamp 1669390400
transform 1 0 51072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__I0
timestamp 1669390400
transform -1 0 44800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__I1
timestamp 1669390400
transform -1 0 45696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__S
timestamp 1669390400
transform -1 0 48272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__I1
timestamp 1669390400
transform 1 0 48720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__S
timestamp 1669390400
transform -1 0 48496 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__I
timestamp 1669390400
transform 1 0 62272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__I0
timestamp 1669390400
transform -1 0 36736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__I1
timestamp 1669390400
transform -1 0 39536 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__S
timestamp 1669390400
transform -1 0 39088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__I1
timestamp 1669390400
transform 1 0 39200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__S
timestamp 1669390400
transform -1 0 39872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__I0
timestamp 1669390400
transform -1 0 35840 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__I1
timestamp 1669390400
transform -1 0 42112 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__S
timestamp 1669390400
transform -1 0 40880 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__I1
timestamp 1669390400
transform -1 0 40208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__S
timestamp 1669390400
transform 1 0 40432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__I0
timestamp 1669390400
transform 1 0 29232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__I1
timestamp 1669390400
transform -1 0 32368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__S
timestamp 1669390400
transform 1 0 32592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__I
timestamp 1669390400
transform 1 0 20720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__I1
timestamp 1669390400
transform -1 0 31584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__S
timestamp 1669390400
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__I0
timestamp 1669390400
transform -1 0 29456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__I1
timestamp 1669390400
transform -1 0 31920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__S
timestamp 1669390400
transform 1 0 30800 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__I1
timestamp 1669390400
transform 1 0 29120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__S
timestamp 1669390400
transform 1 0 26320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__I1
timestamp 1669390400
transform -1 0 22848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__S
timestamp 1669390400
transform -1 0 22176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__I1
timestamp 1669390400
transform 1 0 21952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__S
timestamp 1669390400
transform -1 0 17920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__I0
timestamp 1669390400
transform -1 0 17920 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__I1
timestamp 1669390400
transform -1 0 20832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__S
timestamp 1669390400
transform -1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__I1
timestamp 1669390400
transform -1 0 20048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__S
timestamp 1669390400
transform 1 0 20272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__A1
timestamp 1669390400
transform 1 0 14896 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__A2
timestamp 1669390400
transform -1 0 14000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__288__I
timestamp 1669390400
transform 1 0 52640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__A1
timestamp 1669390400
transform 1 0 69664 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__A2
timestamp 1669390400
transform -1 0 68992 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A1
timestamp 1669390400
transform 1 0 51296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A2
timestamp 1669390400
transform -1 0 52640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__I
timestamp 1669390400
transform -1 0 56560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__I
timestamp 1669390400
transform 1 0 58800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__I
timestamp 1669390400
transform 1 0 30016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__I
timestamp 1669390400
transform 1 0 22176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__I
timestamp 1669390400
transform -1 0 21280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__I
timestamp 1669390400
transform 1 0 30688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__I
timestamp 1669390400
transform 1 0 32480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__I
timestamp 1669390400
transform 1 0 55888 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__I
timestamp 1669390400
transform 1 0 57232 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__I
timestamp 1669390400
transform -1 0 40992 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__I
timestamp 1669390400
transform -1 0 42336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__I
timestamp 1669390400
transform -1 0 48160 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__I
timestamp 1669390400
transform -1 0 54208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__I
timestamp 1669390400
transform 1 0 71904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__I
timestamp 1669390400
transform -1 0 64400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__I
timestamp 1669390400
transform 1 0 69888 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__I
timestamp 1669390400
transform 1 0 71680 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__I
timestamp 1669390400
transform -1 0 64736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__I
timestamp 1669390400
transform -1 0 92512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__I
timestamp 1669390400
transform 1 0 81200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__I
timestamp 1669390400
transform 1 0 81648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__I
timestamp 1669390400
transform 1 0 93072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__314__I
timestamp 1669390400
transform 1 0 92176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__I
timestamp 1669390400
transform 1 0 93632 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__I
timestamp 1669390400
transform 1 0 98336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__I
timestamp 1669390400
transform 1 0 102480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__318__I
timestamp 1669390400
transform 1 0 120960 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__I
timestamp 1669390400
transform -1 0 116032 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__I
timestamp 1669390400
transform 1 0 135408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__I
timestamp 1669390400
transform 1 0 108304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__I
timestamp 1669390400
transform 1 0 134512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__I
timestamp 1669390400
transform 1 0 15792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__I
timestamp 1669390400
transform 1 0 12208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__I
timestamp 1669390400
transform -1 0 12544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__CLK
timestamp 1669390400
transform 1 0 21504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__CLK
timestamp 1669390400
transform 1 0 21504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__CLK
timestamp 1669390400
transform 1 0 29456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__CLK
timestamp 1669390400
transform 1 0 31808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__CLK
timestamp 1669390400
transform 1 0 41440 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__CLK
timestamp 1669390400
transform -1 0 40320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__CLK
timestamp 1669390400
transform -1 0 48944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__CLK
timestamp 1669390400
transform 1 0 54432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__CLK
timestamp 1669390400
transform 1 0 60592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__CLK
timestamp 1669390400
transform -1 0 68768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__CLK
timestamp 1669390400
transform 1 0 72128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__CLK
timestamp 1669390400
transform 1 0 63168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__CLK
timestamp 1669390400
transform -1 0 80528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__CLK
timestamp 1669390400
transform -1 0 76832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__CLK
timestamp 1669390400
transform 1 0 86240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__CLK
timestamp 1669390400
transform 1 0 84448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__CLK
timestamp 1669390400
transform -1 0 94976 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__CLK
timestamp 1669390400
transform 1 0 99008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__CLK
timestamp 1669390400
transform 1 0 116704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__CLK
timestamp 1669390400
transform -1 0 116256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__CLK
timestamp 1669390400
transform 1 0 126784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__D
timestamp 1669390400
transform 1 0 132832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__RN
timestamp 1669390400
transform -1 0 132384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__CLK
timestamp 1669390400
transform -1 0 129360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__D
timestamp 1669390400
transform -1 0 133168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__CLK
timestamp 1669390400
transform 1 0 124208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__D
timestamp 1669390400
transform -1 0 128576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__CLK
timestamp 1669390400
transform 1 0 134176 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__CLK
timestamp 1669390400
transform 1 0 107520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__CLK
timestamp 1669390400
transform 1 0 113008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__CLK
timestamp 1669390400
transform 1 0 117152 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__CLK
timestamp 1669390400
transform 1 0 112000 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__CLK
timestamp 1669390400
transform -1 0 128128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__D
timestamp 1669390400
transform 1 0 136864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__CLK
timestamp 1669390400
transform 1 0 126896 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__D
timestamp 1669390400
transform -1 0 133616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__CLK
timestamp 1669390400
transform 1 0 127344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__CLK
timestamp 1669390400
transform 1 0 127344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__CLK
timestamp 1669390400
transform 1 0 16912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__D
timestamp 1669390400
transform 1 0 12656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__CLK
timestamp 1669390400
transform 1 0 11312 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__372__CLK
timestamp 1669390400
transform 1 0 11200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__I
timestamp 1669390400
transform 1 0 8512 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__I
timestamp 1669390400
transform 1 0 11648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__I
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__I
timestamp 1669390400
transform -1 0 21504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__379__I
timestamp 1669390400
transform 1 0 38416 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__380__I
timestamp 1669390400
transform 1 0 42112 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__I
timestamp 1669390400
transform 1 0 48944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__I
timestamp 1669390400
transform 1 0 49392 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__I
timestamp 1669390400
transform 1 0 46480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__I
timestamp 1669390400
transform 1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__385__I
timestamp 1669390400
transform 1 0 39872 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__I
timestamp 1669390400
transform -1 0 45360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__I
timestamp 1669390400
transform 1 0 59808 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__I
timestamp 1669390400
transform 1 0 57120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__I
timestamp 1669390400
transform 1 0 77616 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__I
timestamp 1669390400
transform 1 0 83776 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__I
timestamp 1669390400
transform 1 0 80528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__I
timestamp 1669390400
transform 1 0 76272 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__393__I
timestamp 1669390400
transform -1 0 6160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__I
timestamp 1669390400
transform -1 0 10080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__I
timestamp 1669390400
transform 1 0 14896 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__I
timestamp 1669390400
transform 1 0 19712 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__I
timestamp 1669390400
transform -1 0 31584 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__I
timestamp 1669390400
transform 1 0 37632 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__I
timestamp 1669390400
transform 1 0 34496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__I
timestamp 1669390400
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__I
timestamp 1669390400
transform 1 0 46928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__I
timestamp 1669390400
transform 1 0 48496 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__I
timestamp 1669390400
transform 1 0 51968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__I
timestamp 1669390400
transform -1 0 41216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__I
timestamp 1669390400
transform 1 0 52416 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__I
timestamp 1669390400
transform -1 0 53760 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__I
timestamp 1669390400
transform 1 0 73696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__I
timestamp 1669390400
transform -1 0 59584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__I
timestamp 1669390400
transform 1 0 57792 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__I
timestamp 1669390400
transform 1 0 54880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__I
timestamp 1669390400
transform -1 0 56336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__I
timestamp 1669390400
transform 1 0 70784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__I
timestamp 1669390400
transform 1 0 61824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__I
timestamp 1669390400
transform 1 0 84560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__415__I
timestamp 1669390400
transform -1 0 88256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__I
timestamp 1669390400
transform 1 0 100240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__I
timestamp 1669390400
transform 1 0 110432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__418__I
timestamp 1669390400
transform 1 0 118496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__I
timestamp 1669390400
transform 1 0 120064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__I
timestamp 1669390400
transform 1 0 127904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__I
timestamp 1669390400
transform -1 0 138096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__I
timestamp 1669390400
transform 1 0 124880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__I
timestamp 1669390400
transform 1 0 79408 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__424__I
timestamp 1669390400
transform 1 0 74144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__I
timestamp 1669390400
transform 1 0 15568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__I
timestamp 1669390400
transform 1 0 21504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__I
timestamp 1669390400
transform 1 0 35616 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__I
timestamp 1669390400
transform 1 0 41552 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__I
timestamp 1669390400
transform 1 0 58240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__I
timestamp 1669390400
transform 1 0 64288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__431__I
timestamp 1669390400
transform 1 0 87584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__I
timestamp 1669390400
transform 1 0 98560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__I
timestamp 1669390400
transform 1 0 93520 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__I
timestamp 1669390400
transform 1 0 91952 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__I
timestamp 1669390400
transform 1 0 84896 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__I
timestamp 1669390400
transform 1 0 97216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__I
timestamp 1669390400
transform 1 0 105504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__I
timestamp 1669390400
transform 1 0 108640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__I
timestamp 1669390400
transform 1 0 111328 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__I
timestamp 1669390400
transform 1 0 116928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__I
timestamp 1669390400
transform 1 0 117376 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__I
timestamp 1669390400
transform 1 0 122080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__I
timestamp 1669390400
transform 1 0 124768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__I
timestamp 1669390400
transform 1 0 107968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__I
timestamp 1669390400
transform 1 0 114016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__I
timestamp 1669390400
transform 1 0 117824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__I
timestamp 1669390400
transform 1 0 128912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__I
timestamp 1669390400
transform 1 0 133952 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__449__I
timestamp 1669390400
transform 1 0 131376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__I
timestamp 1669390400
transform 1 0 131936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__I
timestamp 1669390400
transform 1 0 133168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__I
timestamp 1669390400
transform 1 0 134736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__453__I
timestamp 1669390400
transform 1 0 140896 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__I
timestamp 1669390400
transform 1 0 139552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__I
timestamp 1669390400
transform 1 0 145712 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__456__I
timestamp 1669390400
transform 1 0 145600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__I
timestamp 1669390400
transform 1 0 9856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__I
timestamp 1669390400
transform 1 0 15008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__I
timestamp 1669390400
transform 1 0 18816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__I
timestamp 1669390400
transform -1 0 17920 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__461__I
timestamp 1669390400
transform 1 0 38080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__I
timestamp 1669390400
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__I
timestamp 1669390400
transform 1 0 28336 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__I
timestamp 1669390400
transform 1 0 41216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_io_wbs_clk_I
timestamp 1669390400
transform 1 0 70672 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_io_wbs_clk_I
timestamp 1669390400
transform 1 0 72576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_io_wbs_clk_I
timestamp 1669390400
transform -1 0 68320 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_io_wbs_clk_I
timestamp 1669390400
transform 1 0 73472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_io_wbs_clk_I
timestamp 1669390400
transform -1 0 76384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform 1 0 9632 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 36960 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 37520 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform -1 0 41664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 42784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform -1 0 43680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform -1 0 45584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform 1 0 47600 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform 1 0 49840 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform -1 0 49280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform -1 0 53536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1669390400
transform 1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1669390400
transform -1 0 53200 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1669390400
transform -1 0 56896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1669390400
transform 1 0 59584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1669390400
transform -1 0 60256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1669390400
transform -1 0 57120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1669390400
transform 1 0 64848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1669390400
transform -1 0 60928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1669390400
transform 1 0 67648 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1669390400
transform -1 0 68544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1669390400
transform -1 0 71456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1669390400
transform -1 0 14000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1669390400
transform -1 0 72800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1669390400
transform -1 0 71792 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1669390400
transform -1 0 19488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1669390400
transform -1 0 21504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1669390400
transform -1 0 25312 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1669390400
transform -1 0 28000 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1669390400
transform -1 0 27776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1669390400
transform -1 0 33488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1669390400
transform -1 0 33600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1669390400
transform 1 0 82992 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1669390400
transform 1 0 109536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1669390400
transform -1 0 110208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1669390400
transform 1 0 114352 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1669390400
transform 1 0 116032 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1669390400
transform 1 0 118272 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1669390400
transform -1 0 117152 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1669390400
transform 1 0 122192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1669390400
transform -1 0 121184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1669390400
transform 1 0 126112 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1669390400
transform 1 0 125216 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1669390400
transform -1 0 82656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1669390400
transform -1 0 126336 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1669390400
transform 1 0 130368 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1669390400
transform 1 0 132160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1669390400
transform -1 0 131040 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1669390400
transform 1 0 134288 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1669390400
transform -1 0 135408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1669390400
transform -1 0 136864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1669390400
transform 1 0 140112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1669390400
transform -1 0 140224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1669390400
transform -1 0 142800 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1669390400
transform 1 0 89040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1669390400
transform -1 0 143360 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1669390400
transform 1 0 146832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1669390400
transform 1 0 92400 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1669390400
transform -1 0 94192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1669390400
transform 1 0 99008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1669390400
transform 1 0 103600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1669390400
transform -1 0 101696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1669390400
transform -1 0 104160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1669390400
transform 1 0 108864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1669390400
transform -1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1669390400
transform -1 0 61936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1669390400
transform 1 0 25200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1669390400
transform -1 0 27552 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1669390400
transform -1 0 33824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1669390400
transform -1 0 37856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1669390400
transform -1 0 41888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1669390400
transform -1 0 45920 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1669390400
transform -1 0 49952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1669390400
transform -1 0 53984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1669390400
transform -1 0 6944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1669390400
transform 1 0 19376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1669390400
transform -1 0 60592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1669390400
transform -1 0 60928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1669390400
transform 1 0 69888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1669390400
transform -1 0 72688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1669390400
transform -1 0 72688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1669390400
transform 1 0 84000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1669390400
transform 1 0 87920 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input84_I
timestamp 1669390400
transform 1 0 91840 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input85_I
timestamp 1669390400
transform 1 0 96208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input86_I
timestamp 1669390400
transform -1 0 96992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input87_I
timestamp 1669390400
transform 1 0 22176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input88_I
timestamp 1669390400
transform -1 0 101024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input89_I
timestamp 1669390400
transform -1 0 105056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input90_I
timestamp 1669390400
transform -1 0 108976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input91_I
timestamp 1669390400
transform 1 0 119952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input92_I
timestamp 1669390400
transform 1 0 123200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input93_I
timestamp 1669390400
transform 1 0 123648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input94_I
timestamp 1669390400
transform 1 0 127120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input95_I
timestamp 1669390400
transform 1 0 135632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input96_I
timestamp 1669390400
transform 1 0 137984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input97_I
timestamp 1669390400
transform -1 0 137536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input98_I
timestamp 1669390400
transform -1 0 25760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input99_I
timestamp 1669390400
transform -1 0 141344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input100_I
timestamp 1669390400
transform 1 0 147168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input101_I
timestamp 1669390400
transform 1 0 33488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input102_I
timestamp 1669390400
transform 1 0 36960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input103_I
timestamp 1669390400
transform 1 0 41216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input104_I
timestamp 1669390400
transform -1 0 45360 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input105_I
timestamp 1669390400
transform 1 0 49168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input106_I
timestamp 1669390400
transform -1 0 52640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input107_I
timestamp 1669390400
transform -1 0 57568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input108_I
timestamp 1669390400
transform 1 0 10080 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input109_I
timestamp 1669390400
transform -1 0 17808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input110_I
timestamp 1669390400
transform -1 0 21952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input111_I
timestamp 1669390400
transform -1 0 26656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input112_I
timestamp 1669390400
transform 1 0 33040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input113_I
timestamp 1669390400
transform -1 0 9856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input114_I
timestamp 1669390400
transform -1 0 11984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output119_I
timestamp 1669390400
transform -1 0 23296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output120_I
timestamp 1669390400
transform 1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output121_I
timestamp 1669390400
transform -1 0 27440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output122_I
timestamp 1669390400
transform 1 0 28784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output123_I
timestamp 1669390400
transform 1 0 33488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output124_I
timestamp 1669390400
transform -1 0 78064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output125_I
timestamp 1669390400
transform 1 0 82096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output126_I
timestamp 1669390400
transform -1 0 85232 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output127_I
timestamp 1669390400
transform -1 0 87808 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output128_I
timestamp 1669390400
transform 1 0 94192 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output129_I
timestamp 1669390400
transform 1 0 95088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output130_I
timestamp 1669390400
transform 1 0 96432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output131_I
timestamp 1669390400
transform 1 0 100240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output132_I
timestamp 1669390400
transform -1 0 102816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output134_I
timestamp 1669390400
transform 1 0 36064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output136_I
timestamp 1669390400
transform -1 0 41888 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output137_I
timestamp 1669390400
transform -1 0 43232 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output138_I
timestamp 1669390400
transform -1 0 44352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output139_I
timestamp 1669390400
transform -1 0 46032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output140_I
timestamp 1669390400
transform -1 0 48832 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output143_I
timestamp 1669390400
transform -1 0 53984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output146_I
timestamp 1669390400
transform -1 0 56448 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output147_I
timestamp 1669390400
transform -1 0 59248 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output148_I
timestamp 1669390400
transform -1 0 60816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output149_I
timestamp 1669390400
transform -1 0 62944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output150_I
timestamp 1669390400
transform -1 0 65520 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output151_I
timestamp 1669390400
transform -1 0 66752 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output152_I
timestamp 1669390400
transform -1 0 68208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output153_I
timestamp 1669390400
transform 1 0 71456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output154_I
timestamp 1669390400
transform 1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output159_I
timestamp 1669390400
transform -1 0 23744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output160_I
timestamp 1669390400
transform 1 0 24416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output162_I
timestamp 1669390400
transform -1 0 31472 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output163_I
timestamp 1669390400
transform 1 0 33936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output164_I
timestamp 1669390400
transform 1 0 35168 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output165_I
timestamp 1669390400
transform -1 0 79184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output166_I
timestamp 1669390400
transform -1 0 106848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output167_I
timestamp 1669390400
transform -1 0 109312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output175_I
timestamp 1669390400
transform -1 0 122976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output176_I
timestamp 1669390400
transform -1 0 81536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output177_I
timestamp 1669390400
transform 1 0 125664 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output178_I
timestamp 1669390400
transform 1 0 126560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output187_I
timestamp 1669390400
transform 1 0 88256 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output190_I
timestamp 1669390400
transform -1 0 89824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output191_I
timestamp 1669390400
transform -1 0 94864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output192_I
timestamp 1669390400
transform 1 0 95984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output193_I
timestamp 1669390400
transform 1 0 98896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output195_I
timestamp 1669390400
transform 1 0 102592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output196_I
timestamp 1669390400
transform -1 0 105056 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output197_I
timestamp 1669390400
transform -1 0 6496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output199_I
timestamp 1669390400
transform 1 0 59920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output203_I
timestamp 1669390400
transform -1 0 75152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output204_I
timestamp 1669390400
transform 1 0 81536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output205_I
timestamp 1669390400
transform 1 0 85568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output206_I
timestamp 1669390400
transform -1 0 86912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output207_I
timestamp 1669390400
transform -1 0 95984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output208_I
timestamp 1669390400
transform 1 0 97104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output210_I
timestamp 1669390400
transform 1 0 101696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output211_I
timestamp 1669390400
transform 1 0 105728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output212_I
timestamp 1669390400
transform 1 0 111104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output213_I
timestamp 1669390400
transform -1 0 114240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output214_I
timestamp 1669390400
transform 1 0 120400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output217_I
timestamp 1669390400
transform 1 0 126448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output218_I
timestamp 1669390400
transform 1 0 134960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output219_I
timestamp 1669390400
transform -1 0 139104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output221_I
timestamp 1669390400
transform -1 0 140000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output222_I
timestamp 1669390400
transform 1 0 146496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output228_I
timestamp 1669390400
transform 1 0 53312 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output229_I
timestamp 1669390400
transform -1 0 55104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output230_I
timestamp 1669390400
transform 1 0 7168 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output236_I
timestamp 1669390400
transform 1 0 79744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output237_I
timestamp 1669390400
transform 1 0 85456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output238_I
timestamp 1669390400
transform -1 0 87136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output239_I
timestamp 1669390400
transform 1 0 92176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41
timestamp 1669390400
transform 1 0 5936 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83
timestamp 1669390400
transform 1 0 10640 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87
timestamp 1669390400
transform 1 0 11088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113
timestamp 1669390400
transform 1 0 14000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121
timestamp 1669390400
transform 1 0 14896 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_159
timestamp 1669390400
transform 1 0 19152 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_163 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 19600 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_171
timestamp 1669390400
transform 1 0 20496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_181
timestamp 1669390400
transform 1 0 21616 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_184
timestamp 1669390400
transform 1 0 21952 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188
timestamp 1669390400
transform 1 0 22400 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_192
timestamp 1669390400
transform 1 0 22848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_215
timestamp 1669390400
transform 1 0 25424 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_223
timestamp 1669390400
transform 1 0 26320 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_226
timestamp 1669390400
transform 1 0 26656 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_254
timestamp 1669390400
transform 1 0 29792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_258
timestamp 1669390400
transform 1 0 30240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_262
timestamp 1669390400
transform 1 0 30688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1669390400
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_285
timestamp 1669390400
transform 1 0 33264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_293
timestamp 1669390400
transform 1 0 34160 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_297
timestamp 1669390400
transform 1 0 34608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1669390400
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_320
timestamp 1669390400
transform 1 0 37184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_326
timestamp 1669390400
transform 1 0 37856 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_344
timestamp 1669390400
transform 1 0 39872 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_348
timestamp 1669390400
transform 1 0 40320 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_358
timestamp 1669390400
transform 1 0 41440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_362
timestamp 1669390400
transform 1 0 41888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_380
timestamp 1669390400
transform 1 0 43904 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1669390400
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_395
timestamp 1669390400
transform 1 0 45584 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_398
timestamp 1669390400
transform 1 0 45920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_416
timestamp 1669390400
transform 1 0 47936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_425
timestamp 1669390400
transform 1 0 48944 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_429
timestamp 1669390400
transform 1 0 49392 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_431
timestamp 1669390400
transform 1 0 49616 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_434
timestamp 1669390400
transform 1 0 49952 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_452
timestamp 1669390400
transform 1 0 51968 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1669390400
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_465
timestamp 1669390400
transform 1 0 53424 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_467
timestamp 1669390400
transform 1 0 53648 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_470
timestamp 1669390400
transform 1 0 53984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_488
timestamp 1669390400
transform 1 0 56000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_499
timestamp 1669390400
transform 1 0 57232 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_503
timestamp 1669390400
transform 1 0 57680 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_506
timestamp 1669390400
transform 1 0 58016 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_524
timestamp 1669390400
transform 1 0 60032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_527
timestamp 1669390400
transform 1 0 60368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_529
timestamp 1669390400
transform 1 0 60592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_532
timestamp 1669390400
transform 1 0 60928 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_559
timestamp 1669390400
transform 1 0 63952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_562
timestamp 1669390400
transform 1 0 64288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_566
timestamp 1669390400
transform 1 0 64736 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_593
timestamp 1669390400
transform 1 0 67760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1669390400
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_602
timestamp 1669390400
transform 1 0 68768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_629
timestamp 1669390400
transform 1 0 71792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_632
timestamp 1669390400
transform 1 0 72128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_634
timestamp 1669390400
transform 1 0 72352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_637
timestamp 1669390400
transform 1 0 72688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1669390400
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1669390400
transform 1 0 76048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_670
timestamp 1669390400
transform 1 0 76384 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_674
timestamp 1669390400
transform 1 0 76832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_692
timestamp 1669390400
transform 1 0 78848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_698
timestamp 1669390400
transform 1 0 79520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_702
timestamp 1669390400
transform 1 0 79968 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_707
timestamp 1669390400
transform 1 0 80528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_734
timestamp 1669390400
transform 1 0 83552 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_737
timestamp 1669390400
transform 1 0 83888 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_740
timestamp 1669390400
transform 1 0 84224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_769
timestamp 1669390400
transform 1 0 87472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_772
timestamp 1669390400
transform 1 0 87808 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_775
timestamp 1669390400
transform 1 0 88144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_804
timestamp 1669390400
transform 1 0 91392 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_807
timestamp 1669390400
transform 1 0 91728 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_810
timestamp 1669390400
transform 1 0 92064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_839
timestamp 1669390400
transform 1 0 95312 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_842
timestamp 1669390400
transform 1 0 95648 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_845
timestamp 1669390400
transform 1 0 95984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_849
timestamp 1669390400
transform 1 0 96432 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_851
timestamp 1669390400
transform 1 0 96656 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_854
timestamp 1669390400
transform 1 0 96992 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_872
timestamp 1669390400
transform 1 0 99008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_874
timestamp 1669390400
transform 1 0 99232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_877
timestamp 1669390400
transform 1 0 99568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_885
timestamp 1669390400
transform 1 0 100464 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_887
timestamp 1669390400
transform 1 0 100688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_890
timestamp 1669390400
transform 1 0 101024 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_908
timestamp 1669390400
transform 1 0 103040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_912
timestamp 1669390400
transform 1 0 103488 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_920
timestamp 1669390400
transform 1 0 104384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_926
timestamp 1669390400
transform 1 0 105056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_944
timestamp 1669390400
transform 1 0 107072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_947
timestamp 1669390400
transform 1 0 107408 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_957
timestamp 1669390400
transform 1 0 108528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_961
timestamp 1669390400
transform 1 0 108976 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_979
timestamp 1669390400
transform 1 0 110992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_982
timestamp 1669390400
transform 1 0 111328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_988
timestamp 1669390400
transform 1 0 112000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_996
timestamp 1669390400
transform 1 0 112896 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1014
timestamp 1669390400
transform 1 0 114912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1017
timestamp 1669390400
transform 1 0 115248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1022
timestamp 1669390400
transform 1 0 115808 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1028
timestamp 1669390400
transform 1 0 116480 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1032
timestamp 1669390400
transform 1 0 116928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1049
timestamp 1669390400
transform 1 0 118832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1052
timestamp 1669390400
transform 1 0 119168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1057
timestamp 1669390400
transform 1 0 119728 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1061
timestamp 1669390400
transform 1 0 120176 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1065
timestamp 1669390400
transform 1 0 120624 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1067
timestamp 1669390400
transform 1 0 120848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1084
timestamp 1669390400
transform 1 0 122752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1087
timestamp 1669390400
transform 1 0 123088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1090
timestamp 1669390400
transform 1 0 123424 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1094
timestamp 1669390400
transform 1 0 123872 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1102
timestamp 1669390400
transform 1 0 124768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1119
timestamp 1669390400
transform 1 0 126672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1122
timestamp 1669390400
transform 1 0 127008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1125
timestamp 1669390400
transform 1 0 127344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1129
timestamp 1669390400
transform 1 0 127792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1132
timestamp 1669390400
transform 1 0 128128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1136
timestamp 1669390400
transform 1 0 128576 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1154
timestamp 1669390400
transform 1 0 130592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1157
timestamp 1669390400
transform 1 0 130928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1165
timestamp 1669390400
transform 1 0 131824 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1171
timestamp 1669390400
transform 1 0 132496 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1189
timestamp 1669390400
transform 1 0 134512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1192
timestamp 1669390400
transform 1 0 134848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1197
timestamp 1669390400
transform 1 0 135408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1201
timestamp 1669390400
transform 1 0 135856 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1203
timestamp 1669390400
transform 1 0 136080 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1218
timestamp 1669390400
transform 1 0 137760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1222
timestamp 1669390400
transform 1 0 138208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1224
timestamp 1669390400
transform 1 0 138432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1227
timestamp 1669390400
transform 1 0 138768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1230
timestamp 1669390400
transform 1 0 139104 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1234
timestamp 1669390400
transform 1 0 139552 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1238
timestamp 1669390400
transform 1 0 140000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1254
timestamp 1669390400
transform 1 0 141792 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1258
timestamp 1669390400
transform 1 0 142240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1262
timestamp 1669390400
transform 1 0 142688 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1276
timestamp 1669390400
transform 1 0 144256 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1294
timestamp 1669390400
transform 1 0 146272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1297
timestamp 1669390400
transform 1 0 146608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1312
timestamp 1669390400
transform 1 0 148288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_18
timestamp 1669390400
transform 1 0 3360 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_26
timestamp 1669390400
transform 1 0 4256 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_42
timestamp 1669390400
transform 1 0 6048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_46
timestamp 1669390400
transform 1 0 6496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_50
timestamp 1669390400
transform 1 0 6944 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_68
timestamp 1669390400
transform 1 0 8960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_75
timestamp 1669390400
transform 1 0 9744 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_92
timestamp 1669390400
transform 1 0 11648 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_98
timestamp 1669390400
transform 1 0 12320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_102
timestamp 1669390400
transform 1 0 12768 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_137
timestamp 1669390400
transform 1 0 16688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_147
timestamp 1669390400
transform 1 0 17808 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_149
timestamp 1669390400
transform 1 0 18032 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_164
timestamp 1669390400
transform 1 0 19712 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_182
timestamp 1669390400
transform 1 0 21728 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_200
timestamp 1669390400
transform 1 0 23744 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1669390400
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_218
timestamp 1669390400
transform 1 0 25760 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_236
timestamp 1669390400
transform 1 0 27776 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_242
timestamp 1669390400
transform 1 0 28448 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_260
timestamp 1669390400
transform 1 0 30464 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_264
timestamp 1669390400
transform 1 0 30912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_266
timestamp 1669390400
transform 1 0 31136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_289
timestamp 1669390400
transform 1 0 33712 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_297
timestamp 1669390400
transform 1 0 34608 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_301
timestamp 1669390400
transform 1 0 35056 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_303
timestamp 1669390400
transform 1 0 35280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_338
timestamp 1669390400
transform 1 0 39200 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_374
timestamp 1669390400
transform 1 0 43232 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_390
timestamp 1669390400
transform 1 0 45024 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_445
timestamp 1669390400
transform 1 0 51184 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_449
timestamp 1669390400
transform 1 0 51632 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_453
timestamp 1669390400
transform 1 0 52080 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_455
timestamp 1669390400
transform 1 0 52304 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_458
timestamp 1669390400
transform 1 0 52640 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_476
timestamp 1669390400
transform 1 0 54656 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_480
timestamp 1669390400
transform 1 0 55104 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1669390400
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_516
timestamp 1669390400
transform 1 0 59136 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_524
timestamp 1669390400
transform 1 0 60032 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_528
timestamp 1669390400
transform 1 0 60480 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_531
timestamp 1669390400
transform 1 0 60816 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1669390400
transform 1 0 64848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1669390400
transform 1 0 65184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_621
timestamp 1669390400
transform 1 0 70896 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_623
timestamp 1669390400
transform 1 0 71120 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_638
timestamp 1669390400
transform 1 0 72800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_641
timestamp 1669390400
transform 1 0 73136 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_657
timestamp 1669390400
transform 1 0 74928 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_709
timestamp 1669390400
transform 1 0 80752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_712
timestamp 1669390400
transform 1 0 81088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_715
timestamp 1669390400
transform 1 0 81424 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_719
timestamp 1669390400
transform 1 0 81872 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_735
timestamp 1669390400
transform 1 0 83664 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_750
timestamp 1669390400
transform 1 0 85344 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_754
timestamp 1669390400
transform 1 0 85792 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_760
timestamp 1669390400
transform 1 0 86464 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_764
timestamp 1669390400
transform 1 0 86912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_780
timestamp 1669390400
transform 1 0 88704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_783
timestamp 1669390400
transform 1 0 89040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_818
timestamp 1669390400
transform 1 0 92960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_834
timestamp 1669390400
transform 1 0 94752 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_836
timestamp 1669390400
transform 1 0 94976 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_851
timestamp 1669390400
transform 1 0 96656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_854
timestamp 1669390400
transform 1 0 96992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_857
timestamp 1669390400
transform 1 0 97328 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_859
timestamp 1669390400
transform 1 0 97552 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_864
timestamp 1669390400
transform 1 0 98112 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_868
timestamp 1669390400
transform 1 0 98560 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_874
timestamp 1669390400
transform 1 0 99232 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_910
timestamp 1669390400
transform 1 0 103264 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_918
timestamp 1669390400
transform 1 0 104160 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_922
timestamp 1669390400
transform 1 0 104608 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_925
timestamp 1669390400
transform 1 0 104944 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_941
timestamp 1669390400
transform 1 0 106736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_945
timestamp 1669390400
transform 1 0 107184 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_947
timestamp 1669390400
transform 1 0 107408 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_950
timestamp 1669390400
transform 1 0 107744 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_986
timestamp 1669390400
transform 1 0 111776 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_990
timestamp 1669390400
transform 1 0 112224 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_996
timestamp 1669390400
transform 1 0 112896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1031
timestamp 1669390400
transform 1 0 116816 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1047
timestamp 1669390400
transform 1 0 118608 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1055
timestamp 1669390400
transform 1 0 119504 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1061
timestamp 1669390400
transform 1 0 120176 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1067
timestamp 1669390400
transform 1 0 120848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1082
timestamp 1669390400
transform 1 0 122528 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1090
timestamp 1669390400
transform 1 0 123424 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1094
timestamp 1669390400
transform 1 0 123872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1096
timestamp 1669390400
transform 1 0 124096 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1099
timestamp 1669390400
transform 1 0 124432 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1135
timestamp 1669390400
transform 1 0 128464 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1138
timestamp 1669390400
transform 1 0 128800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1173
timestamp 1669390400
transform 1 0 132720 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1189
timestamp 1669390400
transform 1 0 134512 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1197
timestamp 1669390400
transform 1 0 135408 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1199
timestamp 1669390400
transform 1 0 135632 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1206
timestamp 1669390400
transform 1 0 136416 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1209
timestamp 1669390400
transform 1 0 136752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1212
timestamp 1669390400
transform 1 0 137088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1232
timestamp 1669390400
transform 1 0 139328 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1250
timestamp 1669390400
transform 1 0 141344 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1268
timestamp 1669390400
transform 1 0 143360 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1276
timestamp 1669390400
transform 1 0 144256 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1280
timestamp 1669390400
transform 1 0 144704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1296
timestamp 1669390400
transform 1 0 146496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1300
timestamp 1669390400
transform 1 0 146944 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1304
timestamp 1669390400
transform 1 0 147392 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1312
timestamp 1669390400
transform 1 0 148288 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_89
timestamp 1669390400
transform 1 0 11312 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_95
timestamp 1669390400
transform 1 0 11984 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_99
timestamp 1669390400
transform 1 0 12432 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_103
timestamp 1669390400
transform 1 0 12880 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_126
timestamp 1669390400
transform 1 0 15456 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_128
timestamp 1669390400
transform 1 0 15680 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_131
timestamp 1669390400
transform 1 0 16016 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_137
timestamp 1669390400
transform 1 0 16688 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_175
timestamp 1669390400
transform 1 0 20944 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_184
timestamp 1669390400
transform 1 0 21952 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_188
timestamp 1669390400
transform 1 0 22400 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_204
timestamp 1669390400
transform 1 0 24192 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_208
timestamp 1669390400
transform 1 0 24640 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_210
timestamp 1669390400
transform 1 0 24864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_245
timestamp 1669390400
transform 1 0 28784 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_253
timestamp 1669390400
transform 1 0 29680 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_255
timestamp 1669390400
transform 1 0 29904 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_270
timestamp 1669390400
transform 1 0 31584 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_276
timestamp 1669390400
transform 1 0 32256 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_280
timestamp 1669390400
transform 1 0 32704 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_290
timestamp 1669390400
transform 1 0 33824 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_308
timestamp 1669390400
transform 1 0 35840 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_356
timestamp 1669390400
transform 1 0 41216 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_362
timestamp 1669390400
transform 1 0 41888 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_366
timestamp 1669390400
transform 1 0 42336 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_374
timestamp 1669390400
transform 1 0 43232 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_409
timestamp 1669390400
transform 1 0 47152 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_413
timestamp 1669390400
transform 1 0 47600 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_415
timestamp 1669390400
transform 1 0 47824 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_418
timestamp 1669390400
transform 1 0 48160 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_424
timestamp 1669390400
transform 1 0 48832 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1669390400
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_468
timestamp 1669390400
transform 1 0 53760 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_472
timestamp 1669390400
transform 1 0 54208 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_476
timestamp 1669390400
transform 1 0 54656 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_484
timestamp 1669390400
transform 1 0 55552 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_486
timestamp 1669390400
transform 1 0 55776 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_489
timestamp 1669390400
transform 1 0 56112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_497
timestamp 1669390400
transform 1 0 57008 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_501
timestamp 1669390400
transform 1 0 57456 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_509
timestamp 1669390400
transform 1 0 58352 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_515
timestamp 1669390400
transform 1 0 59024 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1669390400
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_534
timestamp 1669390400
transform 1 0 61152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_585
timestamp 1669390400
transform 1 0 66864 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_602
timestamp 1669390400
transform 1 0 68768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1669390400
transform 1 0 69104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_620
timestamp 1669390400
transform 1 0 70784 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_628
timestamp 1669390400
transform 1 0 71680 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_632
timestamp 1669390400
transform 1 0 72128 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_634
timestamp 1669390400
transform 1 0 72352 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_637
timestamp 1669390400
transform 1 0 72688 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1669390400
transform 1 0 76720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_676
timestamp 1669390400
transform 1 0 77056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_727
timestamp 1669390400
transform 1 0 82768 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_735
timestamp 1669390400
transform 1 0 83664 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_739
timestamp 1669390400
transform 1 0 84112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_741
timestamp 1669390400
transform 1 0 84336 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_744
timestamp 1669390400
transform 1 0 84672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_747
timestamp 1669390400
transform 1 0 85008 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_783
timestamp 1669390400
transform 1 0 89040 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_789
timestamp 1669390400
transform 1 0 89712 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_791
timestamp 1669390400
transform 1 0 89936 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_794
timestamp 1669390400
transform 1 0 90272 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_796
timestamp 1669390400
transform 1 0 90496 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_803
timestamp 1669390400
transform 1 0 91280 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_809
timestamp 1669390400
transform 1 0 91952 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_813
timestamp 1669390400
transform 1 0 92400 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_815
timestamp 1669390400
transform 1 0 92624 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_818
timestamp 1669390400
transform 1 0 92960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_821
timestamp 1669390400
transform 1 0 93296 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_823
timestamp 1669390400
transform 1 0 93520 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_826
timestamp 1669390400
transform 1 0 93856 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_834
timestamp 1669390400
transform 1 0 94752 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_870
timestamp 1669390400
transform 1 0 98784 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_886
timestamp 1669390400
transform 1 0 100576 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_889
timestamp 1669390400
transform 1 0 100912 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_901
timestamp 1669390400
transform 1 0 102256 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_905
timestamp 1669390400
transform 1 0 102704 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_913
timestamp 1669390400
transform 1 0 103600 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_915
timestamp 1669390400
transform 1 0 103824 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_930
timestamp 1669390400
transform 1 0 105504 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_934
timestamp 1669390400
transform 1 0 105952 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_950
timestamp 1669390400
transform 1 0 107744 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_957
timestamp 1669390400
transform 1 0 108528 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_960
timestamp 1669390400
transform 1 0 108864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_975
timestamp 1669390400
transform 1 0 110544 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_977
timestamp 1669390400
transform 1 0 110768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_984
timestamp 1669390400
transform 1 0 111552 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1020
timestamp 1669390400
transform 1 0 115584 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1028
timestamp 1669390400
transform 1 0 116480 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1031
timestamp 1669390400
transform 1 0 116816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1066
timestamp 1669390400
transform 1 0 120736 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1070
timestamp 1669390400
transform 1 0 121184 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1086
timestamp 1669390400
transform 1 0 122976 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1094
timestamp 1669390400
transform 1 0 123872 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1098
timestamp 1669390400
transform 1 0 124320 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1102
timestamp 1669390400
transform 1 0 124768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1117
timestamp 1669390400
transform 1 0 126448 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1123
timestamp 1669390400
transform 1 0 127120 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1127
timestamp 1669390400
transform 1 0 127568 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1163
timestamp 1669390400
transform 1 0 131600 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1169
timestamp 1669390400
transform 1 0 132272 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1173
timestamp 1669390400
transform 1 0 132720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1208
timestamp 1669390400
transform 1 0 136640 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1216
timestamp 1669390400
transform 1 0 137536 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1233
timestamp 1669390400
transform 1 0 139440 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1237
timestamp 1669390400
transform 1 0 139888 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1241
timestamp 1669390400
transform 1 0 140336 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1244
timestamp 1669390400
transform 1 0 140672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1247
timestamp 1669390400
transform 1 0 141008 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1251
timestamp 1669390400
transform 1 0 141456 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1255
timestamp 1669390400
transform 1 0 141904 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1265
timestamp 1669390400
transform 1 0 143024 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1271
timestamp 1669390400
transform 1 0 143696 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1288
timestamp 1669390400
transform 1 0 145600 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1292
timestamp 1669390400
transform 1 0 146048 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1298
timestamp 1669390400
transform 1 0 146720 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1306
timestamp 1669390400
transform 1 0 147616 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1310
timestamp 1669390400
transform 1 0 148064 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1312
timestamp 1669390400
transform 1 0 148288 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_34
timestamp 1669390400
transform 1 0 5152 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_50
timestamp 1669390400
transform 1 0 6944 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_58
timestamp 1669390400
transform 1 0 7840 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_65
timestamp 1669390400
transform 1 0 8624 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_69
timestamp 1669390400
transform 1 0 9072 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_76
timestamp 1669390400
transform 1 0 9856 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_80
timestamp 1669390400
transform 1 0 10304 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_88
timestamp 1669390400
transform 1 0 11200 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_91
timestamp 1669390400
transform 1 0 11536 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_95
timestamp 1669390400
transform 1 0 11984 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_97
timestamp 1669390400
transform 1 0 12208 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_100
timestamp 1669390400
transform 1 0 12544 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_116
timestamp 1669390400
transform 1 0 14336 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_120
timestamp 1669390400
transform 1 0 14784 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_123
timestamp 1669390400
transform 1 0 15120 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_133
timestamp 1669390400
transform 1 0 16240 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_148
timestamp 1669390400
transform 1 0 17920 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_165
timestamp 1669390400
transform 1 0 19824 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_169
timestamp 1669390400
transform 1 0 20272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_174
timestamp 1669390400
transform 1 0 20832 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_178
timestamp 1669390400
transform 1 0 21280 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_182
timestamp 1669390400
transform 1 0 21728 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_186
timestamp 1669390400
transform 1 0 22176 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_202
timestamp 1669390400
transform 1 0 23968 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_210
timestamp 1669390400
transform 1 0 24864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_230
timestamp 1669390400
transform 1 0 27104 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_234
timestamp 1669390400
transform 1 0 27552 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_270
timestamp 1669390400
transform 1 0 31584 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_274
timestamp 1669390400
transform 1 0 32032 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_282
timestamp 1669390400
transform 1 0 32928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_302
timestamp 1669390400
transform 1 0 35168 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_318
timestamp 1669390400
transform 1 0 36960 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_320
timestamp 1669390400
transform 1 0 37184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_336
timestamp 1669390400
transform 1 0 38976 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_344
timestamp 1669390400
transform 1 0 39872 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_350
timestamp 1669390400
transform 1 0 40544 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_360
timestamp 1669390400
transform 1 0 41664 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_376
timestamp 1669390400
transform 1 0 43456 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_384
timestamp 1669390400
transform 1 0 44352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_388
timestamp 1669390400
transform 1 0 44800 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_390
timestamp 1669390400
transform 1 0 45024 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_393
timestamp 1669390400
transform 1 0 45360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_401
timestamp 1669390400
transform 1 0 46256 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_409
timestamp 1669390400
transform 1 0 47152 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_430
timestamp 1669390400
transform 1 0 49504 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_439
timestamp 1669390400
transform 1 0 50512 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_443
timestamp 1669390400
transform 1 0 50960 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_446
timestamp 1669390400
transform 1 0 51296 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_462
timestamp 1669390400
transform 1 0 53088 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_466
timestamp 1669390400
transform 1 0 53536 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_482
timestamp 1669390400
transform 1 0 55328 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_490
timestamp 1669390400
transform 1 0 56224 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_493
timestamp 1669390400
transform 1 0 56560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_502
timestamp 1669390400
transform 1 0 57568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_518
timestamp 1669390400
transform 1 0 59360 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_522
timestamp 1669390400
transform 1 0 59808 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_525
timestamp 1669390400
transform 1 0 60144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_529
timestamp 1669390400
transform 1 0 60592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_533
timestamp 1669390400
transform 1 0 61040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_551
timestamp 1669390400
transform 1 0 63056 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1669390400
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_570
timestamp 1669390400
transform 1 0 65184 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_580
timestamp 1669390400
transform 1 0 66304 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_584
timestamp 1669390400
transform 1 0 66752 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_620
timestamp 1669390400
transform 1 0 70784 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_626
timestamp 1669390400
transform 1 0 71456 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_630
timestamp 1669390400
transform 1 0 71904 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_634
timestamp 1669390400
transform 1 0 72352 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1669390400
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_641
timestamp 1669390400
transform 1 0 73136 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_643
timestamp 1669390400
transform 1 0 73360 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_646
timestamp 1669390400
transform 1 0 73696 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_650
timestamp 1669390400
transform 1 0 74144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_667
timestamp 1669390400
transform 1 0 76048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_703
timestamp 1669390400
transform 1 0 80080 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_707
timestamp 1669390400
transform 1 0 80528 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_709
timestamp 1669390400
transform 1 0 80752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_712
timestamp 1669390400
transform 1 0 81088 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_744
timestamp 1669390400
transform 1 0 84672 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_752
timestamp 1669390400
transform 1 0 85568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_762
timestamp 1669390400
transform 1 0 86688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_766
timestamp 1669390400
transform 1 0 87136 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_770
timestamp 1669390400
transform 1 0 87584 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_780
timestamp 1669390400
transform 1 0 88704 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_783
timestamp 1669390400
transform 1 0 89040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_790
timestamp 1669390400
transform 1 0 89824 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_802
timestamp 1669390400
transform 1 0 91168 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_810
timestamp 1669390400
transform 1 0 92064 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_814
timestamp 1669390400
transform 1 0 92512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_830
timestamp 1669390400
transform 1 0 94304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_836
timestamp 1669390400
transform 1 0 94976 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_854
timestamp 1669390400
transform 1 0 96992 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_870
timestamp 1669390400
transform 1 0 98784 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_878
timestamp 1669390400
transform 1 0 99680 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_894
timestamp 1669390400
transform 1 0 101472 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_898
timestamp 1669390400
transform 1 0 101920 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_914
timestamp 1669390400
transform 1 0 103712 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_922
timestamp 1669390400
transform 1 0 104608 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_925
timestamp 1669390400
transform 1 0 104944 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_941
timestamp 1669390400
transform 1 0 106736 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_949
timestamp 1669390400
transform 1 0 107632 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_953
timestamp 1669390400
transform 1 0 108080 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_970
timestamp 1669390400
transform 1 0 109984 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_974
timestamp 1669390400
transform 1 0 110432 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_978
timestamp 1669390400
transform 1 0 110880 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_982
timestamp 1669390400
transform 1 0 111328 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_986
timestamp 1669390400
transform 1 0 111776 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_993
timestamp 1669390400
transform 1 0 112560 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_996
timestamp 1669390400
transform 1 0 112896 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_998
timestamp 1669390400
transform 1 0 113120 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1001
timestamp 1669390400
transform 1 0 113456 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1018
timestamp 1669390400
transform 1 0 115360 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1022
timestamp 1669390400
transform 1 0 115808 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1026
timestamp 1669390400
transform 1 0 116256 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1062
timestamp 1669390400
transform 1 0 120288 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1064
timestamp 1669390400
transform 1 0 120512 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1067
timestamp 1669390400
transform 1 0 120848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_1070
timestamp 1669390400
transform 1 0 121184 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1102
timestamp 1669390400
transform 1 0 124768 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1110
timestamp 1669390400
transform 1 0 125664 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1114
timestamp 1669390400
transform 1 0 126112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1116
timestamp 1669390400
transform 1 0 126336 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1119
timestamp 1669390400
transform 1 0 126672 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1135
timestamp 1669390400
transform 1 0 128464 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1138
timestamp 1669390400
transform 1 0 128800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1173
timestamp 1669390400
transform 1 0 132720 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1181
timestamp 1669390400
transform 1 0 133616 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1187
timestamp 1669390400
transform 1 0 134288 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1191
timestamp 1669390400
transform 1 0 134736 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1195
timestamp 1669390400
transform 1 0 135184 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1199
timestamp 1669390400
transform 1 0 135632 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1209
timestamp 1669390400
transform 1 0 136752 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1213
timestamp 1669390400
transform 1 0 137200 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1216
timestamp 1669390400
transform 1 0 137536 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1218
timestamp 1669390400
transform 1 0 137760 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1221
timestamp 1669390400
transform 1 0 138096 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1238
timestamp 1669390400
transform 1 0 140000 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1242
timestamp 1669390400
transform 1 0 140448 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1244
timestamp 1669390400
transform 1 0 140672 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1247
timestamp 1669390400
transform 1 0 141008 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1257
timestamp 1669390400
transform 1 0 142128 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1274
timestamp 1669390400
transform 1 0 144032 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1280
timestamp 1669390400
transform 1 0 144704 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1283
timestamp 1669390400
transform 1 0 145040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1287
timestamp 1669390400
transform 1 0 145488 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1303
timestamp 1669390400
transform 1 0 147280 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1311
timestamp 1669390400
transform 1 0 148176 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_45
timestamp 1669390400
transform 1 0 6384 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_49
timestamp 1669390400
transform 1 0 6832 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_51
timestamp 1669390400
transform 1 0 7056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_86
timestamp 1669390400
transform 1 0 10976 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_90
timestamp 1669390400
transform 1 0 11424 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_124
timestamp 1669390400
transform 1 0 15232 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_166
timestamp 1669390400
transform 1 0 19936 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_182
timestamp 1669390400
transform 1 0 21728 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_214
timestamp 1669390400
transform 1 0 25312 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_216
timestamp 1669390400
transform 1 0 25536 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_223
timestamp 1669390400
transform 1 0 26320 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_240
timestamp 1669390400
transform 1 0 28224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_244
timestamp 1669390400
transform 1 0 28672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_266
timestamp 1669390400
transform 1 0 31136 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_270
timestamp 1669390400
transform 1 0 31584 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_302
timestamp 1669390400
transform 1 0 35168 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_325
timestamp 1669390400
transform 1 0 37744 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_327
timestamp 1669390400
transform 1 0 37968 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_343
timestamp 1669390400
transform 1 0 39760 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_347
timestamp 1669390400
transform 1 0 40208 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_351
timestamp 1669390400
transform 1 0 40656 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_383
timestamp 1669390400
transform 1 0 44240 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_387
timestamp 1669390400
transform 1 0 44688 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_408
timestamp 1669390400
transform 1 0 47040 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_425
timestamp 1669390400
transform 1 0 48944 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_442
timestamp 1669390400
transform 1 0 50848 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_450
timestamp 1669390400
transform 1 0 51744 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_458
timestamp 1669390400
transform 1 0 52640 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1669390400
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_463 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 53200 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1669390400
transform 1 0 60368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1669390400
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_534
timestamp 1669390400
transform 1 0 61152 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_538
timestamp 1669390400
transform 1 0 61600 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_541
timestamp 1669390400
transform 1 0 61936 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_577
timestamp 1669390400
transform 1 0 65968 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_585
timestamp 1669390400
transform 1 0 66864 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1669390400
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_605
timestamp 1669390400
transform 1 0 69104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_610
timestamp 1669390400
transform 1 0 69664 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_614
timestamp 1669390400
transform 1 0 70112 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_618
timestamp 1669390400
transform 1 0 70560 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_621
timestamp 1669390400
transform 1 0 70896 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1669390400
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_676
timestamp 1669390400
transform 1 0 77056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_683
timestamp 1669390400
transform 1 0 77840 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_691
timestamp 1669390400
transform 1 0 78736 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_699
timestamp 1669390400
transform 1 0 79632 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_714
timestamp 1669390400
transform 1 0 81312 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_718
timestamp 1669390400
transform 1 0 81760 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_734
timestamp 1669390400
transform 1 0 83552 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_742
timestamp 1669390400
transform 1 0 84448 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_744
timestamp 1669390400
transform 1 0 84672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_747
timestamp 1669390400
transform 1 0 85008 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_778
timestamp 1669390400
transform 1 0 88480 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_795
timestamp 1669390400
transform 1 0 90384 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_812
timestamp 1669390400
transform 1 0 92288 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_818
timestamp 1669390400
transform 1 0 92960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_821
timestamp 1669390400
transform 1 0 93296 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_825
timestamp 1669390400
transform 1 0 93744 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_857
timestamp 1669390400
transform 1 0 97328 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_865
timestamp 1669390400
transform 1 0 98224 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_869
timestamp 1669390400
transform 1 0 98672 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_886
timestamp 1669390400
transform 1 0 100576 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_889
timestamp 1669390400
transform 1 0 100912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_892
timestamp 1669390400
transform 1 0 101248 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_896
timestamp 1669390400
transform 1 0 101696 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_928
timestamp 1669390400
transform 1 0 105280 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_944
timestamp 1669390400
transform 1 0 107072 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_952
timestamp 1669390400
transform 1 0 107968 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_956
timestamp 1669390400
transform 1 0 108416 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_960
timestamp 1669390400
transform 1 0 108864 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_968
timestamp 1669390400
transform 1 0 109760 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_972
timestamp 1669390400
transform 1 0 110208 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_976
timestamp 1669390400
transform 1 0 110656 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_986
timestamp 1669390400
transform 1 0 111776 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1002
timestamp 1669390400
transform 1 0 113568 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1019
timestamp 1669390400
transform 1 0 115472 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1023
timestamp 1669390400
transform 1 0 115920 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1027
timestamp 1669390400
transform 1 0 116368 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1031
timestamp 1669390400
transform 1 0 116816 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1033
timestamp 1669390400
transform 1 0 117040 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1036
timestamp 1669390400
transform 1 0 117376 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1072
timestamp 1669390400
transform 1 0 121408 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1080
timestamp 1669390400
transform 1 0 122304 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1096
timestamp 1669390400
transform 1 0 124096 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1102
timestamp 1669390400
transform 1 0 124768 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1118
timestamp 1669390400
transform 1 0 126560 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1120
timestamp 1669390400
transform 1 0 126784 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1123
timestamp 1669390400
transform 1 0 127120 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1127
timestamp 1669390400
transform 1 0 127568 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1163
timestamp 1669390400
transform 1 0 131600 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1169
timestamp 1669390400
transform 1 0 132272 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1173
timestamp 1669390400
transform 1 0 132720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1178
timestamp 1669390400
transform 1 0 133280 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1184
timestamp 1669390400
transform 1 0 133952 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_1188
timestamp 1669390400
transform 1 0 134400 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1220
timestamp 1669390400
transform 1 0 137984 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1236
timestamp 1669390400
transform 1 0 139776 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1240
timestamp 1669390400
transform 1 0 140224 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1244
timestamp 1669390400
transform 1 0 140672 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1250
timestamp 1669390400
transform 1 0 141344 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1267
timestamp 1669390400
transform 1 0 143248 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1271
timestamp 1669390400
transform 1 0 143696 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_1275
timestamp 1669390400
transform 1 0 144144 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1307
timestamp 1669390400
transform 1 0 147728 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1311
timestamp 1669390400
transform 1 0 148176 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1669390400
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1669390400
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_163
timestamp 1669390400
transform 1 0 19600 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_167
timestamp 1669390400
transform 1 0 20048 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_171
timestamp 1669390400
transform 1 0 20496 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_175
timestamp 1669390400
transform 1 0 20944 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_207
timestamp 1669390400
transform 1 0 24528 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_211
timestamp 1669390400
transform 1 0 24976 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_225
timestamp 1669390400
transform 1 0 26544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_233
timestamp 1669390400
transform 1 0 27440 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_237
timestamp 1669390400
transform 1 0 27888 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_239
timestamp 1669390400
transform 1 0 28112 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_246
timestamp 1669390400
transform 1 0 28896 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_250
timestamp 1669390400
transform 1 0 29344 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_282
timestamp 1669390400
transform 1 0 32928 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_318
timestamp 1669390400
transform 1 0 36960 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_334
timestamp 1669390400
transform 1 0 38752 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_340
timestamp 1669390400
transform 1 0 39424 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_344
timestamp 1669390400
transform 1 0 39872 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_352
timestamp 1669390400
transform 1 0 40768 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_389
timestamp 1669390400
transform 1 0 44912 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_405
timestamp 1669390400
transform 1 0 46704 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_413
timestamp 1669390400
transform 1 0 47600 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_417
timestamp 1669390400
transform 1 0 48048 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_421
timestamp 1669390400
transform 1 0 48496 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_434
timestamp 1669390400
transform 1 0 49952 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_442
timestamp 1669390400
transform 1 0 50848 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_446
timestamp 1669390400
transform 1 0 51296 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_450
timestamp 1669390400
transform 1 0 51744 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_482
timestamp 1669390400
transform 1 0 55328 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_490
timestamp 1669390400
transform 1 0 56224 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_494
timestamp 1669390400
transform 1 0 56672 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_531
timestamp 1669390400
transform 1 0 60816 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_539
timestamp 1669390400
transform 1 0 61712 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_543
timestamp 1669390400
transform 1 0 62160 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_551
timestamp 1669390400
transform 1 0 63056 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_553
timestamp 1669390400
transform 1 0 63280 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_560
timestamp 1669390400
transform 1 0 64064 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_562
timestamp 1669390400
transform 1 0 64288 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1669390400
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_570
timestamp 1669390400
transform 1 0 65184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_586
timestamp 1669390400
transform 1 0 66976 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_590
timestamp 1669390400
transform 1 0 67424 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_598
timestamp 1669390400
transform 1 0 68320 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_602
timestamp 1669390400
transform 1 0 68768 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_606
timestamp 1669390400
transform 1 0 69216 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_610
timestamp 1669390400
transform 1 0 69664 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_614
timestamp 1669390400
transform 1 0 70112 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_630
timestamp 1669390400
transform 1 0 71904 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1669390400
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_641
timestamp 1669390400
transform 1 0 73136 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_659
timestamp 1669390400
transform 1 0 75152 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_661
timestamp 1669390400
transform 1 0 75376 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_664
timestamp 1669390400
transform 1 0 75712 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_681
timestamp 1669390400
transform 1 0 77616 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_685
timestamp 1669390400
transform 1 0 78064 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_689
timestamp 1669390400
transform 1 0 78512 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_705
timestamp 1669390400
transform 1 0 80304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_709
timestamp 1669390400
transform 1 0 80752 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_712
timestamp 1669390400
transform 1 0 81088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_776
timestamp 1669390400
transform 1 0 88256 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_780
timestamp 1669390400
transform 1 0 88704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_783
timestamp 1669390400
transform 1 0 89040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_786
timestamp 1669390400
transform 1 0 89376 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_790
timestamp 1669390400
transform 1 0 89824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_794
timestamp 1669390400
transform 1 0 90272 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_797
timestamp 1669390400
transform 1 0 90608 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_801
timestamp 1669390400
transform 1 0 91056 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_805
timestamp 1669390400
transform 1 0 91504 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_837
timestamp 1669390400
transform 1 0 95088 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_845
timestamp 1669390400
transform 1 0 95984 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_849
timestamp 1669390400
transform 1 0 96432 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_851
timestamp 1669390400
transform 1 0 96656 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_854
timestamp 1669390400
transform 1 0 96992 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_870
timestamp 1669390400
transform 1 0 98784 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_872
timestamp 1669390400
transform 1 0 99008 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_879
timestamp 1669390400
transform 1 0 99792 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_911
timestamp 1669390400
transform 1 0 103376 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_919
timestamp 1669390400
transform 1 0 104272 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_925
timestamp 1669390400
transform 1 0 104944 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_989
timestamp 1669390400
transform 1 0 112112 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_993
timestamp 1669390400
transform 1 0 112560 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_996
timestamp 1669390400
transform 1 0 112896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_999
timestamp 1669390400
transform 1 0 113232 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1001
timestamp 1669390400
transform 1 0 113456 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1004
timestamp 1669390400
transform 1 0 113792 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1008
timestamp 1669390400
transform 1 0 114240 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1016
timestamp 1669390400
transform 1 0 115136 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1020
timestamp 1669390400
transform 1 0 115584 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1024
timestamp 1669390400
transform 1 0 116032 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1028
timestamp 1669390400
transform 1 0 116480 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1032
timestamp 1669390400
transform 1 0 116928 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1036
timestamp 1669390400
transform 1 0 117376 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1039
timestamp 1669390400
transform 1 0 117712 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1047
timestamp 1669390400
transform 1 0 118608 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1064
timestamp 1669390400
transform 1 0 120512 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1067
timestamp 1669390400
transform 1 0 120848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1083
timestamp 1669390400
transform 1 0 122640 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1087
timestamp 1669390400
transform 1 0 123088 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_1091
timestamp 1669390400
transform 1 0 123536 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1107
timestamp 1669390400
transform 1 0 125328 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1111
timestamp 1669390400
transform 1 0 125776 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1114
timestamp 1669390400
transform 1 0 126112 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1118
timestamp 1669390400
transform 1 0 126560 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1135
timestamp 1669390400
transform 1 0 128464 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1138
timestamp 1669390400
transform 1 0 128800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1173
timestamp 1669390400
transform 1 0 132720 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1177
timestamp 1669390400
transform 1 0 133168 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_1181
timestamp 1669390400
transform 1 0 133616 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1197
timestamp 1669390400
transform 1 0 135408 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1205
timestamp 1669390400
transform 1 0 136304 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_1209
timestamp 1669390400
transform 1 0 136752 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1241
timestamp 1669390400
transform 1 0 140336 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1249
timestamp 1669390400
transform 1 0 141232 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1256
timestamp 1669390400
transform 1 0 142016 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1264
timestamp 1669390400
transform 1 0 142912 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1272
timestamp 1669390400
transform 1 0 143808 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1276
timestamp 1669390400
transform 1 0 144256 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_1280
timestamp 1669390400
transform 1 0 144704 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1312
timestamp 1669390400
transform 1 0 148288 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1669390400
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1669390400
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1669390400
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1669390400
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1669390400
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1669390400
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1669390400
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_534
timestamp 1669390400
transform 1 0 61152 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_550
timestamp 1669390400
transform 1 0 62944 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_554
timestamp 1669390400
transform 1 0 63392 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_590
timestamp 1669390400
transform 1 0 67424 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_594
timestamp 1669390400
transform 1 0 67872 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_598
timestamp 1669390400
transform 1 0 68320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1669390400
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1669390400
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_669
timestamp 1669390400
transform 1 0 76272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1669390400
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_676
timestamp 1669390400
transform 1 0 77056 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_740
timestamp 1669390400
transform 1 0 84224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_744
timestamp 1669390400
transform 1 0 84672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_747
timestamp 1669390400
transform 1 0 85008 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_779
timestamp 1669390400
transform 1 0 88592 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_781
timestamp 1669390400
transform 1 0 88816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_784
timestamp 1669390400
transform 1 0 89152 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_818
timestamp 1669390400
transform 1 0 92960 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_882
timestamp 1669390400
transform 1 0 100128 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_886
timestamp 1669390400
transform 1 0 100576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_889
timestamp 1669390400
transform 1 0 100912 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_953
timestamp 1669390400
transform 1 0 108080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_957
timestamp 1669390400
transform 1 0 108528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_960
timestamp 1669390400
transform 1 0 108864 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1024
timestamp 1669390400
transform 1 0 116032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1028
timestamp 1669390400
transform 1 0 116480 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1031
timestamp 1669390400
transform 1 0 116816 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1039
timestamp 1669390400
transform 1 0 117712 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1045
timestamp 1669390400
transform 1 0 118384 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1062
timestamp 1669390400
transform 1 0 120288 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1066
timestamp 1669390400
transform 1 0 120736 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1070
timestamp 1669390400
transform 1 0 121184 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_1074
timestamp 1669390400
transform 1 0 121632 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1090
timestamp 1669390400
transform 1 0 123424 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1098
timestamp 1669390400
transform 1 0 124320 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_1102
timestamp 1669390400
transform 1 0 124768 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1118
timestamp 1669390400
transform 1 0 126560 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1122
timestamp 1669390400
transform 1 0 127008 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1130
timestamp 1669390400
transform 1 0 127904 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1166
timestamp 1669390400
transform 1 0 131936 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1170
timestamp 1669390400
transform 1 0 132384 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1173
timestamp 1669390400
transform 1 0 132720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1176
timestamp 1669390400
transform 1 0 133056 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1240
timestamp 1669390400
transform 1 0 140224 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1244
timestamp 1669390400
transform 1 0 140672 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1308
timestamp 1669390400
transform 1 0 147840 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1312
timestamp 1669390400
transform 1 0 148288 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1669390400
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1669390400
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1669390400
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1669390400
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1669390400
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1669390400
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_531
timestamp 1669390400
transform 1 0 60816 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_547
timestamp 1669390400
transform 1 0 62608 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_555
timestamp 1669390400
transform 1 0 63504 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_559
timestamp 1669390400
transform 1 0 63952 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_563
timestamp 1669390400
transform 1 0 64400 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1669390400
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_570
timestamp 1669390400
transform 1 0 65184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_586
timestamp 1669390400
transform 1 0 66976 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_590
timestamp 1669390400
transform 1 0 67424 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_622
timestamp 1669390400
transform 1 0 71008 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1669390400
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_641
timestamp 1669390400
transform 1 0 73136 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_705
timestamp 1669390400
transform 1 0 80304 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_709
timestamp 1669390400
transform 1 0 80752 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_712
timestamp 1669390400
transform 1 0 81088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_776
timestamp 1669390400
transform 1 0 88256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_780
timestamp 1669390400
transform 1 0 88704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_783
timestamp 1669390400
transform 1 0 89040 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_847
timestamp 1669390400
transform 1 0 96208 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_851
timestamp 1669390400
transform 1 0 96656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_854
timestamp 1669390400
transform 1 0 96992 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_918
timestamp 1669390400
transform 1 0 104160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_922
timestamp 1669390400
transform 1 0 104608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_925
timestamp 1669390400
transform 1 0 104944 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_989
timestamp 1669390400
transform 1 0 112112 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_993
timestamp 1669390400
transform 1 0 112560 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_996
timestamp 1669390400
transform 1 0 112896 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1060
timestamp 1669390400
transform 1 0 120064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1064
timestamp 1669390400
transform 1 0 120512 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_1067
timestamp 1669390400
transform 1 0 120848 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_1099
timestamp 1669390400
transform 1 0 124432 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_1115
timestamp 1669390400
transform 1 0 126224 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1123
timestamp 1669390400
transform 1 0 127120 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1127
timestamp 1669390400
transform 1 0 127568 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1135
timestamp 1669390400
transform 1 0 128464 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1138
timestamp 1669390400
transform 1 0 128800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1154
timestamp 1669390400
transform 1 0 130592 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1158
timestamp 1669390400
transform 1 0 131040 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_1162
timestamp 1669390400
transform 1 0 131488 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_1194
timestamp 1669390400
transform 1 0 135072 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1202
timestamp 1669390400
transform 1 0 135968 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1206
timestamp 1669390400
transform 1 0 136416 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1209
timestamp 1669390400
transform 1 0 136752 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1273
timestamp 1669390400
transform 1 0 143920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1277
timestamp 1669390400
transform 1 0 144368 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_1280
timestamp 1669390400
transform 1 0 144704 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1312
timestamp 1669390400
transform 1 0 148288 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1669390400
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1669390400
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1669390400
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1669390400
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1669390400
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1669390400
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1669390400
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1669390400
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_598
timestamp 1669390400
transform 1 0 68320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1669390400
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1669390400
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_669
timestamp 1669390400
transform 1 0 76272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1669390400
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_676
timestamp 1669390400
transform 1 0 77056 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_740
timestamp 1669390400
transform 1 0 84224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_744
timestamp 1669390400
transform 1 0 84672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_747
timestamp 1669390400
transform 1 0 85008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_811
timestamp 1669390400
transform 1 0 92176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_815
timestamp 1669390400
transform 1 0 92624 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_818
timestamp 1669390400
transform 1 0 92960 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_882
timestamp 1669390400
transform 1 0 100128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_886
timestamp 1669390400
transform 1 0 100576 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_889
timestamp 1669390400
transform 1 0 100912 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_953
timestamp 1669390400
transform 1 0 108080 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_957
timestamp 1669390400
transform 1 0 108528 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_960
timestamp 1669390400
transform 1 0 108864 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1024
timestamp 1669390400
transform 1 0 116032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1028
timestamp 1669390400
transform 1 0 116480 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1031
timestamp 1669390400
transform 1 0 116816 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1095
timestamp 1669390400
transform 1 0 123984 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1099
timestamp 1669390400
transform 1 0 124432 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_1102
timestamp 1669390400
transform 1 0 124768 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1134
timestamp 1669390400
transform 1 0 128352 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1136
timestamp 1669390400
transform 1 0 128576 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1139
timestamp 1669390400
transform 1 0 128912 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_1143
timestamp 1669390400
transform 1 0 129360 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_1159
timestamp 1669390400
transform 1 0 131152 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1167
timestamp 1669390400
transform 1 0 132048 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1173
timestamp 1669390400
transform 1 0 132720 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1237
timestamp 1669390400
transform 1 0 139888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1241
timestamp 1669390400
transform 1 0 140336 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1244
timestamp 1669390400
transform 1 0 140672 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1308
timestamp 1669390400
transform 1 0 147840 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1312
timestamp 1669390400
transform 1 0 148288 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1669390400
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1669390400
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1669390400
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1669390400
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1669390400
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_563
timestamp 1669390400
transform 1 0 64400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1669390400
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1669390400
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1669390400
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1669390400
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_641
timestamp 1669390400
transform 1 0 73136 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_705
timestamp 1669390400
transform 1 0 80304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_709
timestamp 1669390400
transform 1 0 80752 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_712
timestamp 1669390400
transform 1 0 81088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_776
timestamp 1669390400
transform 1 0 88256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_780
timestamp 1669390400
transform 1 0 88704 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_783
timestamp 1669390400
transform 1 0 89040 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_847
timestamp 1669390400
transform 1 0 96208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_851
timestamp 1669390400
transform 1 0 96656 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_854
timestamp 1669390400
transform 1 0 96992 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_918
timestamp 1669390400
transform 1 0 104160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_922
timestamp 1669390400
transform 1 0 104608 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_925
timestamp 1669390400
transform 1 0 104944 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_989
timestamp 1669390400
transform 1 0 112112 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_993
timestamp 1669390400
transform 1 0 112560 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_996
timestamp 1669390400
transform 1 0 112896 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1060
timestamp 1669390400
transform 1 0 120064 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1064
timestamp 1669390400
transform 1 0 120512 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1067
timestamp 1669390400
transform 1 0 120848 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1131
timestamp 1669390400
transform 1 0 128016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1135
timestamp 1669390400
transform 1 0 128464 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1138
timestamp 1669390400
transform 1 0 128800 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1202
timestamp 1669390400
transform 1 0 135968 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1206
timestamp 1669390400
transform 1 0 136416 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1209
timestamp 1669390400
transform 1 0 136752 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1273
timestamp 1669390400
transform 1 0 143920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1277
timestamp 1669390400
transform 1 0 144368 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_1280
timestamp 1669390400
transform 1 0 144704 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1312
timestamp 1669390400
transform 1 0 148288 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1669390400
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1669390400
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1669390400
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1669390400
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1669390400
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1669390400
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1669390400
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_598
timestamp 1669390400
transform 1 0 68320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1669390400
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_605
timestamp 1669390400
transform 1 0 69104 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_669
timestamp 1669390400
transform 1 0 76272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1669390400
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_676
timestamp 1669390400
transform 1 0 77056 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_740
timestamp 1669390400
transform 1 0 84224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_744
timestamp 1669390400
transform 1 0 84672 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_747
timestamp 1669390400
transform 1 0 85008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_811
timestamp 1669390400
transform 1 0 92176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_815
timestamp 1669390400
transform 1 0 92624 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_818
timestamp 1669390400
transform 1 0 92960 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_882
timestamp 1669390400
transform 1 0 100128 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_886
timestamp 1669390400
transform 1 0 100576 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_889
timestamp 1669390400
transform 1 0 100912 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_953
timestamp 1669390400
transform 1 0 108080 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_957
timestamp 1669390400
transform 1 0 108528 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_960
timestamp 1669390400
transform 1 0 108864 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1024
timestamp 1669390400
transform 1 0 116032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1028
timestamp 1669390400
transform 1 0 116480 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1031
timestamp 1669390400
transform 1 0 116816 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1095
timestamp 1669390400
transform 1 0 123984 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1099
timestamp 1669390400
transform 1 0 124432 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1102
timestamp 1669390400
transform 1 0 124768 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1166
timestamp 1669390400
transform 1 0 131936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1170
timestamp 1669390400
transform 1 0 132384 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1173
timestamp 1669390400
transform 1 0 132720 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1237
timestamp 1669390400
transform 1 0 139888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1241
timestamp 1669390400
transform 1 0 140336 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1244
timestamp 1669390400
transform 1 0 140672 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1308
timestamp 1669390400
transform 1 0 147840 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1312
timestamp 1669390400
transform 1 0 148288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1669390400
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1669390400
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1669390400
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1669390400
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1669390400
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_563
timestamp 1669390400
transform 1 0 64400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1669390400
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1669390400
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1669390400
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1669390400
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_641
timestamp 1669390400
transform 1 0 73136 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_705
timestamp 1669390400
transform 1 0 80304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_709
timestamp 1669390400
transform 1 0 80752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_712
timestamp 1669390400
transform 1 0 81088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_776
timestamp 1669390400
transform 1 0 88256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_780
timestamp 1669390400
transform 1 0 88704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_783
timestamp 1669390400
transform 1 0 89040 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_847
timestamp 1669390400
transform 1 0 96208 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_851
timestamp 1669390400
transform 1 0 96656 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_854
timestamp 1669390400
transform 1 0 96992 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_918
timestamp 1669390400
transform 1 0 104160 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_922
timestamp 1669390400
transform 1 0 104608 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_925
timestamp 1669390400
transform 1 0 104944 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_989
timestamp 1669390400
transform 1 0 112112 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_993
timestamp 1669390400
transform 1 0 112560 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_996
timestamp 1669390400
transform 1 0 112896 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1060
timestamp 1669390400
transform 1 0 120064 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1064
timestamp 1669390400
transform 1 0 120512 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1067
timestamp 1669390400
transform 1 0 120848 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1131
timestamp 1669390400
transform 1 0 128016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1135
timestamp 1669390400
transform 1 0 128464 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1138
timestamp 1669390400
transform 1 0 128800 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1202
timestamp 1669390400
transform 1 0 135968 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1206
timestamp 1669390400
transform 1 0 136416 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1209
timestamp 1669390400
transform 1 0 136752 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1273
timestamp 1669390400
transform 1 0 143920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1277
timestamp 1669390400
transform 1 0 144368 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_1280
timestamp 1669390400
transform 1 0 144704 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1312
timestamp 1669390400
transform 1 0 148288 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1669390400
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1669390400
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1669390400
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1669390400
transform 1 0 60368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1669390400
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1669390400
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_598
timestamp 1669390400
transform 1 0 68320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1669390400
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1669390400
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_669
timestamp 1669390400
transform 1 0 76272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1669390400
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_676
timestamp 1669390400
transform 1 0 77056 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_740
timestamp 1669390400
transform 1 0 84224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_744
timestamp 1669390400
transform 1 0 84672 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_747
timestamp 1669390400
transform 1 0 85008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_811
timestamp 1669390400
transform 1 0 92176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_815
timestamp 1669390400
transform 1 0 92624 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_818
timestamp 1669390400
transform 1 0 92960 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_882
timestamp 1669390400
transform 1 0 100128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_886
timestamp 1669390400
transform 1 0 100576 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_889
timestamp 1669390400
transform 1 0 100912 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_953
timestamp 1669390400
transform 1 0 108080 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_957
timestamp 1669390400
transform 1 0 108528 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_960
timestamp 1669390400
transform 1 0 108864 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1024
timestamp 1669390400
transform 1 0 116032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1028
timestamp 1669390400
transform 1 0 116480 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1031
timestamp 1669390400
transform 1 0 116816 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1095
timestamp 1669390400
transform 1 0 123984 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1099
timestamp 1669390400
transform 1 0 124432 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1102
timestamp 1669390400
transform 1 0 124768 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1166
timestamp 1669390400
transform 1 0 131936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1170
timestamp 1669390400
transform 1 0 132384 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1173
timestamp 1669390400
transform 1 0 132720 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1237
timestamp 1669390400
transform 1 0 139888 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1241
timestamp 1669390400
transform 1 0 140336 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1244
timestamp 1669390400
transform 1 0 140672 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1308
timestamp 1669390400
transform 1 0 147840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1312
timestamp 1669390400
transform 1 0 148288 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1669390400
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1669390400
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1669390400
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1669390400
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1669390400
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1669390400
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1669390400
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_563
timestamp 1669390400
transform 1 0 64400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1669390400
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1669390400
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1669390400
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1669390400
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_641
timestamp 1669390400
transform 1 0 73136 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_705
timestamp 1669390400
transform 1 0 80304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_709
timestamp 1669390400
transform 1 0 80752 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_712
timestamp 1669390400
transform 1 0 81088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_776
timestamp 1669390400
transform 1 0 88256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_780
timestamp 1669390400
transform 1 0 88704 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_783
timestamp 1669390400
transform 1 0 89040 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_847
timestamp 1669390400
transform 1 0 96208 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_851
timestamp 1669390400
transform 1 0 96656 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_854
timestamp 1669390400
transform 1 0 96992 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_918
timestamp 1669390400
transform 1 0 104160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_922
timestamp 1669390400
transform 1 0 104608 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_925
timestamp 1669390400
transform 1 0 104944 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_989
timestamp 1669390400
transform 1 0 112112 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_993
timestamp 1669390400
transform 1 0 112560 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_996
timestamp 1669390400
transform 1 0 112896 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1060
timestamp 1669390400
transform 1 0 120064 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1064
timestamp 1669390400
transform 1 0 120512 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1067
timestamp 1669390400
transform 1 0 120848 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1131
timestamp 1669390400
transform 1 0 128016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1135
timestamp 1669390400
transform 1 0 128464 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1138
timestamp 1669390400
transform 1 0 128800 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1202
timestamp 1669390400
transform 1 0 135968 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1206
timestamp 1669390400
transform 1 0 136416 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1209
timestamp 1669390400
transform 1 0 136752 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1273
timestamp 1669390400
transform 1 0 143920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1277
timestamp 1669390400
transform 1 0 144368 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_1280
timestamp 1669390400
transform 1 0 144704 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1312
timestamp 1669390400
transform 1 0 148288 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1669390400
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1669390400
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1669390400
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1669390400
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1669390400
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1669390400
transform 1 0 60368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1669390400
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1669390400
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1669390400
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1669390400
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1669390400
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_669
timestamp 1669390400
transform 1 0 76272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1669390400
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_676
timestamp 1669390400
transform 1 0 77056 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_740
timestamp 1669390400
transform 1 0 84224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_744
timestamp 1669390400
transform 1 0 84672 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_747
timestamp 1669390400
transform 1 0 85008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_811
timestamp 1669390400
transform 1 0 92176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_815
timestamp 1669390400
transform 1 0 92624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_818
timestamp 1669390400
transform 1 0 92960 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_882
timestamp 1669390400
transform 1 0 100128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_886
timestamp 1669390400
transform 1 0 100576 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_889
timestamp 1669390400
transform 1 0 100912 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_953
timestamp 1669390400
transform 1 0 108080 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_957
timestamp 1669390400
transform 1 0 108528 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_960
timestamp 1669390400
transform 1 0 108864 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1024
timestamp 1669390400
transform 1 0 116032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1028
timestamp 1669390400
transform 1 0 116480 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1031
timestamp 1669390400
transform 1 0 116816 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1095
timestamp 1669390400
transform 1 0 123984 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1099
timestamp 1669390400
transform 1 0 124432 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1102
timestamp 1669390400
transform 1 0 124768 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1166
timestamp 1669390400
transform 1 0 131936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1170
timestamp 1669390400
transform 1 0 132384 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1173
timestamp 1669390400
transform 1 0 132720 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1237
timestamp 1669390400
transform 1 0 139888 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1241
timestamp 1669390400
transform 1 0 140336 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1244
timestamp 1669390400
transform 1 0 140672 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1308
timestamp 1669390400
transform 1 0 147840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1312
timestamp 1669390400
transform 1 0 148288 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1669390400
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1669390400
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1669390400
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1669390400
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1669390400
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1669390400
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1669390400
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1669390400
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_641
timestamp 1669390400
transform 1 0 73136 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_705
timestamp 1669390400
transform 1 0 80304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_709
timestamp 1669390400
transform 1 0 80752 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_712
timestamp 1669390400
transform 1 0 81088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_776
timestamp 1669390400
transform 1 0 88256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_780
timestamp 1669390400
transform 1 0 88704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_783
timestamp 1669390400
transform 1 0 89040 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_847
timestamp 1669390400
transform 1 0 96208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_851
timestamp 1669390400
transform 1 0 96656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_854
timestamp 1669390400
transform 1 0 96992 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_918
timestamp 1669390400
transform 1 0 104160 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_922
timestamp 1669390400
transform 1 0 104608 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_925
timestamp 1669390400
transform 1 0 104944 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_989
timestamp 1669390400
transform 1 0 112112 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_993
timestamp 1669390400
transform 1 0 112560 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_996
timestamp 1669390400
transform 1 0 112896 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1060
timestamp 1669390400
transform 1 0 120064 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1064
timestamp 1669390400
transform 1 0 120512 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1067
timestamp 1669390400
transform 1 0 120848 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1131
timestamp 1669390400
transform 1 0 128016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1135
timestamp 1669390400
transform 1 0 128464 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1138
timestamp 1669390400
transform 1 0 128800 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1202
timestamp 1669390400
transform 1 0 135968 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1206
timestamp 1669390400
transform 1 0 136416 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1209
timestamp 1669390400
transform 1 0 136752 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1273
timestamp 1669390400
transform 1 0 143920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1277
timestamp 1669390400
transform 1 0 144368 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_1280
timestamp 1669390400
transform 1 0 144704 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1312
timestamp 1669390400
transform 1 0 148288 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1669390400
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1669390400
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1669390400
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1669390400
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1669390400
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1669390400
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1669390400
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_598
timestamp 1669390400
transform 1 0 68320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1669390400
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_605
timestamp 1669390400
transform 1 0 69104 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_669
timestamp 1669390400
transform 1 0 76272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_673
timestamp 1669390400
transform 1 0 76720 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_676
timestamp 1669390400
transform 1 0 77056 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_740
timestamp 1669390400
transform 1 0 84224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_744
timestamp 1669390400
transform 1 0 84672 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_747
timestamp 1669390400
transform 1 0 85008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_811
timestamp 1669390400
transform 1 0 92176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_815
timestamp 1669390400
transform 1 0 92624 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_818
timestamp 1669390400
transform 1 0 92960 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_882
timestamp 1669390400
transform 1 0 100128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_886
timestamp 1669390400
transform 1 0 100576 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_889
timestamp 1669390400
transform 1 0 100912 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_953
timestamp 1669390400
transform 1 0 108080 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_957
timestamp 1669390400
transform 1 0 108528 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_960
timestamp 1669390400
transform 1 0 108864 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1024
timestamp 1669390400
transform 1 0 116032 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1028
timestamp 1669390400
transform 1 0 116480 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1031
timestamp 1669390400
transform 1 0 116816 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1095
timestamp 1669390400
transform 1 0 123984 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1099
timestamp 1669390400
transform 1 0 124432 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1102
timestamp 1669390400
transform 1 0 124768 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1166
timestamp 1669390400
transform 1 0 131936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1170
timestamp 1669390400
transform 1 0 132384 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1173
timestamp 1669390400
transform 1 0 132720 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1237
timestamp 1669390400
transform 1 0 139888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1241
timestamp 1669390400
transform 1 0 140336 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1244
timestamp 1669390400
transform 1 0 140672 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1308
timestamp 1669390400
transform 1 0 147840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1312
timestamp 1669390400
transform 1 0 148288 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1669390400
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1669390400
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1669390400
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1669390400
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1669390400
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1669390400
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_563
timestamp 1669390400
transform 1 0 64400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1669390400
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1669390400
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_634
timestamp 1669390400
transform 1 0 72352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1669390400
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_641
timestamp 1669390400
transform 1 0 73136 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_705
timestamp 1669390400
transform 1 0 80304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_709
timestamp 1669390400
transform 1 0 80752 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_712
timestamp 1669390400
transform 1 0 81088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_776
timestamp 1669390400
transform 1 0 88256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_780
timestamp 1669390400
transform 1 0 88704 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_783
timestamp 1669390400
transform 1 0 89040 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_847
timestamp 1669390400
transform 1 0 96208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_851
timestamp 1669390400
transform 1 0 96656 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_854
timestamp 1669390400
transform 1 0 96992 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_918
timestamp 1669390400
transform 1 0 104160 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_922
timestamp 1669390400
transform 1 0 104608 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_925
timestamp 1669390400
transform 1 0 104944 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_989
timestamp 1669390400
transform 1 0 112112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_993
timestamp 1669390400
transform 1 0 112560 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_996
timestamp 1669390400
transform 1 0 112896 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1060
timestamp 1669390400
transform 1 0 120064 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1064
timestamp 1669390400
transform 1 0 120512 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1067
timestamp 1669390400
transform 1 0 120848 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1131
timestamp 1669390400
transform 1 0 128016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1135
timestamp 1669390400
transform 1 0 128464 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1138
timestamp 1669390400
transform 1 0 128800 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1202
timestamp 1669390400
transform 1 0 135968 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1206
timestamp 1669390400
transform 1 0 136416 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1209
timestamp 1669390400
transform 1 0 136752 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1273
timestamp 1669390400
transform 1 0 143920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1277
timestamp 1669390400
transform 1 0 144368 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_1280
timestamp 1669390400
transform 1 0 144704 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1312
timestamp 1669390400
transform 1 0 148288 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1669390400
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1669390400
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1669390400
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_527
timestamp 1669390400
transform 1 0 60368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1669390400
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1669390400
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_598
timestamp 1669390400
transform 1 0 68320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1669390400
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_605
timestamp 1669390400
transform 1 0 69104 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_669
timestamp 1669390400
transform 1 0 76272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_673
timestamp 1669390400
transform 1 0 76720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_676
timestamp 1669390400
transform 1 0 77056 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_740
timestamp 1669390400
transform 1 0 84224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_744
timestamp 1669390400
transform 1 0 84672 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_747
timestamp 1669390400
transform 1 0 85008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_811
timestamp 1669390400
transform 1 0 92176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_815
timestamp 1669390400
transform 1 0 92624 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_818
timestamp 1669390400
transform 1 0 92960 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_882
timestamp 1669390400
transform 1 0 100128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_886
timestamp 1669390400
transform 1 0 100576 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_889
timestamp 1669390400
transform 1 0 100912 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_953
timestamp 1669390400
transform 1 0 108080 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_957
timestamp 1669390400
transform 1 0 108528 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_960
timestamp 1669390400
transform 1 0 108864 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1024
timestamp 1669390400
transform 1 0 116032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1028
timestamp 1669390400
transform 1 0 116480 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1031
timestamp 1669390400
transform 1 0 116816 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1095
timestamp 1669390400
transform 1 0 123984 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1099
timestamp 1669390400
transform 1 0 124432 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1102
timestamp 1669390400
transform 1 0 124768 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1166
timestamp 1669390400
transform 1 0 131936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1170
timestamp 1669390400
transform 1 0 132384 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1173
timestamp 1669390400
transform 1 0 132720 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1237
timestamp 1669390400
transform 1 0 139888 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1241
timestamp 1669390400
transform 1 0 140336 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1244
timestamp 1669390400
transform 1 0 140672 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1308
timestamp 1669390400
transform 1 0 147840 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1312
timestamp 1669390400
transform 1 0 148288 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1669390400
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1669390400
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1669390400
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1669390400
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1669390400
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_563
timestamp 1669390400
transform 1 0 64400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1669390400
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1669390400
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1669390400
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1669390400
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_641
timestamp 1669390400
transform 1 0 73136 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_705
timestamp 1669390400
transform 1 0 80304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_709
timestamp 1669390400
transform 1 0 80752 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_712
timestamp 1669390400
transform 1 0 81088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_776
timestamp 1669390400
transform 1 0 88256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_780
timestamp 1669390400
transform 1 0 88704 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_783
timestamp 1669390400
transform 1 0 89040 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_847
timestamp 1669390400
transform 1 0 96208 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_851
timestamp 1669390400
transform 1 0 96656 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_854
timestamp 1669390400
transform 1 0 96992 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_918
timestamp 1669390400
transform 1 0 104160 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_922
timestamp 1669390400
transform 1 0 104608 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_925
timestamp 1669390400
transform 1 0 104944 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_989
timestamp 1669390400
transform 1 0 112112 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_993
timestamp 1669390400
transform 1 0 112560 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_996
timestamp 1669390400
transform 1 0 112896 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1060
timestamp 1669390400
transform 1 0 120064 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1064
timestamp 1669390400
transform 1 0 120512 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1067
timestamp 1669390400
transform 1 0 120848 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1131
timestamp 1669390400
transform 1 0 128016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1135
timestamp 1669390400
transform 1 0 128464 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1138
timestamp 1669390400
transform 1 0 128800 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1202
timestamp 1669390400
transform 1 0 135968 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1206
timestamp 1669390400
transform 1 0 136416 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1209
timestamp 1669390400
transform 1 0 136752 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1273
timestamp 1669390400
transform 1 0 143920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1277
timestamp 1669390400
transform 1 0 144368 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_1280
timestamp 1669390400
transform 1 0 144704 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1312
timestamp 1669390400
transform 1 0 148288 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1669390400
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1669390400
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1669390400
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_527
timestamp 1669390400
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1669390400
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1669390400
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_598
timestamp 1669390400
transform 1 0 68320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1669390400
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_605
timestamp 1669390400
transform 1 0 69104 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_669
timestamp 1669390400
transform 1 0 76272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_673
timestamp 1669390400
transform 1 0 76720 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_676
timestamp 1669390400
transform 1 0 77056 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_740
timestamp 1669390400
transform 1 0 84224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_744
timestamp 1669390400
transform 1 0 84672 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_747
timestamp 1669390400
transform 1 0 85008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_811
timestamp 1669390400
transform 1 0 92176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_815
timestamp 1669390400
transform 1 0 92624 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_818
timestamp 1669390400
transform 1 0 92960 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_882
timestamp 1669390400
transform 1 0 100128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_886
timestamp 1669390400
transform 1 0 100576 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_889
timestamp 1669390400
transform 1 0 100912 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_953
timestamp 1669390400
transform 1 0 108080 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_957
timestamp 1669390400
transform 1 0 108528 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_960
timestamp 1669390400
transform 1 0 108864 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1024
timestamp 1669390400
transform 1 0 116032 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1028
timestamp 1669390400
transform 1 0 116480 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1031
timestamp 1669390400
transform 1 0 116816 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1095
timestamp 1669390400
transform 1 0 123984 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1099
timestamp 1669390400
transform 1 0 124432 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1102
timestamp 1669390400
transform 1 0 124768 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1166
timestamp 1669390400
transform 1 0 131936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1170
timestamp 1669390400
transform 1 0 132384 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1173
timestamp 1669390400
transform 1 0 132720 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1237
timestamp 1669390400
transform 1 0 139888 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1241
timestamp 1669390400
transform 1 0 140336 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1244
timestamp 1669390400
transform 1 0 140672 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1308
timestamp 1669390400
transform 1 0 147840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1312
timestamp 1669390400
transform 1 0 148288 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1669390400
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1669390400
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1669390400
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1669390400
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1669390400
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_563
timestamp 1669390400
transform 1 0 64400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1669390400
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1669390400
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_634
timestamp 1669390400
transform 1 0 72352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1669390400
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_641
timestamp 1669390400
transform 1 0 73136 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_705
timestamp 1669390400
transform 1 0 80304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_709
timestamp 1669390400
transform 1 0 80752 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_712
timestamp 1669390400
transform 1 0 81088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_776
timestamp 1669390400
transform 1 0 88256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_780
timestamp 1669390400
transform 1 0 88704 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_783
timestamp 1669390400
transform 1 0 89040 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_847
timestamp 1669390400
transform 1 0 96208 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_851
timestamp 1669390400
transform 1 0 96656 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_854
timestamp 1669390400
transform 1 0 96992 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_918
timestamp 1669390400
transform 1 0 104160 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_922
timestamp 1669390400
transform 1 0 104608 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_925
timestamp 1669390400
transform 1 0 104944 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_989
timestamp 1669390400
transform 1 0 112112 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_993
timestamp 1669390400
transform 1 0 112560 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_996
timestamp 1669390400
transform 1 0 112896 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1060
timestamp 1669390400
transform 1 0 120064 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1064
timestamp 1669390400
transform 1 0 120512 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1067
timestamp 1669390400
transform 1 0 120848 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1131
timestamp 1669390400
transform 1 0 128016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1135
timestamp 1669390400
transform 1 0 128464 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1138
timestamp 1669390400
transform 1 0 128800 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1202
timestamp 1669390400
transform 1 0 135968 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1206
timestamp 1669390400
transform 1 0 136416 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1209
timestamp 1669390400
transform 1 0 136752 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1273
timestamp 1669390400
transform 1 0 143920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1277
timestamp 1669390400
transform 1 0 144368 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_1280
timestamp 1669390400
transform 1 0 144704 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1312
timestamp 1669390400
transform 1 0 148288 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1669390400
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1669390400
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1669390400
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_527
timestamp 1669390400
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1669390400
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1669390400
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_598
timestamp 1669390400
transform 1 0 68320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1669390400
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_605
timestamp 1669390400
transform 1 0 69104 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_669
timestamp 1669390400
transform 1 0 76272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_673
timestamp 1669390400
transform 1 0 76720 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_676
timestamp 1669390400
transform 1 0 77056 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_740
timestamp 1669390400
transform 1 0 84224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_744
timestamp 1669390400
transform 1 0 84672 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_747
timestamp 1669390400
transform 1 0 85008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_811
timestamp 1669390400
transform 1 0 92176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_815
timestamp 1669390400
transform 1 0 92624 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_818
timestamp 1669390400
transform 1 0 92960 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_882
timestamp 1669390400
transform 1 0 100128 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_886
timestamp 1669390400
transform 1 0 100576 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_889
timestamp 1669390400
transform 1 0 100912 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_953
timestamp 1669390400
transform 1 0 108080 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_957
timestamp 1669390400
transform 1 0 108528 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_960
timestamp 1669390400
transform 1 0 108864 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1024
timestamp 1669390400
transform 1 0 116032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1028
timestamp 1669390400
transform 1 0 116480 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1031
timestamp 1669390400
transform 1 0 116816 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1095
timestamp 1669390400
transform 1 0 123984 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1099
timestamp 1669390400
transform 1 0 124432 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1102
timestamp 1669390400
transform 1 0 124768 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1166
timestamp 1669390400
transform 1 0 131936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1170
timestamp 1669390400
transform 1 0 132384 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1173
timestamp 1669390400
transform 1 0 132720 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1237
timestamp 1669390400
transform 1 0 139888 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1241
timestamp 1669390400
transform 1 0 140336 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1244
timestamp 1669390400
transform 1 0 140672 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1308
timestamp 1669390400
transform 1 0 147840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1312
timestamp 1669390400
transform 1 0 148288 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1669390400
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1669390400
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1669390400
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1669390400
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_563
timestamp 1669390400
transform 1 0 64400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1669390400
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1669390400
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_634
timestamp 1669390400
transform 1 0 72352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1669390400
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_641
timestamp 1669390400
transform 1 0 73136 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_705
timestamp 1669390400
transform 1 0 80304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_709
timestamp 1669390400
transform 1 0 80752 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_712
timestamp 1669390400
transform 1 0 81088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_776
timestamp 1669390400
transform 1 0 88256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_780
timestamp 1669390400
transform 1 0 88704 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_783
timestamp 1669390400
transform 1 0 89040 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_847
timestamp 1669390400
transform 1 0 96208 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_851
timestamp 1669390400
transform 1 0 96656 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_854
timestamp 1669390400
transform 1 0 96992 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_918
timestamp 1669390400
transform 1 0 104160 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_922
timestamp 1669390400
transform 1 0 104608 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_925
timestamp 1669390400
transform 1 0 104944 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_989
timestamp 1669390400
transform 1 0 112112 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_993
timestamp 1669390400
transform 1 0 112560 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_996
timestamp 1669390400
transform 1 0 112896 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1060
timestamp 1669390400
transform 1 0 120064 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1064
timestamp 1669390400
transform 1 0 120512 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1067
timestamp 1669390400
transform 1 0 120848 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1131
timestamp 1669390400
transform 1 0 128016 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1135
timestamp 1669390400
transform 1 0 128464 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1138
timestamp 1669390400
transform 1 0 128800 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1202
timestamp 1669390400
transform 1 0 135968 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1206
timestamp 1669390400
transform 1 0 136416 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1209
timestamp 1669390400
transform 1 0 136752 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1273
timestamp 1669390400
transform 1 0 143920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1277
timestamp 1669390400
transform 1 0 144368 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_1280
timestamp 1669390400
transform 1 0 144704 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1312
timestamp 1669390400
transform 1 0 148288 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1669390400
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1669390400
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1669390400
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1669390400
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1669390400
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1669390400
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_527
timestamp 1669390400
transform 1 0 60368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1669390400
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1669390400
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_598
timestamp 1669390400
transform 1 0 68320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1669390400
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_605
timestamp 1669390400
transform 1 0 69104 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_669
timestamp 1669390400
transform 1 0 76272 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1669390400
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_676
timestamp 1669390400
transform 1 0 77056 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_740
timestamp 1669390400
transform 1 0 84224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_744
timestamp 1669390400
transform 1 0 84672 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_747
timestamp 1669390400
transform 1 0 85008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_811
timestamp 1669390400
transform 1 0 92176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_815
timestamp 1669390400
transform 1 0 92624 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_818
timestamp 1669390400
transform 1 0 92960 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_882
timestamp 1669390400
transform 1 0 100128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_886
timestamp 1669390400
transform 1 0 100576 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_889
timestamp 1669390400
transform 1 0 100912 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_953
timestamp 1669390400
transform 1 0 108080 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_957
timestamp 1669390400
transform 1 0 108528 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_960
timestamp 1669390400
transform 1 0 108864 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1024
timestamp 1669390400
transform 1 0 116032 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1028
timestamp 1669390400
transform 1 0 116480 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1031
timestamp 1669390400
transform 1 0 116816 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1095
timestamp 1669390400
transform 1 0 123984 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1099
timestamp 1669390400
transform 1 0 124432 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1102
timestamp 1669390400
transform 1 0 124768 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1166
timestamp 1669390400
transform 1 0 131936 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1170
timestamp 1669390400
transform 1 0 132384 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1173
timestamp 1669390400
transform 1 0 132720 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1237
timestamp 1669390400
transform 1 0 139888 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1241
timestamp 1669390400
transform 1 0 140336 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1244
timestamp 1669390400
transform 1 0 140672 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1308
timestamp 1669390400
transform 1 0 147840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1312
timestamp 1669390400
transform 1 0 148288 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1669390400
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1669390400
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1669390400
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1669390400
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_563
timestamp 1669390400
transform 1 0 64400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1669390400
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1669390400
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1669390400
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1669390400
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_641
timestamp 1669390400
transform 1 0 73136 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_705
timestamp 1669390400
transform 1 0 80304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_709
timestamp 1669390400
transform 1 0 80752 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_712
timestamp 1669390400
transform 1 0 81088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_776
timestamp 1669390400
transform 1 0 88256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_780
timestamp 1669390400
transform 1 0 88704 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_783
timestamp 1669390400
transform 1 0 89040 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_847
timestamp 1669390400
transform 1 0 96208 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_851
timestamp 1669390400
transform 1 0 96656 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_854
timestamp 1669390400
transform 1 0 96992 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_918
timestamp 1669390400
transform 1 0 104160 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_922
timestamp 1669390400
transform 1 0 104608 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_925
timestamp 1669390400
transform 1 0 104944 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_989
timestamp 1669390400
transform 1 0 112112 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_993
timestamp 1669390400
transform 1 0 112560 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_996
timestamp 1669390400
transform 1 0 112896 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1060
timestamp 1669390400
transform 1 0 120064 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1064
timestamp 1669390400
transform 1 0 120512 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1067
timestamp 1669390400
transform 1 0 120848 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1131
timestamp 1669390400
transform 1 0 128016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1135
timestamp 1669390400
transform 1 0 128464 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1138
timestamp 1669390400
transform 1 0 128800 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1202
timestamp 1669390400
transform 1 0 135968 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1206
timestamp 1669390400
transform 1 0 136416 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1209
timestamp 1669390400
transform 1 0 136752 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1273
timestamp 1669390400
transform 1 0 143920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1277
timestamp 1669390400
transform 1 0 144368 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_1280
timestamp 1669390400
transform 1 0 144704 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1312
timestamp 1669390400
transform 1 0 148288 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1669390400
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1669390400
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1669390400
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1669390400
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_527
timestamp 1669390400
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1669390400
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1669390400
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_598
timestamp 1669390400
transform 1 0 68320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1669390400
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605
timestamp 1669390400
transform 1 0 69104 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_669
timestamp 1669390400
transform 1 0 76272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1669390400
transform 1 0 76720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_676
timestamp 1669390400
transform 1 0 77056 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_740
timestamp 1669390400
transform 1 0 84224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_744
timestamp 1669390400
transform 1 0 84672 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_747
timestamp 1669390400
transform 1 0 85008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_811
timestamp 1669390400
transform 1 0 92176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_815
timestamp 1669390400
transform 1 0 92624 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_818
timestamp 1669390400
transform 1 0 92960 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_882
timestamp 1669390400
transform 1 0 100128 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_886
timestamp 1669390400
transform 1 0 100576 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_889
timestamp 1669390400
transform 1 0 100912 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_953
timestamp 1669390400
transform 1 0 108080 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_957
timestamp 1669390400
transform 1 0 108528 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_960
timestamp 1669390400
transform 1 0 108864 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1024
timestamp 1669390400
transform 1 0 116032 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1028
timestamp 1669390400
transform 1 0 116480 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1031
timestamp 1669390400
transform 1 0 116816 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1095
timestamp 1669390400
transform 1 0 123984 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1099
timestamp 1669390400
transform 1 0 124432 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1102
timestamp 1669390400
transform 1 0 124768 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1166
timestamp 1669390400
transform 1 0 131936 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1170
timestamp 1669390400
transform 1 0 132384 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1173
timestamp 1669390400
transform 1 0 132720 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1237
timestamp 1669390400
transform 1 0 139888 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1241
timestamp 1669390400
transform 1 0 140336 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1244
timestamp 1669390400
transform 1 0 140672 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1308
timestamp 1669390400
transform 1 0 147840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1312
timestamp 1669390400
transform 1 0 148288 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1669390400
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1669390400
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1669390400
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_563
timestamp 1669390400
transform 1 0 64400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1669390400
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1669390400
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1669390400
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1669390400
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_641
timestamp 1669390400
transform 1 0 73136 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_705
timestamp 1669390400
transform 1 0 80304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_709
timestamp 1669390400
transform 1 0 80752 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_712
timestamp 1669390400
transform 1 0 81088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_776
timestamp 1669390400
transform 1 0 88256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_780
timestamp 1669390400
transform 1 0 88704 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_783
timestamp 1669390400
transform 1 0 89040 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_847
timestamp 1669390400
transform 1 0 96208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_851
timestamp 1669390400
transform 1 0 96656 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_854
timestamp 1669390400
transform 1 0 96992 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_918
timestamp 1669390400
transform 1 0 104160 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_922
timestamp 1669390400
transform 1 0 104608 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_925
timestamp 1669390400
transform 1 0 104944 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_989
timestamp 1669390400
transform 1 0 112112 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_993
timestamp 1669390400
transform 1 0 112560 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_996
timestamp 1669390400
transform 1 0 112896 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1060
timestamp 1669390400
transform 1 0 120064 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1064
timestamp 1669390400
transform 1 0 120512 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1067
timestamp 1669390400
transform 1 0 120848 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1131
timestamp 1669390400
transform 1 0 128016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1135
timestamp 1669390400
transform 1 0 128464 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1138
timestamp 1669390400
transform 1 0 128800 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1202
timestamp 1669390400
transform 1 0 135968 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1206
timestamp 1669390400
transform 1 0 136416 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1209
timestamp 1669390400
transform 1 0 136752 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1273
timestamp 1669390400
transform 1 0 143920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1277
timestamp 1669390400
transform 1 0 144368 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_1280
timestamp 1669390400
transform 1 0 144704 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1312
timestamp 1669390400
transform 1 0 148288 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1669390400
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1669390400
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_527
timestamp 1669390400
transform 1 0 60368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1669390400
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1669390400
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1669390400
transform 1 0 68320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1669390400
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1669390400
transform 1 0 69104 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_669
timestamp 1669390400
transform 1 0 76272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1669390400
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_676
timestamp 1669390400
transform 1 0 77056 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_740
timestamp 1669390400
transform 1 0 84224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_744
timestamp 1669390400
transform 1 0 84672 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_747
timestamp 1669390400
transform 1 0 85008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_811
timestamp 1669390400
transform 1 0 92176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_815
timestamp 1669390400
transform 1 0 92624 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_818
timestamp 1669390400
transform 1 0 92960 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_882
timestamp 1669390400
transform 1 0 100128 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_886
timestamp 1669390400
transform 1 0 100576 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_889
timestamp 1669390400
transform 1 0 100912 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_953
timestamp 1669390400
transform 1 0 108080 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_957
timestamp 1669390400
transform 1 0 108528 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_960
timestamp 1669390400
transform 1 0 108864 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1024
timestamp 1669390400
transform 1 0 116032 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1028
timestamp 1669390400
transform 1 0 116480 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1031
timestamp 1669390400
transform 1 0 116816 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1095
timestamp 1669390400
transform 1 0 123984 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1099
timestamp 1669390400
transform 1 0 124432 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1102
timestamp 1669390400
transform 1 0 124768 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1166
timestamp 1669390400
transform 1 0 131936 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1170
timestamp 1669390400
transform 1 0 132384 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1173
timestamp 1669390400
transform 1 0 132720 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1237
timestamp 1669390400
transform 1 0 139888 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1241
timestamp 1669390400
transform 1 0 140336 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1244
timestamp 1669390400
transform 1 0 140672 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1308
timestamp 1669390400
transform 1 0 147840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1312
timestamp 1669390400
transform 1 0 148288 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1669390400
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1669390400
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1669390400
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1669390400
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_563
timestamp 1669390400
transform 1 0 64400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1669390400
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1669390400
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1669390400
transform 1 0 72352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1669390400
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_641
timestamp 1669390400
transform 1 0 73136 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_705
timestamp 1669390400
transform 1 0 80304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_709
timestamp 1669390400
transform 1 0 80752 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_712
timestamp 1669390400
transform 1 0 81088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_776
timestamp 1669390400
transform 1 0 88256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_780
timestamp 1669390400
transform 1 0 88704 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_783
timestamp 1669390400
transform 1 0 89040 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_847
timestamp 1669390400
transform 1 0 96208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_851
timestamp 1669390400
transform 1 0 96656 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_854
timestamp 1669390400
transform 1 0 96992 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_918
timestamp 1669390400
transform 1 0 104160 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_922
timestamp 1669390400
transform 1 0 104608 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_925
timestamp 1669390400
transform 1 0 104944 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_989
timestamp 1669390400
transform 1 0 112112 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_993
timestamp 1669390400
transform 1 0 112560 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_996
timestamp 1669390400
transform 1 0 112896 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1060
timestamp 1669390400
transform 1 0 120064 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1064
timestamp 1669390400
transform 1 0 120512 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1067
timestamp 1669390400
transform 1 0 120848 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1131
timestamp 1669390400
transform 1 0 128016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1135
timestamp 1669390400
transform 1 0 128464 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1138
timestamp 1669390400
transform 1 0 128800 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1202
timestamp 1669390400
transform 1 0 135968 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1206
timestamp 1669390400
transform 1 0 136416 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1209
timestamp 1669390400
transform 1 0 136752 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1273
timestamp 1669390400
transform 1 0 143920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1277
timestamp 1669390400
transform 1 0 144368 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_1280
timestamp 1669390400
transform 1 0 144704 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1312
timestamp 1669390400
transform 1 0 148288 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1669390400
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1669390400
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1669390400
transform 1 0 60368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1669390400
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1669390400
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1669390400
transform 1 0 68320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1669390400
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1669390400
transform 1 0 69104 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_669
timestamp 1669390400
transform 1 0 76272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1669390400
transform 1 0 76720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_676
timestamp 1669390400
transform 1 0 77056 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_740
timestamp 1669390400
transform 1 0 84224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_744
timestamp 1669390400
transform 1 0 84672 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_747
timestamp 1669390400
transform 1 0 85008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_811
timestamp 1669390400
transform 1 0 92176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_815
timestamp 1669390400
transform 1 0 92624 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_818
timestamp 1669390400
transform 1 0 92960 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_882
timestamp 1669390400
transform 1 0 100128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_886
timestamp 1669390400
transform 1 0 100576 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_889
timestamp 1669390400
transform 1 0 100912 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_953
timestamp 1669390400
transform 1 0 108080 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_957
timestamp 1669390400
transform 1 0 108528 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_960
timestamp 1669390400
transform 1 0 108864 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1024
timestamp 1669390400
transform 1 0 116032 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1028
timestamp 1669390400
transform 1 0 116480 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1031
timestamp 1669390400
transform 1 0 116816 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1095
timestamp 1669390400
transform 1 0 123984 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1099
timestamp 1669390400
transform 1 0 124432 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1102
timestamp 1669390400
transform 1 0 124768 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1166
timestamp 1669390400
transform 1 0 131936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1170
timestamp 1669390400
transform 1 0 132384 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1173
timestamp 1669390400
transform 1 0 132720 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1237
timestamp 1669390400
transform 1 0 139888 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1241
timestamp 1669390400
transform 1 0 140336 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1244
timestamp 1669390400
transform 1 0 140672 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1308
timestamp 1669390400
transform 1 0 147840 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1312
timestamp 1669390400
transform 1 0 148288 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1669390400
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1669390400
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1669390400
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1669390400
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1669390400
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1669390400
transform 1 0 64400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1669390400
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1669390400
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1669390400
transform 1 0 72352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1669390400
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_641
timestamp 1669390400
transform 1 0 73136 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_705
timestamp 1669390400
transform 1 0 80304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_709
timestamp 1669390400
transform 1 0 80752 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_712
timestamp 1669390400
transform 1 0 81088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_776
timestamp 1669390400
transform 1 0 88256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_780
timestamp 1669390400
transform 1 0 88704 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_783
timestamp 1669390400
transform 1 0 89040 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_847
timestamp 1669390400
transform 1 0 96208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_851
timestamp 1669390400
transform 1 0 96656 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_854
timestamp 1669390400
transform 1 0 96992 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_918
timestamp 1669390400
transform 1 0 104160 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_922
timestamp 1669390400
transform 1 0 104608 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_925
timestamp 1669390400
transform 1 0 104944 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_989
timestamp 1669390400
transform 1 0 112112 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_993
timestamp 1669390400
transform 1 0 112560 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_996
timestamp 1669390400
transform 1 0 112896 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1060
timestamp 1669390400
transform 1 0 120064 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1064
timestamp 1669390400
transform 1 0 120512 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1067
timestamp 1669390400
transform 1 0 120848 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1131
timestamp 1669390400
transform 1 0 128016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1135
timestamp 1669390400
transform 1 0 128464 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1138
timestamp 1669390400
transform 1 0 128800 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1202
timestamp 1669390400
transform 1 0 135968 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1206
timestamp 1669390400
transform 1 0 136416 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1209
timestamp 1669390400
transform 1 0 136752 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1273
timestamp 1669390400
transform 1 0 143920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1277
timestamp 1669390400
transform 1 0 144368 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_1280
timestamp 1669390400
transform 1 0 144704 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1312
timestamp 1669390400
transform 1 0 148288 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1669390400
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1669390400
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1669390400
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1669390400
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1669390400
transform 1 0 60368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1669390400
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1669390400
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1669390400
transform 1 0 68320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1669390400
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1669390400
transform 1 0 69104 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_669
timestamp 1669390400
transform 1 0 76272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1669390400
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_676
timestamp 1669390400
transform 1 0 77056 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_740
timestamp 1669390400
transform 1 0 84224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_744
timestamp 1669390400
transform 1 0 84672 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_747
timestamp 1669390400
transform 1 0 85008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_811
timestamp 1669390400
transform 1 0 92176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_815
timestamp 1669390400
transform 1 0 92624 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_818
timestamp 1669390400
transform 1 0 92960 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_882
timestamp 1669390400
transform 1 0 100128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_886
timestamp 1669390400
transform 1 0 100576 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_889
timestamp 1669390400
transform 1 0 100912 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_953
timestamp 1669390400
transform 1 0 108080 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_957
timestamp 1669390400
transform 1 0 108528 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_960
timestamp 1669390400
transform 1 0 108864 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1024
timestamp 1669390400
transform 1 0 116032 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1028
timestamp 1669390400
transform 1 0 116480 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1031
timestamp 1669390400
transform 1 0 116816 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1095
timestamp 1669390400
transform 1 0 123984 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1099
timestamp 1669390400
transform 1 0 124432 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1102
timestamp 1669390400
transform 1 0 124768 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1166
timestamp 1669390400
transform 1 0 131936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1170
timestamp 1669390400
transform 1 0 132384 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1173
timestamp 1669390400
transform 1 0 132720 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1237
timestamp 1669390400
transform 1 0 139888 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1241
timestamp 1669390400
transform 1 0 140336 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1244
timestamp 1669390400
transform 1 0 140672 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1308
timestamp 1669390400
transform 1 0 147840 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1312
timestamp 1669390400
transform 1 0 148288 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1669390400
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1669390400
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1669390400
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1669390400
transform 1 0 64400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1669390400
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1669390400
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1669390400
transform 1 0 72352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1669390400
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_641
timestamp 1669390400
transform 1 0 73136 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_705
timestamp 1669390400
transform 1 0 80304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_709
timestamp 1669390400
transform 1 0 80752 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_712
timestamp 1669390400
transform 1 0 81088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_776
timestamp 1669390400
transform 1 0 88256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_780
timestamp 1669390400
transform 1 0 88704 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_783
timestamp 1669390400
transform 1 0 89040 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_847
timestamp 1669390400
transform 1 0 96208 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_851
timestamp 1669390400
transform 1 0 96656 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_854
timestamp 1669390400
transform 1 0 96992 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_918
timestamp 1669390400
transform 1 0 104160 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_922
timestamp 1669390400
transform 1 0 104608 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_925
timestamp 1669390400
transform 1 0 104944 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_989
timestamp 1669390400
transform 1 0 112112 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_993
timestamp 1669390400
transform 1 0 112560 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_996
timestamp 1669390400
transform 1 0 112896 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1060
timestamp 1669390400
transform 1 0 120064 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1064
timestamp 1669390400
transform 1 0 120512 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1067
timestamp 1669390400
transform 1 0 120848 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1131
timestamp 1669390400
transform 1 0 128016 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1135
timestamp 1669390400
transform 1 0 128464 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1138
timestamp 1669390400
transform 1 0 128800 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1202
timestamp 1669390400
transform 1 0 135968 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1206
timestamp 1669390400
transform 1 0 136416 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1209
timestamp 1669390400
transform 1 0 136752 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1273
timestamp 1669390400
transform 1 0 143920 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1277
timestamp 1669390400
transform 1 0 144368 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_1280
timestamp 1669390400
transform 1 0 144704 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1312
timestamp 1669390400
transform 1 0 148288 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1669390400
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1669390400
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1669390400
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1669390400
transform 1 0 60368 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1669390400
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1669390400
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1669390400
transform 1 0 68320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1669390400
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_605
timestamp 1669390400
transform 1 0 69104 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_669
timestamp 1669390400
transform 1 0 76272 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1669390400
transform 1 0 76720 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_676
timestamp 1669390400
transform 1 0 77056 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_740
timestamp 1669390400
transform 1 0 84224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_744
timestamp 1669390400
transform 1 0 84672 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_747
timestamp 1669390400
transform 1 0 85008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_811
timestamp 1669390400
transform 1 0 92176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_815
timestamp 1669390400
transform 1 0 92624 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_818
timestamp 1669390400
transform 1 0 92960 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_882
timestamp 1669390400
transform 1 0 100128 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_886
timestamp 1669390400
transform 1 0 100576 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_889
timestamp 1669390400
transform 1 0 100912 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_953
timestamp 1669390400
transform 1 0 108080 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_957
timestamp 1669390400
transform 1 0 108528 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_960
timestamp 1669390400
transform 1 0 108864 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1024
timestamp 1669390400
transform 1 0 116032 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1028
timestamp 1669390400
transform 1 0 116480 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1031
timestamp 1669390400
transform 1 0 116816 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1095
timestamp 1669390400
transform 1 0 123984 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1099
timestamp 1669390400
transform 1 0 124432 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1102
timestamp 1669390400
transform 1 0 124768 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1166
timestamp 1669390400
transform 1 0 131936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1170
timestamp 1669390400
transform 1 0 132384 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1173
timestamp 1669390400
transform 1 0 132720 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1237
timestamp 1669390400
transform 1 0 139888 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1241
timestamp 1669390400
transform 1 0 140336 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1244
timestamp 1669390400
transform 1 0 140672 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1308
timestamp 1669390400
transform 1 0 147840 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1312
timestamp 1669390400
transform 1 0 148288 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1669390400
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1669390400
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1669390400
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1669390400
transform 1 0 64400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1669390400
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1669390400
transform 1 0 65184 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1669390400
transform 1 0 72352 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1669390400
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_641
timestamp 1669390400
transform 1 0 73136 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_705
timestamp 1669390400
transform 1 0 80304 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_709
timestamp 1669390400
transform 1 0 80752 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_712
timestamp 1669390400
transform 1 0 81088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_776
timestamp 1669390400
transform 1 0 88256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_780
timestamp 1669390400
transform 1 0 88704 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_783
timestamp 1669390400
transform 1 0 89040 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_847
timestamp 1669390400
transform 1 0 96208 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_851
timestamp 1669390400
transform 1 0 96656 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_854
timestamp 1669390400
transform 1 0 96992 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_918
timestamp 1669390400
transform 1 0 104160 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_922
timestamp 1669390400
transform 1 0 104608 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_925
timestamp 1669390400
transform 1 0 104944 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_989
timestamp 1669390400
transform 1 0 112112 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_993
timestamp 1669390400
transform 1 0 112560 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_996
timestamp 1669390400
transform 1 0 112896 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1060
timestamp 1669390400
transform 1 0 120064 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1064
timestamp 1669390400
transform 1 0 120512 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1067
timestamp 1669390400
transform 1 0 120848 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1131
timestamp 1669390400
transform 1 0 128016 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1135
timestamp 1669390400
transform 1 0 128464 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1138
timestamp 1669390400
transform 1 0 128800 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1202
timestamp 1669390400
transform 1 0 135968 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1206
timestamp 1669390400
transform 1 0 136416 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1209
timestamp 1669390400
transform 1 0 136752 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1273
timestamp 1669390400
transform 1 0 143920 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1277
timestamp 1669390400
transform 1 0 144368 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_1280
timestamp 1669390400
transform 1 0 144704 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1312
timestamp 1669390400
transform 1 0 148288 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1669390400
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1669390400
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_424
timestamp 1669390400
transform 1 0 48832 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_427
timestamp 1669390400
transform 1 0 49168 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_459
timestamp 1669390400
transform 1 0 52752 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1669390400
transform 1 0 60368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1669390400
transform 1 0 60816 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_534
timestamp 1669390400
transform 1 0 61152 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_566
timestamp 1669390400
transform 1 0 64736 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_569
timestamp 1669390400
transform 1 0 65072 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_601
timestamp 1669390400
transform 1 0 68656 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1669390400
transform 1 0 69104 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_669
timestamp 1669390400
transform 1 0 76272 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1669390400
transform 1 0 76720 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_676
timestamp 1669390400
transform 1 0 77056 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_740
timestamp 1669390400
transform 1 0 84224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_744
timestamp 1669390400
transform 1 0 84672 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_747
timestamp 1669390400
transform 1 0 85008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_811
timestamp 1669390400
transform 1 0 92176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_815
timestamp 1669390400
transform 1 0 92624 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_818
timestamp 1669390400
transform 1 0 92960 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_882
timestamp 1669390400
transform 1 0 100128 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_886
timestamp 1669390400
transform 1 0 100576 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_889
timestamp 1669390400
transform 1 0 100912 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_953
timestamp 1669390400
transform 1 0 108080 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_957
timestamp 1669390400
transform 1 0 108528 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_960
timestamp 1669390400
transform 1 0 108864 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1024
timestamp 1669390400
transform 1 0 116032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1028
timestamp 1669390400
transform 1 0 116480 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1031
timestamp 1669390400
transform 1 0 116816 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1095
timestamp 1669390400
transform 1 0 123984 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1099
timestamp 1669390400
transform 1 0 124432 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1102
timestamp 1669390400
transform 1 0 124768 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1166
timestamp 1669390400
transform 1 0 131936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1170
timestamp 1669390400
transform 1 0 132384 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1173
timestamp 1669390400
transform 1 0 132720 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1237
timestamp 1669390400
transform 1 0 139888 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1241
timestamp 1669390400
transform 1 0 140336 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1244
timestamp 1669390400
transform 1 0 140672 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1308
timestamp 1669390400
transform 1 0 147840 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1312
timestamp 1669390400
transform 1 0 148288 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1669390400
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_318
timestamp 1669390400
transform 1 0 36960 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_326
timestamp 1669390400
transform 1 0 37856 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_330
timestamp 1669390400
transform 1 0 38304 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_333
timestamp 1669390400
transform 1 0 38640 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_337
timestamp 1669390400
transform 1 0 39088 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_341
timestamp 1669390400
transform 1 0 39536 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_345
timestamp 1669390400
transform 1 0 39984 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_348
timestamp 1669390400
transform 1 0 40320 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_350
timestamp 1669390400
transform 1 0 40544 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_353
timestamp 1669390400
transform 1 0 40880 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_360
timestamp 1669390400
transform 1 0 41664 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_364
timestamp 1669390400
transform 1 0 42112 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_396
timestamp 1669390400
transform 1 0 45696 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_400
timestamp 1669390400
transform 1 0 46144 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_402
timestamp 1669390400
transform 1 0 46368 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_405
timestamp 1669390400
transform 1 0 46704 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_409
timestamp 1669390400
transform 1 0 47152 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_415
timestamp 1669390400
transform 1 0 47824 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_419
timestamp 1669390400
transform 1 0 48272 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_423
timestamp 1669390400
transform 1 0 48720 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1669390400
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_431
timestamp 1669390400
transform 1 0 49616 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_435
timestamp 1669390400
transform 1 0 50064 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_437
timestamp 1669390400
transform 1 0 50288 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_440
timestamp 1669390400
transform 1 0 50624 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_444
timestamp 1669390400
transform 1 0 51072 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_448
timestamp 1669390400
transform 1 0 51520 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_458
timestamp 1669390400
transform 1 0 52640 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_490
timestamp 1669390400
transform 1 0 56224 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_494
timestamp 1669390400
transform 1 0 56672 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1669390400
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_531
timestamp 1669390400
transform 1 0 60816 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_539
timestamp 1669390400
transform 1 0 61712 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_542
timestamp 1669390400
transform 1 0 62048 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_546
timestamp 1669390400
transform 1 0 62496 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_550
timestamp 1669390400
transform 1 0 62944 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_554
timestamp 1669390400
transform 1 0 63392 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_560
timestamp 1669390400
transform 1 0 64064 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_564
timestamp 1669390400
transform 1 0 64512 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_570
timestamp 1669390400
transform 1 0 65184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_573
timestamp 1669390400
transform 1 0 65520 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_577
timestamp 1669390400
transform 1 0 65968 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_581
timestamp 1669390400
transform 1 0 66416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_585
timestamp 1669390400
transform 1 0 66864 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_588
timestamp 1669390400
transform 1 0 67200 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_620
timestamp 1669390400
transform 1 0 70784 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_636
timestamp 1669390400
transform 1 0 72576 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1669390400
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_641
timestamp 1669390400
transform 1 0 73136 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_705
timestamp 1669390400
transform 1 0 80304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_709
timestamp 1669390400
transform 1 0 80752 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_712
timestamp 1669390400
transform 1 0 81088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_776
timestamp 1669390400
transform 1 0 88256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_780
timestamp 1669390400
transform 1 0 88704 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_783
timestamp 1669390400
transform 1 0 89040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_786
timestamp 1669390400
transform 1 0 89376 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_790
timestamp 1669390400
transform 1 0 89824 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_794
timestamp 1669390400
transform 1 0 90272 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_796
timestamp 1669390400
transform 1 0 90496 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_799
timestamp 1669390400
transform 1 0 90832 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_803
timestamp 1669390400
transform 1 0 91280 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_807
timestamp 1669390400
transform 1 0 91728 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_811
timestamp 1669390400
transform 1 0 92176 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_815
timestamp 1669390400
transform 1 0 92624 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_819
timestamp 1669390400
transform 1 0 93072 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_851
timestamp 1669390400
transform 1 0 96656 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_854
timestamp 1669390400
transform 1 0 96992 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_918
timestamp 1669390400
transform 1 0 104160 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_922
timestamp 1669390400
transform 1 0 104608 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_925
timestamp 1669390400
transform 1 0 104944 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_989
timestamp 1669390400
transform 1 0 112112 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_993
timestamp 1669390400
transform 1 0 112560 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_996
timestamp 1669390400
transform 1 0 112896 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_1028
timestamp 1669390400
transform 1 0 116480 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_1044
timestamp 1669390400
transform 1 0 118272 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1046
timestamp 1669390400
transform 1 0 118496 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_1049
timestamp 1669390400
transform 1 0 118832 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1051
timestamp 1669390400
transform 1 0 119056 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_1054
timestamp 1669390400
transform 1 0 119392 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1058
timestamp 1669390400
transform 1 0 119840 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_1062
timestamp 1669390400
transform 1 0 120288 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1064
timestamp 1669390400
transform 1 0 120512 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1067
timestamp 1669390400
transform 1 0 120848 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1131
timestamp 1669390400
transform 1 0 128016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1135
timestamp 1669390400
transform 1 0 128464 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_1138
timestamp 1669390400
transform 1 0 128800 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_1154
timestamp 1669390400
transform 1 0 130592 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_1158
timestamp 1669390400
transform 1 0 131040 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1160
timestamp 1669390400
transform 1 0 131264 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_1163
timestamp 1669390400
transform 1 0 131600 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_1195
timestamp 1669390400
transform 1 0 135184 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1203
timestamp 1669390400
transform 1 0 136080 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1209
timestamp 1669390400
transform 1 0 136752 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1273
timestamp 1669390400
transform 1 0 143920 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1277
timestamp 1669390400
transform 1 0 144368 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_1280
timestamp 1669390400
transform 1 0 144704 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1312
timestamp 1669390400
transform 1 0 148288 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_116
timestamp 1669390400
transform 1 0 14336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_120
timestamp 1669390400
transform 1 0 14784 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_123
timestamp 1669390400
transform 1 0 15120 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_155
timestamp 1669390400
transform 1 0 18704 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_158
timestamp 1669390400
transform 1 0 19040 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_162
timestamp 1669390400
transform 1 0 19488 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_166
timestamp 1669390400
transform 1 0 19936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_182
timestamp 1669390400
transform 1 0 21728 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_186
timestamp 1669390400
transform 1 0 22176 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_202
timestamp 1669390400
transform 1 0 23968 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_210
timestamp 1669390400
transform 1 0 24864 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_214
timestamp 1669390400
transform 1 0 25312 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_246
timestamp 1669390400
transform 1 0 28896 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_253
timestamp 1669390400
transform 1 0 29680 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_261
timestamp 1669390400
transform 1 0 30576 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_265
timestamp 1669390400
transform 1 0 31024 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_269
timestamp 1669390400
transform 1 0 31472 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_273
timestamp 1669390400
transform 1 0 31920 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_277
timestamp 1669390400
transform 1 0 32368 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_281
timestamp 1669390400
transform 1 0 32816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_287
timestamp 1669390400
transform 1 0 33488 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_303
timestamp 1669390400
transform 1 0 35280 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_311
timestamp 1669390400
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_315
timestamp 1669390400
transform 1 0 36624 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_323
timestamp 1669390400
transform 1 0 37520 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_326
timestamp 1669390400
transform 1 0 37856 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_330
timestamp 1669390400
transform 1 0 38304 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_338
timestamp 1669390400
transform 1 0 39200 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_346
timestamp 1669390400
transform 1 0 40096 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_354
timestamp 1669390400
transform 1 0 40992 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_358
timestamp 1669390400
transform 1 0 41440 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_362
timestamp 1669390400
transform 1 0 41888 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_366
timestamp 1669390400
transform 1 0 42336 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_370
timestamp 1669390400
transform 1 0 42784 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_386
timestamp 1669390400
transform 1 0 44576 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_395
timestamp 1669390400
transform 1 0 45584 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_399
timestamp 1669390400
transform 1 0 46032 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_407
timestamp 1669390400
transform 1 0 46928 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_413
timestamp 1669390400
transform 1 0 47600 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_421
timestamp 1669390400
transform 1 0 48496 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_429
timestamp 1669390400
transform 1 0 49392 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_431
timestamp 1669390400
transform 1 0 49616 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_438
timestamp 1669390400
transform 1 0 50400 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_442
timestamp 1669390400
transform 1 0 50848 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_450
timestamp 1669390400
transform 1 0 51744 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_454
timestamp 1669390400
transform 1 0 52192 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_458
timestamp 1669390400
transform 1 0 52640 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_466
timestamp 1669390400
transform 1 0 53536 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_470
timestamp 1669390400
transform 1 0 53984 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_486
timestamp 1669390400
transform 1 0 55776 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_494
timestamp 1669390400
transform 1 0 56672 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_500
timestamp 1669390400
transform 1 0 57344 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_506
timestamp 1669390400
transform 1 0 58016 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_510
timestamp 1669390400
transform 1 0 58464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_514
timestamp 1669390400
transform 1 0 58912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_517
timestamp 1669390400
transform 1 0 59248 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_519
timestamp 1669390400
transform 1 0 59472 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_522
timestamp 1669390400
transform 1 0 59808 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_526
timestamp 1669390400
transform 1 0 60256 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_528
timestamp 1669390400
transform 1 0 60480 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1669390400
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_534
timestamp 1669390400
transform 1 0 61152 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_544
timestamp 1669390400
transform 1 0 62272 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_552
timestamp 1669390400
transform 1 0 63168 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_556
timestamp 1669390400
transform 1 0 63616 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_560
timestamp 1669390400
transform 1 0 64064 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_564
timestamp 1669390400
transform 1 0 64512 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_580
timestamp 1669390400
transform 1 0 66304 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_584
timestamp 1669390400
transform 1 0 66752 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_588
timestamp 1669390400
transform 1 0 67200 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_590
timestamp 1669390400
transform 1 0 67424 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_593
timestamp 1669390400
transform 1 0 67760 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_597
timestamp 1669390400
transform 1 0 68208 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_601
timestamp 1669390400
transform 1 0 68656 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_605
timestamp 1669390400
transform 1 0 69104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_608
timestamp 1669390400
transform 1 0 69440 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_612
timestamp 1669390400
transform 1 0 69888 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_622
timestamp 1669390400
transform 1 0 71008 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_626
timestamp 1669390400
transform 1 0 71456 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_642
timestamp 1669390400
transform 1 0 73248 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_648
timestamp 1669390400
transform 1 0 73920 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_664
timestamp 1669390400
transform 1 0 75712 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_668
timestamp 1669390400
transform 1 0 76160 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_672
timestamp 1669390400
transform 1 0 76608 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_676
timestamp 1669390400
transform 1 0 77056 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_680
timestamp 1669390400
transform 1 0 77504 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_682
timestamp 1669390400
transform 1 0 77728 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_685
timestamp 1669390400
transform 1 0 78064 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_717
timestamp 1669390400
transform 1 0 81648 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_721
timestamp 1669390400
transform 1 0 82096 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_723
timestamp 1669390400
transform 1 0 82320 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_726
timestamp 1669390400
transform 1 0 82656 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_742
timestamp 1669390400
transform 1 0 84448 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_744
timestamp 1669390400
transform 1 0 84672 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_747
timestamp 1669390400
transform 1 0 85008 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_763
timestamp 1669390400
transform 1 0 86800 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_767
timestamp 1669390400
transform 1 0 87248 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_769
timestamp 1669390400
transform 1 0 87472 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_772
timestamp 1669390400
transform 1 0 87808 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_788
timestamp 1669390400
transform 1 0 89600 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_804
timestamp 1669390400
transform 1 0 91392 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_806
timestamp 1669390400
transform 1 0 91616 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_809
timestamp 1669390400
transform 1 0 91952 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_813
timestamp 1669390400
transform 1 0 92400 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_815
timestamp 1669390400
transform 1 0 92624 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_818
timestamp 1669390400
transform 1 0 92960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_821
timestamp 1669390400
transform 1 0 93296 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_825
timestamp 1669390400
transform 1 0 93744 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_829
timestamp 1669390400
transform 1 0 94192 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_835
timestamp 1669390400
transform 1 0 94864 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_839
timestamp 1669390400
transform 1 0 95312 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_855
timestamp 1669390400
transform 1 0 97104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_858
timestamp 1669390400
transform 1 0 97440 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_862
timestamp 1669390400
transform 1 0 97888 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_866
timestamp 1669390400
transform 1 0 98336 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_870
timestamp 1669390400
transform 1 0 98784 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_874
timestamp 1669390400
transform 1 0 99232 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_881
timestamp 1669390400
transform 1 0 100016 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_885
timestamp 1669390400
transform 1 0 100464 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_889
timestamp 1669390400
transform 1 0 100912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_892
timestamp 1669390400
transform 1 0 101248 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_896
timestamp 1669390400
transform 1 0 101696 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_906
timestamp 1669390400
transform 1 0 102816 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_914
timestamp 1669390400
transform 1 0 103712 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_918
timestamp 1669390400
transform 1 0 104160 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_922
timestamp 1669390400
transform 1 0 104608 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_926
timestamp 1669390400
transform 1 0 105056 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_930
timestamp 1669390400
transform 1 0 105504 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_934
timestamp 1669390400
transform 1 0 105952 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_938
timestamp 1669390400
transform 1 0 106400 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_942
timestamp 1669390400
transform 1 0 106848 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_946
timestamp 1669390400
transform 1 0 107296 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_950
timestamp 1669390400
transform 1 0 107744 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_954
timestamp 1669390400
transform 1 0 108192 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_960
timestamp 1669390400
transform 1 0 108864 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_976
timestamp 1669390400
transform 1 0 110656 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_984
timestamp 1669390400
transform 1 0 111552 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_988
timestamp 1669390400
transform 1 0 112000 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1004
timestamp 1669390400
transform 1 0 113792 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1008
timestamp 1669390400
transform 1 0 114240 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_1012
timestamp 1669390400
transform 1 0 114688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1028
timestamp 1669390400
transform 1 0 116480 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1031
timestamp 1669390400
transform 1 0 116816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1034
timestamp 1669390400
transform 1 0 117152 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1038
timestamp 1669390400
transform 1 0 117600 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1042
timestamp 1669390400
transform 1 0 118048 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1050
timestamp 1669390400
transform 1 0 118944 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1058
timestamp 1669390400
transform 1 0 119840 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1062
timestamp 1669390400
transform 1 0 120288 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1066
timestamp 1669390400
transform 1 0 120736 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1070
timestamp 1669390400
transform 1 0 121184 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1076
timestamp 1669390400
transform 1 0 121856 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1080
timestamp 1669390400
transform 1 0 122304 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1086
timestamp 1669390400
transform 1 0 122976 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1096
timestamp 1669390400
transform 1 0 124096 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1102
timestamp 1669390400
transform 1 0 124768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_1105
timestamp 1669390400
transform 1 0 125104 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_1121
timestamp 1669390400
transform 1 0 126896 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1129
timestamp 1669390400
transform 1 0 127792 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1133
timestamp 1669390400
transform 1 0 128240 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1148
timestamp 1669390400
transform 1 0 129920 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1164
timestamp 1669390400
transform 1 0 131712 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1168
timestamp 1669390400
transform 1 0 132160 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1170
timestamp 1669390400
transform 1 0 132384 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1173
timestamp 1669390400
transform 1 0 132720 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_1179
timestamp 1669390400
transform 1 0 133392 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_1195
timestamp 1669390400
transform 1 0 135184 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1203
timestamp 1669390400
transform 1 0 136080 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1207
timestamp 1669390400
transform 1 0 136528 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1210
timestamp 1669390400
transform 1 0 136864 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1228
timestamp 1669390400
transform 1 0 138880 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1232
timestamp 1669390400
transform 1 0 139328 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1236
timestamp 1669390400
transform 1 0 139776 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1240
timestamp 1669390400
transform 1 0 140224 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_1244
timestamp 1669390400
transform 1 0 140672 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1260
timestamp 1669390400
transform 1 0 142464 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_1263
timestamp 1669390400
transform 1 0 142800 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_1295
timestamp 1669390400
transform 1 0 146384 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1311
timestamp 1669390400
transform 1 0 148176 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_34
timestamp 1669390400
transform 1 0 5152 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_50
timestamp 1669390400
transform 1 0 6944 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_54
timestamp 1669390400
transform 1 0 7392 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_62
timestamp 1669390400
transform 1 0 8288 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_75
timestamp 1669390400
transform 1 0 9744 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_78
timestamp 1669390400
transform 1 0 10080 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_82
timestamp 1669390400
transform 1 0 10528 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_90
timestamp 1669390400
transform 1 0 11424 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_94
timestamp 1669390400
transform 1 0 11872 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_110
timestamp 1669390400
transform 1 0 13664 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_120
timestamp 1669390400
transform 1 0 14784 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_124
timestamp 1669390400
transform 1 0 15232 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_128
timestamp 1669390400
transform 1 0 15680 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_135
timestamp 1669390400
transform 1 0 16464 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_139
timestamp 1669390400
transform 1 0 16912 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_148
timestamp 1669390400
transform 1 0 17920 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_156
timestamp 1669390400
transform 1 0 18816 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_164
timestamp 1669390400
transform 1 0 19712 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_180
timestamp 1669390400
transform 1 0 21504 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_188
timestamp 1669390400
transform 1 0 22400 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_192
timestamp 1669390400
transform 1 0 22848 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_196
timestamp 1669390400
transform 1 0 23296 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_200
timestamp 1669390400
transform 1 0 23744 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_204
timestamp 1669390400
transform 1 0 24192 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_223
timestamp 1669390400
transform 1 0 26320 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_233
timestamp 1669390400
transform 1 0 27440 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_235
timestamp 1669390400
transform 1 0 27664 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_238
timestamp 1669390400
transform 1 0 28000 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_240
timestamp 1669390400
transform 1 0 28224 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_243
timestamp 1669390400
transform 1 0 28560 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_247
timestamp 1669390400
transform 1 0 29008 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_251
timestamp 1669390400
transform 1 0 29456 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_267
timestamp 1669390400
transform 1 0 31248 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_289
timestamp 1669390400
transform 1 0 33712 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_293
timestamp 1669390400
transform 1 0 34160 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_295
timestamp 1669390400
transform 1 0 34384 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_298
timestamp 1669390400
transform 1 0 34720 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_304
timestamp 1669390400
transform 1 0 35392 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_308
timestamp 1669390400
transform 1 0 35840 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_312
timestamp 1669390400
transform 1 0 36288 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_316
timestamp 1669390400
transform 1 0 36736 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_324
timestamp 1669390400
transform 1 0 37632 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_340
timestamp 1669390400
transform 1 0 39424 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_346
timestamp 1669390400
transform 1 0 40096 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_361
timestamp 1669390400
transform 1 0 41776 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_369
timestamp 1669390400
transform 1 0 42672 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_371
timestamp 1669390400
transform 1 0 42896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_374
timestamp 1669390400
transform 1 0 43232 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_384
timestamp 1669390400
transform 1 0 44352 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_388
timestamp 1669390400
transform 1 0 44800 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_404
timestamp 1669390400
transform 1 0 46592 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_420
timestamp 1669390400
transform 1 0 48384 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_424
timestamp 1669390400
transform 1 0 48832 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_443
timestamp 1669390400
transform 1 0 50960 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_445
timestamp 1669390400
transform 1 0 51184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_452
timestamp 1669390400
transform 1 0 51968 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_468
timestamp 1669390400
transform 1 0 53760 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_476
timestamp 1669390400
transform 1 0 54656 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_480
timestamp 1669390400
transform 1 0 55104 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_488
timestamp 1669390400
transform 1 0 56000 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_492
timestamp 1669390400
transform 1 0 56448 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_506
timestamp 1669390400
transform 1 0 58016 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_516
timestamp 1669390400
transform 1 0 59136 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_520
timestamp 1669390400
transform 1 0 59584 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_524
timestamp 1669390400
transform 1 0 60032 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_532
timestamp 1669390400
transform 1 0 60928 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_548
timestamp 1669390400
transform 1 0 62720 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_558
timestamp 1669390400
transform 1 0 63840 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_566
timestamp 1669390400
transform 1 0 64736 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_570
timestamp 1669390400
transform 1 0 65184 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_572
timestamp 1669390400
transform 1 0 65408 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_575
timestamp 1669390400
transform 1 0 65744 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_591
timestamp 1669390400
transform 1 0 67536 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_608
timestamp 1669390400
transform 1 0 69440 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_624
timestamp 1669390400
transform 1 0 71232 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_628
timestamp 1669390400
transform 1 0 71680 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_632
timestamp 1669390400
transform 1 0 72128 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1669390400
transform 1 0 72800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_641
timestamp 1669390400
transform 1 0 73136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_648
timestamp 1669390400
transform 1 0 73920 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_652
timestamp 1669390400
transform 1 0 74368 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_656
timestamp 1669390400
transform 1 0 74816 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_660
timestamp 1669390400
transform 1 0 75264 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_666
timestamp 1669390400
transform 1 0 75936 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_668
timestamp 1669390400
transform 1 0 76160 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_671
timestamp 1669390400
transform 1 0 76496 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_679
timestamp 1669390400
transform 1 0 77392 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_683
timestamp 1669390400
transform 1 0 77840 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_687
timestamp 1669390400
transform 1 0 78288 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_691
timestamp 1669390400
transform 1 0 78736 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_695
timestamp 1669390400
transform 1 0 79184 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_699
timestamp 1669390400
transform 1 0 79632 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_702
timestamp 1669390400
transform 1 0 79968 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_706
timestamp 1669390400
transform 1 0 80416 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_709
timestamp 1669390400
transform 1 0 80752 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_712
timestamp 1669390400
transform 1 0 81088 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_716
timestamp 1669390400
transform 1 0 81536 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_732
timestamp 1669390400
transform 1 0 83328 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_738
timestamp 1669390400
transform 1 0 84000 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_742
timestamp 1669390400
transform 1 0 84448 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_745
timestamp 1669390400
transform 1 0 84784 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_749
timestamp 1669390400
transform 1 0 85232 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_753
timestamp 1669390400
transform 1 0 85680 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_761
timestamp 1669390400
transform 1 0 86576 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_763
timestamp 1669390400
transform 1 0 86800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_766
timestamp 1669390400
transform 1 0 87136 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_772
timestamp 1669390400
transform 1 0 87808 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_776
timestamp 1669390400
transform 1 0 88256 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_780
timestamp 1669390400
transform 1 0 88704 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_783
timestamp 1669390400
transform 1 0 89040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_790
timestamp 1669390400
transform 1 0 89824 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_807
timestamp 1669390400
transform 1 0 91728 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_823
timestamp 1669390400
transform 1 0 93520 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_827
timestamp 1669390400
transform 1 0 93968 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_831
timestamp 1669390400
transform 1 0 94416 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_835
timestamp 1669390400
transform 1 0 94864 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_839
timestamp 1669390400
transform 1 0 95312 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_843
timestamp 1669390400
transform 1 0 95760 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_847
timestamp 1669390400
transform 1 0 96208 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_851
timestamp 1669390400
transform 1 0 96656 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_854
timestamp 1669390400
transform 1 0 96992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_869
timestamp 1669390400
transform 1 0 98672 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_873
timestamp 1669390400
transform 1 0 99120 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_877
timestamp 1669390400
transform 1 0 99568 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_892
timestamp 1669390400
transform 1 0 101248 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_896
timestamp 1669390400
transform 1 0 101696 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_900
timestamp 1669390400
transform 1 0 102144 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_906
timestamp 1669390400
transform 1 0 102816 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_922
timestamp 1669390400
transform 1 0 104608 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_925
timestamp 1669390400
transform 1 0 104944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_940
timestamp 1669390400
transform 1 0 106624 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_956
timestamp 1669390400
transform 1 0 108416 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_960
timestamp 1669390400
transform 1 0 108864 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_964
timestamp 1669390400
transform 1 0 109312 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_968
timestamp 1669390400
transform 1 0 109760 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_972
timestamp 1669390400
transform 1 0 110208 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_976
timestamp 1669390400
transform 1 0 110656 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_980
timestamp 1669390400
transform 1 0 111104 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_984
timestamp 1669390400
transform 1 0 111552 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_986
timestamp 1669390400
transform 1 0 111776 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_989
timestamp 1669390400
transform 1 0 112112 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_993
timestamp 1669390400
transform 1 0 112560 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_996
timestamp 1669390400
transform 1 0 112896 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1013
timestamp 1669390400
transform 1 0 114800 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1017
timestamp 1669390400
transform 1 0 115248 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1021
timestamp 1669390400
transform 1 0 115696 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1036
timestamp 1669390400
transform 1 0 117376 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1044
timestamp 1669390400
transform 1 0 118272 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1048
timestamp 1669390400
transform 1 0 118720 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1064
timestamp 1669390400
transform 1 0 120512 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1067
timestamp 1669390400
transform 1 0 120848 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1069
timestamp 1669390400
transform 1 0 121072 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1084
timestamp 1669390400
transform 1 0 122752 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1100
timestamp 1669390400
transform 1 0 124544 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1104
timestamp 1669390400
transform 1 0 124992 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1108
timestamp 1669390400
transform 1 0 125440 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1112
timestamp 1669390400
transform 1 0 125888 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1116
timestamp 1669390400
transform 1 0 126336 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_1120
timestamp 1669390400
transform 1 0 126784 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1138
timestamp 1669390400
transform 1 0 128800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1141
timestamp 1669390400
transform 1 0 129136 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1145
timestamp 1669390400
transform 1 0 129584 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1149
timestamp 1669390400
transform 1 0 130032 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1166
timestamp 1669390400
transform 1 0 131936 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1174
timestamp 1669390400
transform 1 0 132832 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1178
timestamp 1669390400
transform 1 0 133280 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1185
timestamp 1669390400
transform 1 0 134064 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1189
timestamp 1669390400
transform 1 0 134512 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1193
timestamp 1669390400
transform 1 0 134960 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1197
timestamp 1669390400
transform 1 0 135408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1201
timestamp 1669390400
transform 1 0 135856 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1203
timestamp 1669390400
transform 1 0 136080 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1206
timestamp 1669390400
transform 1 0 136416 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1209
timestamp 1669390400
transform 1 0 136752 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1212
timestamp 1669390400
transform 1 0 137088 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1216
timestamp 1669390400
transform 1 0 137536 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1235
timestamp 1669390400
transform 1 0 139664 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1251
timestamp 1669390400
transform 1 0 141456 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1253
timestamp 1669390400
transform 1 0 141680 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1256
timestamp 1669390400
transform 1 0 142016 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1260
timestamp 1669390400
transform 1 0 142464 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1277
timestamp 1669390400
transform 1 0 144368 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1280
timestamp 1669390400
transform 1 0 144704 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_1295
timestamp 1669390400
transform 1 0 146384 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1311
timestamp 1669390400
transform 1 0 148176 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_52
timestamp 1669390400
transform 1 0 7168 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_68
timestamp 1669390400
transform 1 0 8960 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_76
timestamp 1669390400
transform 1 0 9856 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_92
timestamp 1669390400
transform 1 0 11648 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_100
timestamp 1669390400
transform 1 0 12544 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_102
timestamp 1669390400
transform 1 0 12768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_124
timestamp 1669390400
transform 1 0 15232 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_126
timestamp 1669390400
transform 1 0 15456 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_129
timestamp 1669390400
transform 1 0 15792 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_137
timestamp 1669390400
transform 1 0 16688 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_153
timestamp 1669390400
transform 1 0 18480 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_170
timestamp 1669390400
transform 1 0 20384 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_174
timestamp 1669390400
transform 1 0 20832 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_194
timestamp 1669390400
transform 1 0 23072 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_212
timestamp 1669390400
transform 1 0 25088 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_216
timestamp 1669390400
transform 1 0 25536 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_231
timestamp 1669390400
transform 1 0 27216 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_266
timestamp 1669390400
transform 1 0 31136 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_270
timestamp 1669390400
transform 1 0 31584 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_286
timestamp 1669390400
transform 1 0 33376 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_302
timestamp 1669390400
transform 1 0 35168 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_337
timestamp 1669390400
transform 1 0 39088 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_341
timestamp 1669390400
transform 1 0 39536 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_356
timestamp 1669390400
transform 1 0 41216 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_372
timestamp 1669390400
transform 1 0 43008 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_388
timestamp 1669390400
transform 1 0 44800 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_396
timestamp 1669390400
transform 1 0 45696 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_404
timestamp 1669390400
transform 1 0 46592 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_421
timestamp 1669390400
transform 1 0 48496 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_438
timestamp 1669390400
transform 1 0 50400 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_454
timestamp 1669390400
transform 1 0 52192 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1669390400
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_465
timestamp 1669390400
transform 1 0 53424 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_468
timestamp 1669390400
transform 1 0 53760 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_484
timestamp 1669390400
transform 1 0 55552 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_488
timestamp 1669390400
transform 1 0 56000 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_491
timestamp 1669390400
transform 1 0 56336 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_499
timestamp 1669390400
transform 1 0 57232 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_515
timestamp 1669390400
transform 1 0 59024 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1669390400
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_534
timestamp 1669390400
transform 1 0 61152 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_546
timestamp 1669390400
transform 1 0 62496 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_562
timestamp 1669390400
transform 1 0 64288 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_579
timestamp 1669390400
transform 1 0 66192 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_585
timestamp 1669390400
transform 1 0 66864 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1669390400
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_605
timestamp 1669390400
transform 1 0 69104 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_607
timestamp 1669390400
transform 1 0 69328 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_610
timestamp 1669390400
transform 1 0 69664 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_628
timestamp 1669390400
transform 1 0 71680 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_644
timestamp 1669390400
transform 1 0 73472 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_660
timestamp 1669390400
transform 1 0 75264 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_670
timestamp 1669390400
transform 1 0 76384 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_676
timestamp 1669390400
transform 1 0 77056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_683
timestamp 1669390400
transform 1 0 77840 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_691
timestamp 1669390400
transform 1 0 78736 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_695
timestamp 1669390400
transform 1 0 79184 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_699
timestamp 1669390400
transform 1 0 79632 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_701
timestamp 1669390400
transform 1 0 79856 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_716
timestamp 1669390400
transform 1 0 81536 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_732
timestamp 1669390400
transform 1 0 83328 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_736
timestamp 1669390400
transform 1 0 83776 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_743
timestamp 1669390400
transform 1 0 84560 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_747
timestamp 1669390400
transform 1 0 85008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_762
timestamp 1669390400
transform 1 0 86688 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_780
timestamp 1669390400
transform 1 0 88704 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_784
timestamp 1669390400
transform 1 0 89152 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_801
timestamp 1669390400
transform 1 0 91056 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_805
timestamp 1669390400
transform 1 0 91504 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_815
timestamp 1669390400
transform 1 0 92624 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_818
timestamp 1669390400
transform 1 0 92960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_833
timestamp 1669390400
transform 1 0 94640 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_849
timestamp 1669390400
transform 1 0 96432 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_865
timestamp 1669390400
transform 1 0 98224 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_881
timestamp 1669390400
transform 1 0 100016 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_885
timestamp 1669390400
transform 1 0 100464 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_889
timestamp 1669390400
transform 1 0 100912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_904
timestamp 1669390400
transform 1 0 102592 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_920
timestamp 1669390400
transform 1 0 104384 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_922
timestamp 1669390400
transform 1 0 104608 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_931
timestamp 1669390400
transform 1 0 105616 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_948
timestamp 1669390400
transform 1 0 107520 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_956
timestamp 1669390400
transform 1 0 108416 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_960
timestamp 1669390400
transform 1 0 108864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_975
timestamp 1669390400
transform 1 0 110544 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_991
timestamp 1669390400
transform 1 0 112336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1010
timestamp 1669390400
transform 1 0 114464 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1026
timestamp 1669390400
transform 1 0 116256 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1028
timestamp 1669390400
transform 1 0 116480 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1031
timestamp 1669390400
transform 1 0 116816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1034
timestamp 1669390400
transform 1 0 117152 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1052
timestamp 1669390400
transform 1 0 119168 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1071
timestamp 1669390400
transform 1 0 121296 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1075
timestamp 1669390400
transform 1 0 121744 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1077
timestamp 1669390400
transform 1 0 121968 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1093
timestamp 1669390400
transform 1 0 123760 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1097
timestamp 1669390400
transform 1 0 124208 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1099
timestamp 1669390400
transform 1 0 124432 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1102
timestamp 1669390400
transform 1 0 124768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1117
timestamp 1669390400
transform 1 0 126448 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1133
timestamp 1669390400
transform 1 0 128240 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1137
timestamp 1669390400
transform 1 0 128688 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1140
timestamp 1669390400
transform 1 0 129024 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1144
timestamp 1669390400
transform 1 0 129472 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1161
timestamp 1669390400
transform 1 0 131376 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1169
timestamp 1669390400
transform 1 0 132272 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1173
timestamp 1669390400
transform 1 0 132720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1188
timestamp 1669390400
transform 1 0 134400 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1196
timestamp 1669390400
transform 1 0 135296 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1212
timestamp 1669390400
transform 1 0 137088 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1216
timestamp 1669390400
transform 1 0 137536 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1233
timestamp 1669390400
transform 1 0 139440 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1237
timestamp 1669390400
transform 1 0 139888 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1241
timestamp 1669390400
transform 1 0 140336 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1244
timestamp 1669390400
transform 1 0 140672 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1260
timestamp 1669390400
transform 1 0 142464 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1264
timestamp 1669390400
transform 1 0 142912 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1268
timestamp 1669390400
transform 1 0 143360 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1286
timestamp 1669390400
transform 1 0 145376 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_1290
timestamp 1669390400
transform 1 0 145824 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1306
timestamp 1669390400
transform 1 0 147616 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1310
timestamp 1669390400
transform 1 0 148064 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1312
timestamp 1669390400
transform 1 0 148288 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_34
timestamp 1669390400
transform 1 0 5152 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_38
timestamp 1669390400
transform 1 0 5600 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_54
timestamp 1669390400
transform 1 0 7392 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_76
timestamp 1669390400
transform 1 0 9856 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_78
timestamp 1669390400
transform 1 0 10080 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_93
timestamp 1669390400
transform 1 0 11760 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_109
timestamp 1669390400
transform 1 0 13552 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_125
timestamp 1669390400
transform 1 0 15344 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_159
timestamp 1669390400
transform 1 0 19152 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_176
timestamp 1669390400
transform 1 0 21056 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_180
timestamp 1669390400
transform 1 0 21504 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_196
timestamp 1669390400
transform 1 0 23296 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_218
timestamp 1669390400
transform 1 0 25760 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_236
timestamp 1669390400
transform 1 0 27776 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_254
timestamp 1669390400
transform 1 0 29792 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_273
timestamp 1669390400
transform 1 0 31920 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_303
timestamp 1669390400
transform 1 0 35280 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_305
timestamp 1669390400
transform 1 0 35504 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_308
timestamp 1669390400
transform 1 0 35840 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_316
timestamp 1669390400
transform 1 0 36736 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_334
timestamp 1669390400
transform 1 0 38752 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_351
timestamp 1669390400
transform 1 0 40656 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_374
timestamp 1669390400
transform 1 0 43232 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_378
timestamp 1669390400
transform 1 0 43680 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_396
timestamp 1669390400
transform 1 0 45696 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_414
timestamp 1669390400
transform 1 0 47712 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_418
timestamp 1669390400
transform 1 0 48160 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_446
timestamp 1669390400
transform 1 0 51296 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_456
timestamp 1669390400
transform 1 0 52416 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_460
timestamp 1669390400
transform 1 0 52864 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_478
timestamp 1669390400
transform 1 0 54880 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1669390400
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_516
timestamp 1669390400
transform 1 0 59136 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_524
timestamp 1669390400
transform 1 0 60032 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_542
timestamp 1669390400
transform 1 0 62048 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_546
timestamp 1669390400
transform 1 0 62496 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_549
timestamp 1669390400
transform 1 0 62832 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1669390400
transform 1 0 64848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_570
timestamp 1669390400
transform 1 0 65184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_586
timestamp 1669390400
transform 1 0 66976 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_606
timestamp 1669390400
transform 1 0 69216 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_612
timestamp 1669390400
transform 1 0 69888 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_620
timestamp 1669390400
transform 1 0 70784 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1669390400
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_641
timestamp 1669390400
transform 1 0 73136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_658
timestamp 1669390400
transform 1 0 75040 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_675
timestamp 1669390400
transform 1 0 76944 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_691
timestamp 1669390400
transform 1 0 78736 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_707
timestamp 1669390400
transform 1 0 80528 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_709
timestamp 1669390400
transform 1 0 80752 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_712
timestamp 1669390400
transform 1 0 81088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_719
timestamp 1669390400
transform 1 0 81872 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_723
timestamp 1669390400
transform 1 0 82320 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_725
timestamp 1669390400
transform 1 0 82544 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_742
timestamp 1669390400
transform 1 0 84448 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_758
timestamp 1669390400
transform 1 0 86240 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_774
timestamp 1669390400
transform 1 0 88032 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_778
timestamp 1669390400
transform 1 0 88480 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_780
timestamp 1669390400
transform 1 0 88704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_783
timestamp 1669390400
transform 1 0 89040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_799
timestamp 1669390400
transform 1 0 90832 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_816
timestamp 1669390400
transform 1 0 92736 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_833
timestamp 1669390400
transform 1 0 94640 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_849
timestamp 1669390400
transform 1 0 96432 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_851
timestamp 1669390400
transform 1 0 96656 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_854
timestamp 1669390400
transform 1 0 96992 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_864
timestamp 1669390400
transform 1 0 98112 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_881
timestamp 1669390400
transform 1 0 100016 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_891
timestamp 1669390400
transform 1 0 101136 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_893
timestamp 1669390400
transform 1 0 101360 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_910
timestamp 1669390400
transform 1 0 103264 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_912
timestamp 1669390400
transform 1 0 103488 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_919
timestamp 1669390400
transform 1 0 104272 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_925
timestamp 1669390400
transform 1 0 104944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_928
timestamp 1669390400
transform 1 0 105280 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_932
timestamp 1669390400
transform 1 0 105728 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_950
timestamp 1669390400
transform 1 0 107744 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_958
timestamp 1669390400
transform 1 0 108640 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_962
timestamp 1669390400
transform 1 0 109088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_982
timestamp 1669390400
transform 1 0 111328 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_990
timestamp 1669390400
transform 1 0 112224 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_996
timestamp 1669390400
transform 1 0 112896 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1014
timestamp 1669390400
transform 1 0 114912 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1022
timestamp 1669390400
transform 1 0 115808 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1026
timestamp 1669390400
transform 1 0 116256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1046
timestamp 1669390400
transform 1 0 118496 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1048
timestamp 1669390400
transform 1 0 118720 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1064
timestamp 1669390400
transform 1 0 120512 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1067
timestamp 1669390400
transform 1 0 120848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1084
timestamp 1669390400
transform 1 0 122752 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1092
timestamp 1669390400
transform 1 0 123648 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1110
timestamp 1669390400
transform 1 0 125664 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1128
timestamp 1669390400
transform 1 0 127680 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1132
timestamp 1669390400
transform 1 0 128128 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1138
timestamp 1669390400
transform 1 0 128800 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1158
timestamp 1669390400
transform 1 0 131040 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1166
timestamp 1669390400
transform 1 0 131936 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1170
timestamp 1669390400
transform 1 0 132384 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1190
timestamp 1669390400
transform 1 0 134624 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1206
timestamp 1669390400
transform 1 0 136416 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1209
timestamp 1669390400
transform 1 0 136752 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1226
timestamp 1669390400
transform 1 0 138656 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1234
timestamp 1669390400
transform 1 0 139552 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1254
timestamp 1669390400
transform 1 0 141792 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1271
timestamp 1669390400
transform 1 0 143696 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1275
timestamp 1669390400
transform 1 0 144144 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1277
timestamp 1669390400
transform 1 0 144368 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1280
timestamp 1669390400
transform 1 0 144704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1297
timestamp 1669390400
transform 1 0 146608 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_1301
timestamp 1669390400
transform 1 0 147056 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1309
timestamp 1669390400
transform 1 0 147952 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_18
timestamp 1669390400
transform 1 0 3360 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_26
timestamp 1669390400
transform 1 0 4256 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_43
timestamp 1669390400
transform 1 0 6160 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_51
timestamp 1669390400
transform 1 0 7056 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_69
timestamp 1669390400
transform 1 0 9072 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_72
timestamp 1669390400
transform 1 0 9408 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_78
timestamp 1669390400
transform 1 0 10080 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_86
timestamp 1669390400
transform 1 0 10976 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_104
timestamp 1669390400
transform 1 0 12992 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_107
timestamp 1669390400
transform 1 0 13328 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_113
timestamp 1669390400
transform 1 0 14000 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_121
timestamp 1669390400
transform 1 0 14896 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_139
timestamp 1669390400
transform 1 0 16912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_142
timestamp 1669390400
transform 1 0 17248 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_148
timestamp 1669390400
transform 1 0 17920 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_156
timestamp 1669390400
transform 1 0 18816 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_174
timestamp 1669390400
transform 1 0 20832 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_177
timestamp 1669390400
transform 1 0 21168 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_180
timestamp 1669390400
transform 1 0 21504 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_188
timestamp 1669390400
transform 1 0 22400 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_206
timestamp 1669390400
transform 1 0 24416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_212
timestamp 1669390400
transform 1 0 25088 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_230
timestamp 1669390400
transform 1 0 27104 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_236
timestamp 1669390400
transform 1 0 27776 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_244
timestamp 1669390400
transform 1 0 28672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_251
timestamp 1669390400
transform 1 0 29456 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_259
timestamp 1669390400
transform 1 0 30352 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_261
timestamp 1669390400
transform 1 0 30576 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_278
timestamp 1669390400
transform 1 0 32480 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_282
timestamp 1669390400
transform 1 0 32928 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_288
timestamp 1669390400
transform 1 0 33600 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_296
timestamp 1669390400
transform 1 0 34496 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_314
timestamp 1669390400
transform 1 0 36512 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_317
timestamp 1669390400
transform 1 0 36848 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_323
timestamp 1669390400
transform 1 0 37520 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_331
timestamp 1669390400
transform 1 0 38416 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_349
timestamp 1669390400
transform 1 0 40432 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_352
timestamp 1669390400
transform 1 0 40768 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_356
timestamp 1669390400
transform 1 0 41216 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_364
timestamp 1669390400
transform 1 0 42112 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_382
timestamp 1669390400
transform 1 0 44128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_384
timestamp 1669390400
transform 1 0 44352 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_387
timestamp 1669390400
transform 1 0 44688 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_393
timestamp 1669390400
transform 1 0 45360 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_401
timestamp 1669390400
transform 1 0 46256 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_419
timestamp 1669390400
transform 1 0 48272 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_422
timestamp 1669390400
transform 1 0 48608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_428
timestamp 1669390400
transform 1 0 49280 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_436
timestamp 1669390400
transform 1 0 50176 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_454
timestamp 1669390400
transform 1 0 52192 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_457
timestamp 1669390400
transform 1 0 52528 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_471
timestamp 1669390400
transform 1 0 54096 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_489
timestamp 1669390400
transform 1 0 56112 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_492
timestamp 1669390400
transform 1 0 56448 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_498
timestamp 1669390400
transform 1 0 57120 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_506
timestamp 1669390400
transform 1 0 58016 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_524
timestamp 1669390400
transform 1 0 60032 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_527
timestamp 1669390400
transform 1 0 60368 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_529
timestamp 1669390400
transform 1 0 60592 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_532
timestamp 1669390400
transform 1 0 60928 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_540
timestamp 1669390400
transform 1 0 61824 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_558
timestamp 1669390400
transform 1 0 63840 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_562
timestamp 1669390400
transform 1 0 64288 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_572
timestamp 1669390400
transform 1 0 65408 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_590
timestamp 1669390400
transform 1 0 67424 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_594
timestamp 1669390400
transform 1 0 67872 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_597
timestamp 1669390400
transform 1 0 68208 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_600
timestamp 1669390400
transform 1 0 68544 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_604
timestamp 1669390400
transform 1 0 68992 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_622
timestamp 1669390400
transform 1 0 71008 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_626
timestamp 1669390400
transform 1 0 71456 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_629
timestamp 1669390400
transform 1 0 71792 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_632
timestamp 1669390400
transform 1 0 72128 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_638
timestamp 1669390400
transform 1 0 72800 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_646
timestamp 1669390400
transform 1 0 73696 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_664
timestamp 1669390400
transform 1 0 75712 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_667
timestamp 1669390400
transform 1 0 76048 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_683
timestamp 1669390400
transform 1 0 77840 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_699
timestamp 1669390400
transform 1 0 79632 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_702
timestamp 1669390400
transform 1 0 79968 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_719
timestamp 1669390400
transform 1 0 81872 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_727
timestamp 1669390400
transform 1 0 82768 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_731
timestamp 1669390400
transform 1 0 83216 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_737
timestamp 1669390400
transform 1 0 83888 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_744
timestamp 1669390400
transform 1 0 84672 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_748
timestamp 1669390400
transform 1 0 85120 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_752
timestamp 1669390400
transform 1 0 85568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_769
timestamp 1669390400
transform 1 0 87472 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_772
timestamp 1669390400
transform 1 0 87808 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_774
timestamp 1669390400
transform 1 0 88032 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_781
timestamp 1669390400
transform 1 0 88816 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_785
timestamp 1669390400
transform 1 0 89264 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_787
timestamp 1669390400
transform 1 0 89488 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_804
timestamp 1669390400
transform 1 0 91392 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_807
timestamp 1669390400
transform 1 0 91728 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_814
timestamp 1669390400
transform 1 0 92512 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_818
timestamp 1669390400
transform 1 0 92960 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_838
timestamp 1669390400
transform 1 0 95200 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_842
timestamp 1669390400
transform 1 0 95648 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_862
timestamp 1669390400
transform 1 0 97888 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_870
timestamp 1669390400
transform 1 0 98784 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_874
timestamp 1669390400
transform 1 0 99232 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_877
timestamp 1669390400
transform 1 0 99568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_894
timestamp 1669390400
transform 1 0 101472 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_898
timestamp 1669390400
transform 1 0 101920 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_907
timestamp 1669390400
transform 1 0 102928 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_909
timestamp 1669390400
transform 1 0 103152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_912
timestamp 1669390400
transform 1 0 103488 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_915
timestamp 1669390400
transform 1 0 103824 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_917
timestamp 1669390400
transform 1 0 104048 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_934
timestamp 1669390400
transform 1 0 105952 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_944
timestamp 1669390400
transform 1 0 107072 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_947
timestamp 1669390400
transform 1 0 107408 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_949
timestamp 1669390400
transform 1 0 107632 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_966
timestamp 1669390400
transform 1 0 109536 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_974
timestamp 1669390400
transform 1 0 110432 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_978
timestamp 1669390400
transform 1 0 110880 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_982
timestamp 1669390400
transform 1 0 111328 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_999
timestamp 1669390400
transform 1 0 113232 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1007
timestamp 1669390400
transform 1 0 114128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1011
timestamp 1669390400
transform 1 0 114576 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1017
timestamp 1669390400
transform 1 0 115248 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1034
timestamp 1669390400
transform 1 0 117152 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1042
timestamp 1669390400
transform 1 0 118048 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1046
timestamp 1669390400
transform 1 0 118496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1052
timestamp 1669390400
transform 1 0 119168 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1069
timestamp 1669390400
transform 1 0 121072 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1077
timestamp 1669390400
transform 1 0 121968 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1081
timestamp 1669390400
transform 1 0 122416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1087
timestamp 1669390400
transform 1 0 123088 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1104
timestamp 1669390400
transform 1 0 124992 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1112
timestamp 1669390400
transform 1 0 125888 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1116
timestamp 1669390400
transform 1 0 126336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1122
timestamp 1669390400
transform 1 0 127008 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1142
timestamp 1669390400
transform 1 0 129248 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1150
timestamp 1669390400
transform 1 0 130144 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1154
timestamp 1669390400
transform 1 0 130592 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1157
timestamp 1669390400
transform 1 0 130928 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1174
timestamp 1669390400
transform 1 0 132832 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1182
timestamp 1669390400
transform 1 0 133728 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1186
timestamp 1669390400
transform 1 0 134176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1192
timestamp 1669390400
transform 1 0 134848 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1209
timestamp 1669390400
transform 1 0 136752 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1217
timestamp 1669390400
transform 1 0 137648 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1221
timestamp 1669390400
transform 1 0 138096 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1227
timestamp 1669390400
transform 1 0 138768 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1244
timestamp 1669390400
transform 1 0 140672 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1248
timestamp 1669390400
transform 1 0 141120 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1252
timestamp 1669390400
transform 1 0 141568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1259
timestamp 1669390400
transform 1 0 142352 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1262
timestamp 1669390400
transform 1 0 142688 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1279
timestamp 1669390400
transform 1 0 144592 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1287
timestamp 1669390400
transform 1 0 145488 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1291
timestamp 1669390400
transform 1 0 145936 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1297
timestamp 1669390400
transform 1 0 146608 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1312
timestamp 1669390400
transform 1 0 148288 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 148624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 148624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 148624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 148624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 148624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 148624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 148624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 148624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 148624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 148624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 148624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 148624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 148624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 148624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 148624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 148624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 148624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 148624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 148624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 148624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 148624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 148624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 148624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 148624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 148624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 148624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 148624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 148624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 148624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 148624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 148624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 148624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 148624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 148624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 148624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 148624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 148624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 148624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 148624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 148624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 148624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 148624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 148624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1669390400
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1669390400
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1669390400
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1669390400
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1669390400
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1669390400
transform 1 0 79744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1669390400
transform 1 0 83664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1669390400
transform 1 0 87584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1669390400
transform 1 0 91504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1669390400
transform 1 0 95424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1669390400
transform 1 0 99344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1669390400
transform 1 0 103264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1669390400
transform 1 0 107184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1669390400
transform 1 0 111104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1669390400
transform 1 0 115024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1669390400
transform 1 0 118944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1669390400
transform 1 0 122864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1669390400
transform 1 0 126784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1669390400
transform 1 0 130704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1669390400
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1669390400
transform 1 0 138544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1669390400
transform 1 0 142464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1669390400
transform 1 0 146384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1669390400
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1669390400
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1669390400
transform 1 0 80864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1669390400
transform 1 0 88816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1669390400
transform 1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1669390400
transform 1 0 104720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1669390400
transform 1 0 112672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1669390400
transform 1 0 120624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1669390400
transform 1 0 128576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1669390400
transform 1 0 136528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1669390400
transform 1 0 144480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 84784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 92736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 100688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 108640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 116592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 124544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 132496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 140448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 80864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 88816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 96768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 104720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 112672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 120624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 128576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 136528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 144480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 84784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 92736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 100688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 108640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 116592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 124544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 132496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 140448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 80864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 88816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 96768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 104720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 112672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 120624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 128576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 136528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 144480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 84784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 92736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 100688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 108640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 116592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 124544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 132496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 140448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 88816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 104720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 112672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 120624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 128576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 136528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 144480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 84784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 92736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 100688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 108640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 116592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 124544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 132496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 140448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 80864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 88816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 96768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 104720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 112672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 120624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 128576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 136528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 144480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 84784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 92736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 100688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 108640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 116592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 124544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 132496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 140448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 80864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 88816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 96768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 104720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 112672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 120624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 128576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 136528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 144480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 84784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 92736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 100688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 108640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 116592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 124544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 132496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 140448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 80864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 88816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 96768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 104720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 112672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 120624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 128576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 136528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 144480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 84784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 92736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 100688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 108640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 116592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 124544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 132496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 140448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 80864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 88816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 96768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 104720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 112672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 120624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 128576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 136528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 144480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 84784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 92736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 100688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 108640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 116592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 124544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 132496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 140448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 80864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 88816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 96768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 104720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 112672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 120624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 128576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 136528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 144480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 84784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 92736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 100688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 108640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 116592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 124544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 132496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 140448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 80864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 88816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 96768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 104720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 112672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 120624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 128576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 136528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 144480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 84784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 92736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 100688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 108640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 116592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 124544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 132496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 140448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 80864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 88816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 96768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 104720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 112672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 120624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 128576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 136528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 144480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 84784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 92736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 100688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 108640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 116592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 124544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 132496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 140448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 80864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 88816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 96768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 104720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 112672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 120624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 128576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 136528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 144480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 84784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 92736 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 100688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 108640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 116592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 124544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 132496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 140448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 80864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 88816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 96768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 104720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 112672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 120624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 128576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 136528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 144480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 84784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 92736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 100688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 108640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 116592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 124544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 132496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 140448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 80864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 88816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 96768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 104720 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 112672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 120624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 128576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 136528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 144480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 84784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 92736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 100688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 108640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 116592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 124544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 132496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1669390400
transform 1 0 140448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1669390400
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1669390400
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1669390400
transform 1 0 80864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1669390400
transform 1 0 88816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1669390400
transform 1 0 96768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1669390400
transform 1 0 104720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1669390400
transform 1 0 112672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1669390400
transform 1 0 120624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1669390400
transform 1 0 128576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1669390400
transform 1 0 136528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1669390400
transform 1 0 144480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1669390400
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1669390400
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1669390400
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1669390400
transform 1 0 84784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1669390400
transform 1 0 92736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1669390400
transform 1 0 100688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1669390400
transform 1 0 108640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1669390400
transform 1 0 116592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1669390400
transform 1 0 124544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1669390400
transform 1 0 132496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1669390400
transform 1 0 140448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1669390400
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1669390400
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1669390400
transform 1 0 80864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1669390400
transform 1 0 88816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1669390400
transform 1 0 96768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1669390400
transform 1 0 104720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1669390400
transform 1 0 112672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1669390400
transform 1 0 120624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1669390400
transform 1 0 128576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1669390400
transform 1 0 136528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1669390400
transform 1 0 144480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1669390400
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1669390400
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1669390400
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1669390400
transform 1 0 84784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1669390400
transform 1 0 92736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1669390400
transform 1 0 100688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1669390400
transform 1 0 108640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1669390400
transform 1 0 116592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1669390400
transform 1 0 124544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1669390400
transform 1 0 132496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1669390400
transform 1 0 140448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1669390400
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1669390400
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1669390400
transform 1 0 80864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1669390400
transform 1 0 88816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1669390400
transform 1 0 96768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1669390400
transform 1 0 104720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1669390400
transform 1 0 112672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1669390400
transform 1 0 120624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1669390400
transform 1 0 128576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1669390400
transform 1 0 136528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1669390400
transform 1 0 144480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1669390400
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1669390400
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1669390400
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1669390400
transform 1 0 84784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1669390400
transform 1 0 92736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1669390400
transform 1 0 100688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1669390400
transform 1 0 108640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1669390400
transform 1 0 116592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1669390400
transform 1 0 124544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1669390400
transform 1 0 132496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1669390400
transform 1 0 140448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1669390400
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1669390400
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1669390400
transform 1 0 80864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1669390400
transform 1 0 88816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1669390400
transform 1 0 96768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1669390400
transform 1 0 104720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1669390400
transform 1 0 112672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1669390400
transform 1 0 120624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1669390400
transform 1 0 128576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1669390400
transform 1 0 136528 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1669390400
transform 1 0 144480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1669390400
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1669390400
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1669390400
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1669390400
transform 1 0 84784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1669390400
transform 1 0 92736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1669390400
transform 1 0 100688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1669390400
transform 1 0 108640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1669390400
transform 1 0 116592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1669390400
transform 1 0 124544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1669390400
transform 1 0 132496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1669390400
transform 1 0 140448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1669390400
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1669390400
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1669390400
transform 1 0 80864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1669390400
transform 1 0 88816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1669390400
transform 1 0 96768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1669390400
transform 1 0 104720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1669390400
transform 1 0 112672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1669390400
transform 1 0 120624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1669390400
transform 1 0 128576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1669390400
transform 1 0 136528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1669390400
transform 1 0 144480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1669390400
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1669390400
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1669390400
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1669390400
transform 1 0 84784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1669390400
transform 1 0 92736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1669390400
transform 1 0 100688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1669390400
transform 1 0 108640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1669390400
transform 1 0 116592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1669390400
transform 1 0 124544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1669390400
transform 1 0 132496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1669390400
transform 1 0 140448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1669390400
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1669390400
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1669390400
transform 1 0 80864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1669390400
transform 1 0 88816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1669390400
transform 1 0 96768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1669390400
transform 1 0 104720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1669390400
transform 1 0 112672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1669390400
transform 1 0 120624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1669390400
transform 1 0 128576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1669390400
transform 1 0 136528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1669390400
transform 1 0 144480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1669390400
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1669390400
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1669390400
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1669390400
transform 1 0 84784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1669390400
transform 1 0 92736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1669390400
transform 1 0 100688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1669390400
transform 1 0 108640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1669390400
transform 1 0 116592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1669390400
transform 1 0 124544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1669390400
transform 1 0 132496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1669390400
transform 1 0 140448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1669390400
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1669390400
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1669390400
transform 1 0 80864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1669390400
transform 1 0 88816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1669390400
transform 1 0 96768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1669390400
transform 1 0 104720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1669390400
transform 1 0 112672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1669390400
transform 1 0 120624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1669390400
transform 1 0 128576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1669390400
transform 1 0 136528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1669390400
transform 1 0 144480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1669390400
transform 1 0 9184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1669390400
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1669390400
transform 1 0 17024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1669390400
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1669390400
transform 1 0 24864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1669390400
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1669390400
transform 1 0 32704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1669390400
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1669390400
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1669390400
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1669390400
transform 1 0 48384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1669390400
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1669390400
transform 1 0 56224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1669390400
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1669390400
transform 1 0 64064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1669390400
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1669390400
transform 1 0 71904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1669390400
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1669390400
transform 1 0 79744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1669390400
transform 1 0 83664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1669390400
transform 1 0 87584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1669390400
transform 1 0 91504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1669390400
transform 1 0 95424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1669390400
transform 1 0 99344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1669390400
transform 1 0 103264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1669390400
transform 1 0 107184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1669390400
transform 1 0 111104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1669390400
transform 1 0 115024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1669390400
transform 1 0 118944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1669390400
transform 1 0 122864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1669390400
transform 1 0 126784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1669390400
transform 1 0 130704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1669390400
transform 1 0 134624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1669390400
transform 1 0 138544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1669390400
transform 1 0 142464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1669390400
transform 1 0 146384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _168_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 62496 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _169_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 92736 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _170_
timestamp 1669390400
transform -1 0 50848 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _171_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 141232 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _172_
timestamp 1669390400
transform 1 0 128912 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _173_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 127792 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _174_
timestamp 1669390400
transform -1 0 91728 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _175_
timestamp 1669390400
transform 1 0 126784 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _176_
timestamp 1669390400
transform 1 0 127232 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _177_
timestamp 1669390400
transform -1 0 62496 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _178_
timestamp 1669390400
transform 1 0 106176 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _179_
timestamp 1669390400
transform -1 0 144368 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _180_
timestamp 1669390400
transform -1 0 144032 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _181_
timestamp 1669390400
transform -1 0 142912 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _182_
timestamp 1669390400
transform 1 0 142016 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _183_
timestamp 1669390400
transform 1 0 141568 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _184_
timestamp 1669390400
transform -1 0 142016 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _185_
timestamp 1669390400
transform -1 0 114464 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _186_
timestamp 1669390400
transform 1 0 110880 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _187_
timestamp 1669390400
transform 1 0 113792 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _188_
timestamp 1669390400
transform 1 0 111888 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _189_
timestamp 1669390400
transform -1 0 120512 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _190_
timestamp 1669390400
transform 1 0 118608 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _191_
timestamp 1669390400
transform -1 0 119504 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _192_
timestamp 1669390400
transform 1 0 104720 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _193_
timestamp 1669390400
transform -1 0 114800 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _194_
timestamp 1669390400
transform 1 0 113680 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _195_
timestamp 1669390400
transform 1 0 110880 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _196_
timestamp 1669390400
transform -1 0 107520 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _197_
timestamp 1669390400
transform 1 0 108304 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _198_
timestamp 1669390400
transform 1 0 107856 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _199_
timestamp 1669390400
transform -1 0 139440 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _200_
timestamp 1669390400
transform 1 0 142128 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _201_
timestamp 1669390400
transform 1 0 137760 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _202_
timestamp 1669390400
transform -1 0 136416 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _203_
timestamp 1669390400
transform -1 0 139664 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _204_
timestamp 1669390400
transform -1 0 140000 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _205_
timestamp 1669390400
transform -1 0 137536 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _206_
timestamp 1669390400
transform 1 0 63168 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _207_
timestamp 1669390400
transform 1 0 102032 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _208_
timestamp 1669390400
transform -1 0 131376 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _209_
timestamp 1669390400
transform 1 0 143920 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _210_
timestamp 1669390400
transform -1 0 144256 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _211_
timestamp 1669390400
transform -1 0 131936 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _212_
timestamp 1669390400
transform 1 0 144816 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _213_
timestamp 1669390400
transform -1 0 144256 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _214_
timestamp 1669390400
transform -1 0 123760 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _215_
timestamp 1669390400
transform 1 0 51072 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _216_
timestamp 1669390400
transform 1 0 90272 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _217_
timestamp 1669390400
transform -1 0 122640 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _218_
timestamp 1669390400
transform -1 0 122304 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _219_
timestamp 1669390400
transform -1 0 121296 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _220_
timestamp 1669390400
transform 1 0 118832 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _221_
timestamp 1669390400
transform -1 0 118608 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _222_
timestamp 1669390400
transform 1 0 100240 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _223_
timestamp 1669390400
transform -1 0 100016 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _224_
timestamp 1669390400
transform 1 0 98896 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _225_
timestamp 1669390400
transform 1 0 99120 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _226_
timestamp 1669390400
transform -1 0 90832 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _227_
timestamp 1669390400
transform 1 0 90608 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _228_
timestamp 1669390400
transform 1 0 91392 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _229_
timestamp 1669390400
transform 1 0 89376 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _230_
timestamp 1669390400
transform -1 0 88704 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _231_
timestamp 1669390400
transform 1 0 86800 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _232_
timestamp 1669390400
transform -1 0 86688 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _233_
timestamp 1669390400
transform -1 0 94640 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _234_
timestamp 1669390400
transform -1 0 90384 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _235_
timestamp 1669390400
transform 1 0 89152 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _236_
timestamp 1669390400
transform 1 0 75488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _237_
timestamp 1669390400
transform -1 0 76944 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _238_
timestamp 1669390400
transform -1 0 76048 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _239_
timestamp 1669390400
transform -1 0 77840 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _240_
timestamp 1669390400
transform -1 0 77840 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _241_
timestamp 1669390400
transform -1 0 77616 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _242_
timestamp 1669390400
transform 1 0 78064 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _243_
timestamp 1669390400
transform -1 0 68768 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _244_
timestamp 1669390400
transform 1 0 65408 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _245_
timestamp 1669390400
transform 1 0 67088 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _246_
timestamp 1669390400
transform -1 0 66864 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _247_
timestamp 1669390400
transform -1 0 69440 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _248_
timestamp 1669390400
transform -1 0 68768 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _249_
timestamp 1669390400
transform -1 0 68320 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _250_
timestamp 1669390400
transform -1 0 65408 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _251_
timestamp 1669390400
transform -1 0 66976 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _252_
timestamp 1669390400
transform 1 0 65296 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _253_
timestamp 1669390400
transform -1 0 64064 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _254_
timestamp 1669390400
transform -1 0 66192 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _255_
timestamp 1669390400
transform 1 0 65296 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _256_
timestamp 1669390400
transform -1 0 63056 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _257_
timestamp 1669390400
transform -1 0 50400 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _258_
timestamp 1669390400
transform -1 0 50512 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _259_
timestamp 1669390400
transform -1 0 50848 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _260_
timestamp 1669390400
transform 1 0 51968 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _261_
timestamp 1669390400
transform -1 0 48496 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _262_
timestamp 1669390400
transform 1 0 47264 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _263_
timestamp 1669390400
transform -1 0 47152 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _264_
timestamp 1669390400
transform -1 0 62272 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _265_
timestamp 1669390400
transform -1 0 39088 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _266_
timestamp 1669390400
transform 1 0 37296 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _267_
timestamp 1669390400
transform -1 0 36960 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _268_
timestamp 1669390400
transform -1 0 40656 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _269_
timestamp 1669390400
transform -1 0 39760 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _270_
timestamp 1669390400
transform 1 0 39200 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _271_
timestamp 1669390400
transform -1 0 31920 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _272_
timestamp 1669390400
transform 1 0 20160 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _273_
timestamp 1669390400
transform 1 0 29456 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _274_
timestamp 1669390400
transform -1 0 28896 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _275_
timestamp 1669390400
transform 1 0 29456 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _276_
timestamp 1669390400
transform 1 0 26544 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _277_
timestamp 1669390400
transform -1 0 26320 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _278_
timestamp 1669390400
transform -1 0 21056 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _279_
timestamp 1669390400
transform 1 0 18144 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _280_
timestamp 1669390400
transform 1 0 15568 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _281_
timestamp 1669390400
transform -1 0 20384 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _282_
timestamp 1669390400
transform 1 0 17920 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _283_
timestamp 1669390400
transform 1 0 16464 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _284_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 14224 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _285_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 10640 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _286_
timestamp 1669390400
transform -1 0 8624 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _287_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6048 0 1 3136
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _288_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 52416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _289_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 72240 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _290_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 52416 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _291_
timestamp 1669390400
transform -1 0 50400 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _292_
timestamp 1669390400
transform 1 0 56560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _293_
timestamp 1669390400
transform -1 0 60032 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _294_
timestamp 1669390400
transform -1 0 29792 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _295_
timestamp 1669390400
transform -1 0 21952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _296_
timestamp 1669390400
transform -1 0 20832 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _297_
timestamp 1669390400
transform -1 0 28448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _298_
timestamp 1669390400
transform -1 0 32256 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _299_
timestamp 1669390400
transform 1 0 56336 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _300_
timestamp 1669390400
transform -1 0 58352 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _301_
timestamp 1669390400
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _302_
timestamp 1669390400
transform -1 0 41888 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _303_
timestamp 1669390400
transform -1 0 48832 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _304_
timestamp 1669390400
transform -1 0 53760 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _305_
timestamp 1669390400
transform -1 0 71680 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _306_
timestamp 1669390400
transform -1 0 64848 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _307_
timestamp 1669390400
transform -1 0 69664 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _308_
timestamp 1669390400
transform -1 0 71456 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _309_
timestamp 1669390400
transform -1 0 68768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _310_
timestamp 1669390400
transform -1 0 91280 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _311_
timestamp 1669390400
transform -1 0 79520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _312_
timestamp 1669390400
transform -1 0 80528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _313_
timestamp 1669390400
transform 1 0 91504 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _314_
timestamp 1669390400
transform -1 0 89712 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _315_
timestamp 1669390400
transform 1 0 94080 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _316_
timestamp 1669390400
transform 1 0 97664 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _317_
timestamp 1669390400
transform 1 0 101808 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _318_
timestamp 1669390400
transform 1 0 119728 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _319_
timestamp 1669390400
transform 1 0 116032 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _320_
timestamp 1669390400
transform -1 0 135408 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _321_
timestamp 1669390400
transform -1 0 135408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _322_
timestamp 1669390400
transform -1 0 133952 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _323_
timestamp 1669390400
transform -1 0 131824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _324_
timestamp 1669390400
transform 1 0 132048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _325_
timestamp 1669390400
transform -1 0 112896 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _326_
timestamp 1669390400
transform -1 0 112000 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _327_
timestamp 1669390400
transform -1 0 116480 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _328_
timestamp 1669390400
transform 1 0 119280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _329_
timestamp 1669390400
transform -1 0 115808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _330_
timestamp 1669390400
transform -1 0 133616 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _331_
timestamp 1669390400
transform -1 0 134288 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _332_
timestamp 1669390400
transform -1 0 133280 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _333_
timestamp 1669390400
transform -1 0 132272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _334_
timestamp 1669390400
transform -1 0 132272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _335_
timestamp 1669390400
transform -1 0 16688 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _336_
timestamp 1669390400
transform -1 0 11984 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _337_
timestamp 1669390400
transform -1 0 12320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _338_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17136 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _339_
timestamp 1669390400
transform 1 0 16128 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _340_
timestamp 1669390400
transform 1 0 24976 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _341_
timestamp 1669390400
transform 1 0 27776 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _342_
timestamp 1669390400
transform -1 0 41216 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _343_
timestamp 1669390400
transform 1 0 35392 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _344_
timestamp 1669390400
transform 1 0 45136 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _345_
timestamp 1669390400
transform -1 0 52864 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _346_
timestamp 1669390400
transform 1 0 61040 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _347_
timestamp 1669390400
transform 1 0 62160 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _348_
timestamp 1669390400
transform 1 0 66976 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _349_
timestamp 1669390400
transform 1 0 63616 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _350_
timestamp 1669390400
transform -1 0 80080 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _351_
timestamp 1669390400
transform -1 0 76720 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _352_
timestamp 1669390400
transform 1 0 89152 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _353_
timestamp 1669390400
transform 1 0 85232 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _354_
timestamp 1669390400
transform 1 0 94976 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _355_
timestamp 1669390400
transform 1 0 99456 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _356_
timestamp 1669390400
transform 1 0 116928 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _357_
timestamp 1669390400
transform -1 0 120288 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _358_
timestamp 1669390400
transform -1 0 131936 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _359_
timestamp 1669390400
transform -1 0 132720 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _360_
timestamp 1669390400
transform 1 0 124656 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _361_
timestamp 1669390400
transform -1 0 136640 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _362_
timestamp 1669390400
transform 1 0 107968 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _363_
timestamp 1669390400
transform 1 0 113008 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _364_
timestamp 1669390400
transform 1 0 117600 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _365_
timestamp 1669390400
transform 1 0 111776 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _366_
timestamp 1669390400
transform 1 0 128912 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _367_
timestamp 1669390400
transform 1 0 128912 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _368_
timestamp 1669390400
transform 1 0 127792 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _369_
timestamp 1669390400
transform 1 0 127792 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _370_
timestamp 1669390400
transform 1 0 12880 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _371_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7280 0 1 4704
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _372_
timestamp 1669390400
transform 1 0 7168 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _375_
timestamp 1669390400
transform -1 0 8288 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _376_
timestamp 1669390400
transform -1 0 11424 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _377_
timestamp 1669390400
transform -1 0 16464 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _378_
timestamp 1669390400
transform -1 0 22400 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _379_
timestamp 1669390400
transform -1 0 38416 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _380_
timestamp 1669390400
transform -1 0 42112 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _381_
timestamp 1669390400
transform -1 0 48944 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _382_
timestamp 1669390400
transform -1 0 49392 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _383_
timestamp 1669390400
transform -1 0 46592 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _384_
timestamp 1669390400
transform 1 0 29680 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _385_
timestamp 1669390400
transform 1 0 40320 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _386_
timestamp 1669390400
transform 1 0 49504 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _387_
timestamp 1669390400
transform 1 0 60256 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _388_
timestamp 1669390400
transform 1 0 57344 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _389_
timestamp 1669390400
transform 1 0 77168 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _390_
timestamp 1669390400
transform 1 0 84000 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _391_
timestamp 1669390400
transform 1 0 81200 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _392_
timestamp 1669390400
transform 1 0 76720 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _393_
timestamp 1669390400
transform 1 0 6384 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _394_
timestamp 1669390400
transform -1 0 10976 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _395_
timestamp 1669390400
transform -1 0 14896 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _396_
timestamp 1669390400
transform -1 0 19712 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _397_
timestamp 1669390400
transform -1 0 33040 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _398_
timestamp 1669390400
transform -1 0 37632 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _399_
timestamp 1669390400
transform -1 0 34496 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _400_
timestamp 1669390400
transform -1 0 40096 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _401_
timestamp 1669390400
transform -1 0 46928 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _402_
timestamp 1669390400
transform -1 0 48496 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _403_
timestamp 1669390400
transform -1 0 51744 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _404_
timestamp 1669390400
transform -1 0 46256 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _405_
timestamp 1669390400
transform -1 0 51968 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _406_
timestamp 1669390400
transform -1 0 54096 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _407_
timestamp 1669390400
transform -1 0 73696 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _408_
timestamp 1669390400
transform -1 0 60032 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _409_
timestamp 1669390400
transform -1 0 58016 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _410_
timestamp 1669390400
transform -1 0 54656 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _411_
timestamp 1669390400
transform -1 0 57232 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _412_
timestamp 1669390400
transform -1 0 70784 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _413_
timestamp 1669390400
transform -1 0 61824 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _414_
timestamp 1669390400
transform -1 0 84560 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _415_
timestamp 1669390400
transform -1 0 89824 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _416_
timestamp 1669390400
transform -1 0 100016 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _417_
timestamp 1669390400
transform -1 0 110432 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _418_
timestamp 1669390400
transform -1 0 118272 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _419_
timestamp 1669390400
transform -1 0 119840 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _420_
timestamp 1669390400
transform -1 0 125888 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _421_
timestamp 1669390400
transform -1 0 133728 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _422_
timestamp 1669390400
transform -1 0 124096 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _423_
timestamp 1669390400
transform -1 0 78736 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _424_
timestamp 1669390400
transform 1 0 73248 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _425_
timestamp 1669390400
transform 1 0 16016 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _426_
timestamp 1669390400
transform 1 0 21728 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _427_
timestamp 1669390400
transform 1 0 36064 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _428_
timestamp 1669390400
transform 1 0 42000 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _429_
timestamp 1669390400
transform 1 0 58464 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _430_
timestamp 1669390400
transform 1 0 64064 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _431_
timestamp 1669390400
transform 1 0 88144 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _432_
timestamp 1669390400
transform 1 0 98112 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _433_
timestamp 1669390400
transform 1 0 91840 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _434_
timestamp 1669390400
transform 1 0 91952 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _435_
timestamp 1669390400
transform 1 0 82096 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _436_
timestamp 1669390400
transform 1 0 97440 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _437_
timestamp 1669390400
transform 1 0 103600 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _438_
timestamp 1669390400
transform 1 0 107744 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _439_
timestamp 1669390400
transform 1 0 111552 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _440_
timestamp 1669390400
transform 1 0 115136 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _441_
timestamp 1669390400
transform 1 0 117376 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _442_
timestamp 1669390400
transform -1 0 121968 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _443_
timestamp 1669390400
transform -1 0 123648 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _444_
timestamp 1669390400
transform 1 0 107968 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _445_
timestamp 1669390400
transform 1 0 113456 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _446_
timestamp 1669390400
transform 1 0 118272 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _447_
timestamp 1669390400
transform -1 0 130144 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _448_
timestamp 1669390400
transform -1 0 131936 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _449_
timestamp 1669390400
transform 1 0 131600 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _450_
timestamp 1669390400
transform 1 0 132160 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _451_
timestamp 1669390400
transform 1 0 133392 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _452_
timestamp 1669390400
transform 1 0 134624 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _453_
timestamp 1669390400
transform 1 0 136976 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _454_
timestamp 1669390400
transform 1 0 138880 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _455_
timestamp 1669390400
transform 1 0 141680 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _456_
timestamp 1669390400
transform -1 0 145488 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _457_
timestamp 1669390400
transform -1 0 9856 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _458_
timestamp 1669390400
transform -1 0 14784 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _459_
timestamp 1669390400
transform -1 0 18816 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _460_
timestamp 1669390400
transform 1 0 18144 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _461_
timestamp 1669390400
transform 1 0 38528 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _462_
timestamp 1669390400
transform 1 0 25648 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _463_
timestamp 1669390400
transform 1 0 28000 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _464_
timestamp 1669390400
transform 1 0 40320 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_io_wbs_clk dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 71120 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_io_wbs_clk
timestamp 1669390400
transform -1 0 70896 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_io_wbs_clk
timestamp 1669390400
transform -1 0 66864 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_io_wbs_clk
timestamp 1669390400
transform 1 0 75152 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_io_wbs_clk
timestamp 1669390400
transform 1 0 77168 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7280 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform 1 0 36960 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform 1 0 38640 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input4
timestamp 1669390400
transform 1 0 41440 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input5
timestamp 1669390400
transform 1 0 42336 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input6
timestamp 1669390400
transform 1 0 43904 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input7
timestamp 1669390400
transform 1 0 45920 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input8
timestamp 1669390400
transform 1 0 46480 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input9
timestamp 1669390400
transform 1 0 49504 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input10
timestamp 1669390400
transform 1 0 50400 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input11
timestamp 1669390400
transform 1 0 53088 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input12
timestamp 1669390400
transform 1 0 11200 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input13
timestamp 1669390400
transform 1 0 54320 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input14
timestamp 1669390400
transform 1 0 57344 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input15
timestamp 1669390400
transform 1 0 58240 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input16
timestamp 1669390400
transform 1 0 60256 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input17
timestamp 1669390400
transform 1 0 62048 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input18
timestamp 1669390400
transform 1 0 63056 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input19
timestamp 1669390400
transform 1 0 65632 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input20
timestamp 1669390400
transform 1 0 67424 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input21
timestamp 1669390400
transform 1 0 69216 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input22
timestamp 1669390400
transform 1 0 71008 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input23
timestamp 1669390400
transform 1 0 15120 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input24
timestamp 1669390400
transform 1 0 73248 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input25
timestamp 1669390400
transform 1 0 73920 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input26
timestamp 1669390400
transform 1 0 19040 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input27
timestamp 1669390400
transform 1 0 22624 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input28
timestamp 1669390400
transform 1 0 25312 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input29
timestamp 1669390400
transform 1 0 28000 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input30
timestamp 1669390400
transform 1 0 30688 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input31
timestamp 1669390400
transform 1 0 33488 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input32
timestamp 1669390400
transform 1 0 34720 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input33
timestamp 1669390400
transform -1 0 81872 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input34
timestamp 1669390400
transform -1 0 109536 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input35
timestamp 1669390400
transform -1 0 111328 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input36
timestamp 1669390400
transform -1 0 113232 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input37
timestamp 1669390400
transform -1 0 114912 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input38
timestamp 1669390400
transform -1 0 117152 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input39
timestamp 1669390400
transform -1 0 118496 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input40
timestamp 1669390400
transform -1 0 121072 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input41
timestamp 1669390400
transform -1 0 122752 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input42
timestamp 1669390400
transform -1 0 124992 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input43
timestamp 1669390400
transform -1 0 125664 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input44
timestamp 1669390400
transform -1 0 84448 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input45
timestamp 1669390400
transform 1 0 125888 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input46
timestamp 1669390400
transform 1 0 127456 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input47
timestamp 1669390400
transform 1 0 129248 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input48
timestamp 1669390400
transform 1 0 131040 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input49
timestamp 1669390400
transform -1 0 134624 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input50
timestamp 1669390400
transform -1 0 136752 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input51
timestamp 1669390400
transform -1 0 138656 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input52
timestamp 1669390400
transform -1 0 140672 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input53
timestamp 1669390400
transform 1 0 140000 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input54
timestamp 1669390400
transform 1 0 142800 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input55
timestamp 1669390400
transform -1 0 87472 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input56
timestamp 1669390400
transform -1 0 145376 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input57
timestamp 1669390400
transform -1 0 146608 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input58
timestamp 1669390400
transform -1 0 91392 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input59
timestamp 1669390400
transform -1 0 95200 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input60
timestamp 1669390400
transform -1 0 97888 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input61
timestamp 1669390400
transform -1 0 101472 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input62
timestamp 1669390400
transform -1 0 103264 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input63
timestamp 1669390400
transform -1 0 105952 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input64
timestamp 1669390400
transform -1 0 107744 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input65
timestamp 1669390400
transform 1 0 58240 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input66 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 61152 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input67
timestamp 1669390400
transform -1 0 24752 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input68
timestamp 1669390400
transform 1 0 28672 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input69
timestamp 1669390400
transform 1 0 34048 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input70
timestamp 1669390400
transform 1 0 38080 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input71
timestamp 1669390400
transform 1 0 42112 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input72
timestamp 1669390400
transform 1 0 46144 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input73
timestamp 1669390400
transform 1 0 50176 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input74
timestamp 1669390400
transform 1 0 54208 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input75
timestamp 1669390400
transform 1 0 7168 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input76
timestamp 1669390400
transform -1 0 16912 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input77
timestamp 1669390400
transform 1 0 61264 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input78
timestamp 1669390400
transform 1 0 64960 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input79
timestamp 1669390400
transform 1 0 68992 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input80
timestamp 1669390400
transform 1 0 72912 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input81
timestamp 1669390400
transform 1 0 77056 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input82
timestamp 1669390400
transform -1 0 83552 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input83
timestamp 1669390400
transform -1 0 87472 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input84
timestamp 1669390400
transform -1 0 91392 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input85
timestamp 1669390400
transform -1 0 95312 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input86
timestamp 1669390400
transform 1 0 97216 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input87
timestamp 1669390400
transform -1 0 21728 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input88
timestamp 1669390400
transform 1 0 101248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input89
timestamp 1669390400
transform 1 0 105280 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input90
timestamp 1669390400
transform 1 0 109200 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input91
timestamp 1669390400
transform -1 0 114912 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input92
timestamp 1669390400
transform -1 0 118832 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input93
timestamp 1669390400
transform -1 0 122752 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input94
timestamp 1669390400
transform -1 0 126672 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input95
timestamp 1669390400
transform -1 0 130592 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input96
timestamp 1669390400
transform 1 0 132720 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input97
timestamp 1669390400
transform 1 0 137536 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input98
timestamp 1669390400
transform 1 0 25984 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input99
timestamp 1669390400
transform 1 0 141568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input100
timestamp 1669390400
transform -1 0 146272 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input101
timestamp 1669390400
transform -1 0 33040 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input102
timestamp 1669390400
transform -1 0 36512 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input103
timestamp 1669390400
transform 1 0 41440 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input104
timestamp 1669390400
transform 1 0 45360 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input105
timestamp 1669390400
transform 1 0 49392 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input106
timestamp 1669390400
transform 1 0 52864 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input107
timestamp 1669390400
transform 1 0 57344 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input108
timestamp 1669390400
transform 1 0 7280 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input109
timestamp 1669390400
transform 1 0 17360 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input110
timestamp 1669390400
transform 1 0 21952 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input111
timestamp 1669390400
transform 1 0 26880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input112
timestamp 1669390400
transform -1 0 32592 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input113
timestamp 1669390400
transform -1 0 11648 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input114
timestamp 1669390400
transform -1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output115 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 7392 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output116
timestamp 1669390400
transform -1 0 11648 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output117
timestamp 1669390400
transform -1 0 15232 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output118
timestamp 1669390400
transform -1 0 18480 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output119
timestamp 1669390400
transform -1 0 23072 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output120
timestamp 1669390400
transform -1 0 25088 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output121
timestamp 1669390400
transform -1 0 27216 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output122
timestamp 1669390400
transform -1 0 29008 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output123
timestamp 1669390400
transform -1 0 33040 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output124
timestamp 1669390400
transform 1 0 78064 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output125
timestamp 1669390400
transform 1 0 81760 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output126
timestamp 1669390400
transform 1 0 85120 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output127
timestamp 1669390400
transform 1 0 88032 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output128
timestamp 1669390400
transform -1 0 94640 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output129
timestamp 1669390400
transform 1 0 94864 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output130
timestamp 1669390400
transform 1 0 97104 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output131
timestamp 1669390400
transform 1 0 99680 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output132
timestamp 1669390400
transform 1 0 102816 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output133
timestamp 1669390400
transform 1 0 7392 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output134
timestamp 1669390400
transform -1 0 36960 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output135
timestamp 1669390400
transform -1 0 39424 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output136
timestamp 1669390400
transform -1 0 41216 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output137
timestamp 1669390400
transform -1 0 43008 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output138
timestamp 1669390400
transform -1 0 44800 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output139
timestamp 1669390400
transform -1 0 46592 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output140
timestamp 1669390400
transform -1 0 48384 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output141
timestamp 1669390400
transform -1 0 50960 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output142
timestamp 1669390400
transform -1 0 52192 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output143
timestamp 1669390400
transform -1 0 53760 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output144
timestamp 1669390400
transform 1 0 10192 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output145
timestamp 1669390400
transform -1 0 55552 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output146
timestamp 1669390400
transform -1 0 56896 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output147
timestamp 1669390400
transform -1 0 59024 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output148
timestamp 1669390400
transform -1 0 60816 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output149
timestamp 1669390400
transform -1 0 62720 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output150
timestamp 1669390400
transform -1 0 64288 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output151
timestamp 1669390400
transform -1 0 66304 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output152
timestamp 1669390400
transform -1 0 67536 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output153
timestamp 1669390400
transform -1 0 71232 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output154
timestamp 1669390400
transform -1 0 71680 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output155
timestamp 1669390400
transform 1 0 13776 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output156
timestamp 1669390400
transform -1 0 73472 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output157
timestamp 1669390400
transform 1 0 73696 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output158
timestamp 1669390400
transform -1 0 19152 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output159
timestamp 1669390400
transform -1 0 23296 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output160
timestamp 1669390400
transform -1 0 25088 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output161
timestamp 1669390400
transform -1 0 27776 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output162
timestamp 1669390400
transform -1 0 31248 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output163
timestamp 1669390400
transform -1 0 33376 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output164
timestamp 1669390400
transform -1 0 35168 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output165
timestamp 1669390400
transform 1 0 78960 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output166
timestamp 1669390400
transform 1 0 106848 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output167
timestamp 1669390400
transform 1 0 108976 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output168
timestamp 1669390400
transform 1 0 110768 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output169
timestamp 1669390400
transform 1 0 112224 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output170
timestamp 1669390400
transform 1 0 114688 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output171
timestamp 1669390400
transform 1 0 115808 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output172
timestamp 1669390400
transform 1 0 117600 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output173
timestamp 1669390400
transform -1 0 120512 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output174
timestamp 1669390400
transform -1 0 122752 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output175
timestamp 1669390400
transform 1 0 122976 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output176
timestamp 1669390400
transform 1 0 81760 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output177
timestamp 1669390400
transform -1 0 126448 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output178
timestamp 1669390400
transform 1 0 126672 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output179
timestamp 1669390400
transform -1 0 129920 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output180
timestamp 1669390400
transform -1 0 131712 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output181
timestamp 1669390400
transform 1 0 132832 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output182
timestamp 1669390400
transform 1 0 134848 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output183
timestamp 1669390400
transform 1 0 135520 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output184
timestamp 1669390400
transform 1 0 137312 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output185
timestamp 1669390400
transform 1 0 139888 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output186
timestamp 1669390400
transform 1 0 140896 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output187
timestamp 1669390400
transform -1 0 88032 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output188
timestamp 1669390400
transform 1 0 146720 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output189
timestamp 1669390400
transform 1 0 144816 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output190
timestamp 1669390400
transform 1 0 89824 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output191
timestamp 1669390400
transform 1 0 94864 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output192
timestamp 1669390400
transform 1 0 96656 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output193
timestamp 1669390400
transform 1 0 98448 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output194
timestamp 1669390400
transform 1 0 101024 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output195
timestamp 1669390400
transform 1 0 103040 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output196
timestamp 1669390400
transform 1 0 105056 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output197
timestamp 1669390400
transform -1 0 6048 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output198
timestamp 1669390400
transform -1 0 15456 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output199
timestamp 1669390400
transform -1 0 60816 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output200
timestamp 1669390400
transform -1 0 64848 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output201
timestamp 1669390400
transform -1 0 70784 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output202
timestamp 1669390400
transform -1 0 72800 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output203
timestamp 1669390400
transform -1 0 74928 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output204
timestamp 1669390400
transform -1 0 81312 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output205
timestamp 1669390400
transform -1 0 85344 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output206
timestamp 1669390400
transform -1 0 88704 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output207
timestamp 1669390400
transform -1 0 94752 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output208
timestamp 1669390400
transform -1 0 96656 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output209
timestamp 1669390400
transform -1 0 19712 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output210
timestamp 1669390400
transform -1 0 101472 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output211
timestamp 1669390400
transform -1 0 105504 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output212
timestamp 1669390400
transform -1 0 110544 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output213
timestamp 1669390400
transform -1 0 113568 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output214
timestamp 1669390400
transform -1 0 118608 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output215
timestamp 1669390400
transform 1 0 120960 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output216
timestamp 1669390400
transform 1 0 124880 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output217
timestamp 1669390400
transform 1 0 126896 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output218
timestamp 1669390400
transform -1 0 134512 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output219
timestamp 1669390400
transform -1 0 137760 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output220
timestamp 1669390400
transform -1 0 27104 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output221
timestamp 1669390400
transform 1 0 140224 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output222
timestamp 1669390400
transform 1 0 146720 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output223
timestamp 1669390400
transform -1 0 31584 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output224
timestamp 1669390400
transform -1 0 36960 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output225
timestamp 1669390400
transform 1 0 39424 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output226
timestamp 1669390400
transform -1 0 44912 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output227
timestamp 1669390400
transform -1 0 48944 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output228
timestamp 1669390400
transform -1 0 53088 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output229
timestamp 1669390400
transform -1 0 56896 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output230
timestamp 1669390400
transform -1 0 7168 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output231
timestamp 1669390400
transform 1 0 77168 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output232
timestamp 1669390400
transform -1 0 9184 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output233
timestamp 1669390400
transform -1 0 13552 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output234
timestamp 1669390400
transform -1 0 17136 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output235
timestamp 1669390400
transform 1 0 19936 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output236
timestamp 1669390400
transform 1 0 79968 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output237
timestamp 1669390400
transform -1 0 86240 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output238
timestamp 1669390400
transform 1 0 87136 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output239
timestamp 1669390400
transform 1 0 91952 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_memory_240 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 5152 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_memory_241
timestamp 1669390400
transform -1 0 75936 0 -1 34496
box -86 -86 534 870
<< labels >>
flabel metal2 s 6384 39200 6496 40000 0 FreeSans 448 90 0 0 addr_mem0[0]
port 0 nsew signal tristate
flabel metal2 s 9968 39200 10080 40000 0 FreeSans 448 90 0 0 addr_mem0[1]
port 1 nsew signal tristate
flabel metal2 s 13552 39200 13664 40000 0 FreeSans 448 90 0 0 addr_mem0[2]
port 2 nsew signal tristate
flabel metal2 s 17136 39200 17248 40000 0 FreeSans 448 90 0 0 addr_mem0[3]
port 3 nsew signal tristate
flabel metal2 s 20720 39200 20832 40000 0 FreeSans 448 90 0 0 addr_mem0[4]
port 4 nsew signal tristate
flabel metal2 s 23408 39200 23520 40000 0 FreeSans 448 90 0 0 addr_mem0[5]
port 5 nsew signal tristate
flabel metal2 s 26096 39200 26208 40000 0 FreeSans 448 90 0 0 addr_mem0[6]
port 6 nsew signal tristate
flabel metal2 s 28784 39200 28896 40000 0 FreeSans 448 90 0 0 addr_mem0[7]
port 7 nsew signal tristate
flabel metal2 s 31472 39200 31584 40000 0 FreeSans 448 90 0 0 addr_mem0[8]
port 8 nsew signal tristate
flabel metal2 s 77168 39200 77280 40000 0 FreeSans 448 90 0 0 addr_mem1[0]
port 9 nsew signal tristate
flabel metal2 s 80752 39200 80864 40000 0 FreeSans 448 90 0 0 addr_mem1[1]
port 10 nsew signal tristate
flabel metal2 s 84336 39200 84448 40000 0 FreeSans 448 90 0 0 addr_mem1[2]
port 11 nsew signal tristate
flabel metal2 s 87920 39200 88032 40000 0 FreeSans 448 90 0 0 addr_mem1[3]
port 12 nsew signal tristate
flabel metal2 s 91504 39200 91616 40000 0 FreeSans 448 90 0 0 addr_mem1[4]
port 13 nsew signal tristate
flabel metal2 s 94192 39200 94304 40000 0 FreeSans 448 90 0 0 addr_mem1[5]
port 14 nsew signal tristate
flabel metal2 s 96880 39200 96992 40000 0 FreeSans 448 90 0 0 addr_mem1[6]
port 15 nsew signal tristate
flabel metal2 s 99568 39200 99680 40000 0 FreeSans 448 90 0 0 addr_mem1[7]
port 16 nsew signal tristate
flabel metal2 s 102256 39200 102368 40000 0 FreeSans 448 90 0 0 addr_mem1[8]
port 17 nsew signal tristate
flabel metal2 s 4592 39200 4704 40000 0 FreeSans 448 90 0 0 csb_mem0
port 18 nsew signal tristate
flabel metal2 s 75376 39200 75488 40000 0 FreeSans 448 90 0 0 csb_mem1
port 19 nsew signal tristate
flabel metal2 s 7280 39200 7392 40000 0 FreeSans 448 90 0 0 din_mem0[0]
port 20 nsew signal tristate
flabel metal2 s 35952 39200 36064 40000 0 FreeSans 448 90 0 0 din_mem0[10]
port 21 nsew signal tristate
flabel metal2 s 37744 39200 37856 40000 0 FreeSans 448 90 0 0 din_mem0[11]
port 22 nsew signal tristate
flabel metal2 s 39536 39200 39648 40000 0 FreeSans 448 90 0 0 din_mem0[12]
port 23 nsew signal tristate
flabel metal2 s 41328 39200 41440 40000 0 FreeSans 448 90 0 0 din_mem0[13]
port 24 nsew signal tristate
flabel metal2 s 43120 39200 43232 40000 0 FreeSans 448 90 0 0 din_mem0[14]
port 25 nsew signal tristate
flabel metal2 s 44912 39200 45024 40000 0 FreeSans 448 90 0 0 din_mem0[15]
port 26 nsew signal tristate
flabel metal2 s 46704 39200 46816 40000 0 FreeSans 448 90 0 0 din_mem0[16]
port 27 nsew signal tristate
flabel metal2 s 48496 39200 48608 40000 0 FreeSans 448 90 0 0 din_mem0[17]
port 28 nsew signal tristate
flabel metal2 s 50288 39200 50400 40000 0 FreeSans 448 90 0 0 din_mem0[18]
port 29 nsew signal tristate
flabel metal2 s 52080 39200 52192 40000 0 FreeSans 448 90 0 0 din_mem0[19]
port 30 nsew signal tristate
flabel metal2 s 10864 39200 10976 40000 0 FreeSans 448 90 0 0 din_mem0[1]
port 31 nsew signal tristate
flabel metal2 s 53872 39200 53984 40000 0 FreeSans 448 90 0 0 din_mem0[20]
port 32 nsew signal tristate
flabel metal2 s 55664 39200 55776 40000 0 FreeSans 448 90 0 0 din_mem0[21]
port 33 nsew signal tristate
flabel metal2 s 57456 39200 57568 40000 0 FreeSans 448 90 0 0 din_mem0[22]
port 34 nsew signal tristate
flabel metal2 s 59248 39200 59360 40000 0 FreeSans 448 90 0 0 din_mem0[23]
port 35 nsew signal tristate
flabel metal2 s 61040 39200 61152 40000 0 FreeSans 448 90 0 0 din_mem0[24]
port 36 nsew signal tristate
flabel metal2 s 62832 39200 62944 40000 0 FreeSans 448 90 0 0 din_mem0[25]
port 37 nsew signal tristate
flabel metal2 s 64624 39200 64736 40000 0 FreeSans 448 90 0 0 din_mem0[26]
port 38 nsew signal tristate
flabel metal2 s 66416 39200 66528 40000 0 FreeSans 448 90 0 0 din_mem0[27]
port 39 nsew signal tristate
flabel metal2 s 68208 39200 68320 40000 0 FreeSans 448 90 0 0 din_mem0[28]
port 40 nsew signal tristate
flabel metal2 s 70000 39200 70112 40000 0 FreeSans 448 90 0 0 din_mem0[29]
port 41 nsew signal tristate
flabel metal2 s 14448 39200 14560 40000 0 FreeSans 448 90 0 0 din_mem0[2]
port 42 nsew signal tristate
flabel metal2 s 71792 39200 71904 40000 0 FreeSans 448 90 0 0 din_mem0[30]
port 43 nsew signal tristate
flabel metal2 s 73584 39200 73696 40000 0 FreeSans 448 90 0 0 din_mem0[31]
port 44 nsew signal tristate
flabel metal2 s 18032 39200 18144 40000 0 FreeSans 448 90 0 0 din_mem0[3]
port 45 nsew signal tristate
flabel metal2 s 21616 39200 21728 40000 0 FreeSans 448 90 0 0 din_mem0[4]
port 46 nsew signal tristate
flabel metal2 s 24304 39200 24416 40000 0 FreeSans 448 90 0 0 din_mem0[5]
port 47 nsew signal tristate
flabel metal2 s 26992 39200 27104 40000 0 FreeSans 448 90 0 0 din_mem0[6]
port 48 nsew signal tristate
flabel metal2 s 29680 39200 29792 40000 0 FreeSans 448 90 0 0 din_mem0[7]
port 49 nsew signal tristate
flabel metal2 s 32368 39200 32480 40000 0 FreeSans 448 90 0 0 din_mem0[8]
port 50 nsew signal tristate
flabel metal2 s 34160 39200 34272 40000 0 FreeSans 448 90 0 0 din_mem0[9]
port 51 nsew signal tristate
flabel metal2 s 78064 39200 78176 40000 0 FreeSans 448 90 0 0 din_mem1[0]
port 52 nsew signal tristate
flabel metal2 s 106736 39200 106848 40000 0 FreeSans 448 90 0 0 din_mem1[10]
port 53 nsew signal tristate
flabel metal2 s 108528 39200 108640 40000 0 FreeSans 448 90 0 0 din_mem1[11]
port 54 nsew signal tristate
flabel metal2 s 110320 39200 110432 40000 0 FreeSans 448 90 0 0 din_mem1[12]
port 55 nsew signal tristate
flabel metal2 s 112112 39200 112224 40000 0 FreeSans 448 90 0 0 din_mem1[13]
port 56 nsew signal tristate
flabel metal2 s 113904 39200 114016 40000 0 FreeSans 448 90 0 0 din_mem1[14]
port 57 nsew signal tristate
flabel metal2 s 115696 39200 115808 40000 0 FreeSans 448 90 0 0 din_mem1[15]
port 58 nsew signal tristate
flabel metal2 s 117488 39200 117600 40000 0 FreeSans 448 90 0 0 din_mem1[16]
port 59 nsew signal tristate
flabel metal2 s 119280 39200 119392 40000 0 FreeSans 448 90 0 0 din_mem1[17]
port 60 nsew signal tristate
flabel metal2 s 121072 39200 121184 40000 0 FreeSans 448 90 0 0 din_mem1[18]
port 61 nsew signal tristate
flabel metal2 s 122864 39200 122976 40000 0 FreeSans 448 90 0 0 din_mem1[19]
port 62 nsew signal tristate
flabel metal2 s 81648 39200 81760 40000 0 FreeSans 448 90 0 0 din_mem1[1]
port 63 nsew signal tristate
flabel metal2 s 124656 39200 124768 40000 0 FreeSans 448 90 0 0 din_mem1[20]
port 64 nsew signal tristate
flabel metal2 s 126448 39200 126560 40000 0 FreeSans 448 90 0 0 din_mem1[21]
port 65 nsew signal tristate
flabel metal2 s 128240 39200 128352 40000 0 FreeSans 448 90 0 0 din_mem1[22]
port 66 nsew signal tristate
flabel metal2 s 130032 39200 130144 40000 0 FreeSans 448 90 0 0 din_mem1[23]
port 67 nsew signal tristate
flabel metal2 s 131824 39200 131936 40000 0 FreeSans 448 90 0 0 din_mem1[24]
port 68 nsew signal tristate
flabel metal2 s 133616 39200 133728 40000 0 FreeSans 448 90 0 0 din_mem1[25]
port 69 nsew signal tristate
flabel metal2 s 135408 39200 135520 40000 0 FreeSans 448 90 0 0 din_mem1[26]
port 70 nsew signal tristate
flabel metal2 s 137200 39200 137312 40000 0 FreeSans 448 90 0 0 din_mem1[27]
port 71 nsew signal tristate
flabel metal2 s 138992 39200 139104 40000 0 FreeSans 448 90 0 0 din_mem1[28]
port 72 nsew signal tristate
flabel metal2 s 140784 39200 140896 40000 0 FreeSans 448 90 0 0 din_mem1[29]
port 73 nsew signal tristate
flabel metal2 s 85232 39200 85344 40000 0 FreeSans 448 90 0 0 din_mem1[2]
port 74 nsew signal tristate
flabel metal2 s 142576 39200 142688 40000 0 FreeSans 448 90 0 0 din_mem1[30]
port 75 nsew signal tristate
flabel metal2 s 144368 39200 144480 40000 0 FreeSans 448 90 0 0 din_mem1[31]
port 76 nsew signal tristate
flabel metal2 s 88816 39200 88928 40000 0 FreeSans 448 90 0 0 din_mem1[3]
port 77 nsew signal tristate
flabel metal2 s 92400 39200 92512 40000 0 FreeSans 448 90 0 0 din_mem1[4]
port 78 nsew signal tristate
flabel metal2 s 95088 39200 95200 40000 0 FreeSans 448 90 0 0 din_mem1[5]
port 79 nsew signal tristate
flabel metal2 s 97776 39200 97888 40000 0 FreeSans 448 90 0 0 din_mem1[6]
port 80 nsew signal tristate
flabel metal2 s 100464 39200 100576 40000 0 FreeSans 448 90 0 0 din_mem1[7]
port 81 nsew signal tristate
flabel metal2 s 103152 39200 103264 40000 0 FreeSans 448 90 0 0 din_mem1[8]
port 82 nsew signal tristate
flabel metal2 s 104944 39200 105056 40000 0 FreeSans 448 90 0 0 din_mem1[9]
port 83 nsew signal tristate
flabel metal2 s 8176 39200 8288 40000 0 FreeSans 448 90 0 0 dout_mem0[0]
port 84 nsew signal input
flabel metal2 s 36848 39200 36960 40000 0 FreeSans 448 90 0 0 dout_mem0[10]
port 85 nsew signal input
flabel metal2 s 38640 39200 38752 40000 0 FreeSans 448 90 0 0 dout_mem0[11]
port 86 nsew signal input
flabel metal2 s 40432 39200 40544 40000 0 FreeSans 448 90 0 0 dout_mem0[12]
port 87 nsew signal input
flabel metal2 s 42224 39200 42336 40000 0 FreeSans 448 90 0 0 dout_mem0[13]
port 88 nsew signal input
flabel metal2 s 44016 39200 44128 40000 0 FreeSans 448 90 0 0 dout_mem0[14]
port 89 nsew signal input
flabel metal2 s 45808 39200 45920 40000 0 FreeSans 448 90 0 0 dout_mem0[15]
port 90 nsew signal input
flabel metal2 s 47600 39200 47712 40000 0 FreeSans 448 90 0 0 dout_mem0[16]
port 91 nsew signal input
flabel metal2 s 49392 39200 49504 40000 0 FreeSans 448 90 0 0 dout_mem0[17]
port 92 nsew signal input
flabel metal2 s 51184 39200 51296 40000 0 FreeSans 448 90 0 0 dout_mem0[18]
port 93 nsew signal input
flabel metal2 s 52976 39200 53088 40000 0 FreeSans 448 90 0 0 dout_mem0[19]
port 94 nsew signal input
flabel metal2 s 11760 39200 11872 40000 0 FreeSans 448 90 0 0 dout_mem0[1]
port 95 nsew signal input
flabel metal2 s 54768 39200 54880 40000 0 FreeSans 448 90 0 0 dout_mem0[20]
port 96 nsew signal input
flabel metal2 s 56560 39200 56672 40000 0 FreeSans 448 90 0 0 dout_mem0[21]
port 97 nsew signal input
flabel metal2 s 58352 39200 58464 40000 0 FreeSans 448 90 0 0 dout_mem0[22]
port 98 nsew signal input
flabel metal2 s 60144 39200 60256 40000 0 FreeSans 448 90 0 0 dout_mem0[23]
port 99 nsew signal input
flabel metal2 s 61936 39200 62048 40000 0 FreeSans 448 90 0 0 dout_mem0[24]
port 100 nsew signal input
flabel metal2 s 63728 39200 63840 40000 0 FreeSans 448 90 0 0 dout_mem0[25]
port 101 nsew signal input
flabel metal2 s 65520 39200 65632 40000 0 FreeSans 448 90 0 0 dout_mem0[26]
port 102 nsew signal input
flabel metal2 s 67312 39200 67424 40000 0 FreeSans 448 90 0 0 dout_mem0[27]
port 103 nsew signal input
flabel metal2 s 69104 39200 69216 40000 0 FreeSans 448 90 0 0 dout_mem0[28]
port 104 nsew signal input
flabel metal2 s 70896 39200 71008 40000 0 FreeSans 448 90 0 0 dout_mem0[29]
port 105 nsew signal input
flabel metal2 s 15344 39200 15456 40000 0 FreeSans 448 90 0 0 dout_mem0[2]
port 106 nsew signal input
flabel metal2 s 72688 39200 72800 40000 0 FreeSans 448 90 0 0 dout_mem0[30]
port 107 nsew signal input
flabel metal2 s 74480 39200 74592 40000 0 FreeSans 448 90 0 0 dout_mem0[31]
port 108 nsew signal input
flabel metal2 s 18928 39200 19040 40000 0 FreeSans 448 90 0 0 dout_mem0[3]
port 109 nsew signal input
flabel metal2 s 22512 39200 22624 40000 0 FreeSans 448 90 0 0 dout_mem0[4]
port 110 nsew signal input
flabel metal2 s 25200 39200 25312 40000 0 FreeSans 448 90 0 0 dout_mem0[5]
port 111 nsew signal input
flabel metal2 s 27888 39200 28000 40000 0 FreeSans 448 90 0 0 dout_mem0[6]
port 112 nsew signal input
flabel metal2 s 30576 39200 30688 40000 0 FreeSans 448 90 0 0 dout_mem0[7]
port 113 nsew signal input
flabel metal2 s 33264 39200 33376 40000 0 FreeSans 448 90 0 0 dout_mem0[8]
port 114 nsew signal input
flabel metal2 s 35056 39200 35168 40000 0 FreeSans 448 90 0 0 dout_mem0[9]
port 115 nsew signal input
flabel metal2 s 78960 39200 79072 40000 0 FreeSans 448 90 0 0 dout_mem1[0]
port 116 nsew signal input
flabel metal2 s 107632 39200 107744 40000 0 FreeSans 448 90 0 0 dout_mem1[10]
port 117 nsew signal input
flabel metal2 s 109424 39200 109536 40000 0 FreeSans 448 90 0 0 dout_mem1[11]
port 118 nsew signal input
flabel metal2 s 111216 39200 111328 40000 0 FreeSans 448 90 0 0 dout_mem1[12]
port 119 nsew signal input
flabel metal2 s 113008 39200 113120 40000 0 FreeSans 448 90 0 0 dout_mem1[13]
port 120 nsew signal input
flabel metal2 s 114800 39200 114912 40000 0 FreeSans 448 90 0 0 dout_mem1[14]
port 121 nsew signal input
flabel metal2 s 116592 39200 116704 40000 0 FreeSans 448 90 0 0 dout_mem1[15]
port 122 nsew signal input
flabel metal2 s 118384 39200 118496 40000 0 FreeSans 448 90 0 0 dout_mem1[16]
port 123 nsew signal input
flabel metal2 s 120176 39200 120288 40000 0 FreeSans 448 90 0 0 dout_mem1[17]
port 124 nsew signal input
flabel metal2 s 121968 39200 122080 40000 0 FreeSans 448 90 0 0 dout_mem1[18]
port 125 nsew signal input
flabel metal2 s 123760 39200 123872 40000 0 FreeSans 448 90 0 0 dout_mem1[19]
port 126 nsew signal input
flabel metal2 s 82544 39200 82656 40000 0 FreeSans 448 90 0 0 dout_mem1[1]
port 127 nsew signal input
flabel metal2 s 125552 39200 125664 40000 0 FreeSans 448 90 0 0 dout_mem1[20]
port 128 nsew signal input
flabel metal2 s 127344 39200 127456 40000 0 FreeSans 448 90 0 0 dout_mem1[21]
port 129 nsew signal input
flabel metal2 s 129136 39200 129248 40000 0 FreeSans 448 90 0 0 dout_mem1[22]
port 130 nsew signal input
flabel metal2 s 130928 39200 131040 40000 0 FreeSans 448 90 0 0 dout_mem1[23]
port 131 nsew signal input
flabel metal2 s 132720 39200 132832 40000 0 FreeSans 448 90 0 0 dout_mem1[24]
port 132 nsew signal input
flabel metal2 s 134512 39200 134624 40000 0 FreeSans 448 90 0 0 dout_mem1[25]
port 133 nsew signal input
flabel metal2 s 136304 39200 136416 40000 0 FreeSans 448 90 0 0 dout_mem1[26]
port 134 nsew signal input
flabel metal2 s 138096 39200 138208 40000 0 FreeSans 448 90 0 0 dout_mem1[27]
port 135 nsew signal input
flabel metal2 s 139888 39200 140000 40000 0 FreeSans 448 90 0 0 dout_mem1[28]
port 136 nsew signal input
flabel metal2 s 141680 39200 141792 40000 0 FreeSans 448 90 0 0 dout_mem1[29]
port 137 nsew signal input
flabel metal2 s 86128 39200 86240 40000 0 FreeSans 448 90 0 0 dout_mem1[2]
port 138 nsew signal input
flabel metal2 s 143472 39200 143584 40000 0 FreeSans 448 90 0 0 dout_mem1[30]
port 139 nsew signal input
flabel metal2 s 145264 39200 145376 40000 0 FreeSans 448 90 0 0 dout_mem1[31]
port 140 nsew signal input
flabel metal2 s 89712 39200 89824 40000 0 FreeSans 448 90 0 0 dout_mem1[3]
port 141 nsew signal input
flabel metal2 s 93296 39200 93408 40000 0 FreeSans 448 90 0 0 dout_mem1[4]
port 142 nsew signal input
flabel metal2 s 95984 39200 96096 40000 0 FreeSans 448 90 0 0 dout_mem1[5]
port 143 nsew signal input
flabel metal2 s 98672 39200 98784 40000 0 FreeSans 448 90 0 0 dout_mem1[6]
port 144 nsew signal input
flabel metal2 s 101360 39200 101472 40000 0 FreeSans 448 90 0 0 dout_mem1[7]
port 145 nsew signal input
flabel metal2 s 104048 39200 104160 40000 0 FreeSans 448 90 0 0 dout_mem1[8]
port 146 nsew signal input
flabel metal2 s 105840 39200 105952 40000 0 FreeSans 448 90 0 0 dout_mem1[9]
port 147 nsew signal input
flabel metal2 s 4368 0 4480 800 0 FreeSans 448 90 0 0 io_wbs_ack
port 148 nsew signal tristate
flabel metal2 s 12432 0 12544 800 0 FreeSans 448 90 0 0 io_wbs_adr[0]
port 149 nsew signal input
flabel metal2 s 58128 0 58240 800 0 FreeSans 448 90 0 0 io_wbs_adr[10]
port 150 nsew signal input
flabel metal2 s 62160 0 62272 800 0 FreeSans 448 90 0 0 io_wbs_adr[11]
port 151 nsew signal input
flabel metal2 s 66192 0 66304 800 0 FreeSans 448 90 0 0 io_wbs_adr[12]
port 152 nsew signal input
flabel metal2 s 70224 0 70336 800 0 FreeSans 448 90 0 0 io_wbs_adr[13]
port 153 nsew signal input
flabel metal2 s 74256 0 74368 800 0 FreeSans 448 90 0 0 io_wbs_adr[14]
port 154 nsew signal input
flabel metal2 s 78288 0 78400 800 0 FreeSans 448 90 0 0 io_wbs_adr[15]
port 155 nsew signal input
flabel metal2 s 82320 0 82432 800 0 FreeSans 448 90 0 0 io_wbs_adr[16]
port 156 nsew signal input
flabel metal2 s 86352 0 86464 800 0 FreeSans 448 90 0 0 io_wbs_adr[17]
port 157 nsew signal input
flabel metal2 s 90384 0 90496 800 0 FreeSans 448 90 0 0 io_wbs_adr[18]
port 158 nsew signal input
flabel metal2 s 94416 0 94528 800 0 FreeSans 448 90 0 0 io_wbs_adr[19]
port 159 nsew signal input
flabel metal2 s 17808 0 17920 800 0 FreeSans 448 90 0 0 io_wbs_adr[1]
port 160 nsew signal input
flabel metal2 s 98448 0 98560 800 0 FreeSans 448 90 0 0 io_wbs_adr[20]
port 161 nsew signal input
flabel metal2 s 102480 0 102592 800 0 FreeSans 448 90 0 0 io_wbs_adr[21]
port 162 nsew signal input
flabel metal2 s 106512 0 106624 800 0 FreeSans 448 90 0 0 io_wbs_adr[22]
port 163 nsew signal input
flabel metal2 s 110544 0 110656 800 0 FreeSans 448 90 0 0 io_wbs_adr[23]
port 164 nsew signal input
flabel metal2 s 114576 0 114688 800 0 FreeSans 448 90 0 0 io_wbs_adr[24]
port 165 nsew signal input
flabel metal2 s 118608 0 118720 800 0 FreeSans 448 90 0 0 io_wbs_adr[25]
port 166 nsew signal input
flabel metal2 s 122640 0 122752 800 0 FreeSans 448 90 0 0 io_wbs_adr[26]
port 167 nsew signal input
flabel metal2 s 126672 0 126784 800 0 FreeSans 448 90 0 0 io_wbs_adr[27]
port 168 nsew signal input
flabel metal2 s 130704 0 130816 800 0 FreeSans 448 90 0 0 io_wbs_adr[28]
port 169 nsew signal input
flabel metal2 s 134736 0 134848 800 0 FreeSans 448 90 0 0 io_wbs_adr[29]
port 170 nsew signal input
flabel metal2 s 23184 0 23296 800 0 FreeSans 448 90 0 0 io_wbs_adr[2]
port 171 nsew signal input
flabel metal2 s 138768 0 138880 800 0 FreeSans 448 90 0 0 io_wbs_adr[30]
port 172 nsew signal input
flabel metal2 s 142800 0 142912 800 0 FreeSans 448 90 0 0 io_wbs_adr[31]
port 173 nsew signal input
flabel metal2 s 28560 0 28672 800 0 FreeSans 448 90 0 0 io_wbs_adr[3]
port 174 nsew signal input
flabel metal2 s 33936 0 34048 800 0 FreeSans 448 90 0 0 io_wbs_adr[4]
port 175 nsew signal input
flabel metal2 s 37968 0 38080 800 0 FreeSans 448 90 0 0 io_wbs_adr[5]
port 176 nsew signal input
flabel metal2 s 42000 0 42112 800 0 FreeSans 448 90 0 0 io_wbs_adr[6]
port 177 nsew signal input
flabel metal2 s 46032 0 46144 800 0 FreeSans 448 90 0 0 io_wbs_adr[7]
port 178 nsew signal input
flabel metal2 s 50064 0 50176 800 0 FreeSans 448 90 0 0 io_wbs_adr[8]
port 179 nsew signal input
flabel metal2 s 54096 0 54208 800 0 FreeSans 448 90 0 0 io_wbs_adr[9]
port 180 nsew signal input
flabel metal2 s 5712 0 5824 800 0 FreeSans 448 90 0 0 io_wbs_clk
port 181 nsew signal input
flabel metal2 s 7056 0 7168 800 0 FreeSans 448 90 0 0 io_wbs_cyc
port 182 nsew signal input
flabel metal2 s 13776 0 13888 800 0 FreeSans 448 90 0 0 io_wbs_datrd[0]
port 183 nsew signal tristate
flabel metal2 s 59472 0 59584 800 0 FreeSans 448 90 0 0 io_wbs_datrd[10]
port 184 nsew signal tristate
flabel metal2 s 63504 0 63616 800 0 FreeSans 448 90 0 0 io_wbs_datrd[11]
port 185 nsew signal tristate
flabel metal2 s 67536 0 67648 800 0 FreeSans 448 90 0 0 io_wbs_datrd[12]
port 186 nsew signal tristate
flabel metal2 s 71568 0 71680 800 0 FreeSans 448 90 0 0 io_wbs_datrd[13]
port 187 nsew signal tristate
flabel metal2 s 75600 0 75712 800 0 FreeSans 448 90 0 0 io_wbs_datrd[14]
port 188 nsew signal tristate
flabel metal2 s 79632 0 79744 800 0 FreeSans 448 90 0 0 io_wbs_datrd[15]
port 189 nsew signal tristate
flabel metal2 s 83664 0 83776 800 0 FreeSans 448 90 0 0 io_wbs_datrd[16]
port 190 nsew signal tristate
flabel metal2 s 87696 0 87808 800 0 FreeSans 448 90 0 0 io_wbs_datrd[17]
port 191 nsew signal tristate
flabel metal2 s 91728 0 91840 800 0 FreeSans 448 90 0 0 io_wbs_datrd[18]
port 192 nsew signal tristate
flabel metal2 s 95760 0 95872 800 0 FreeSans 448 90 0 0 io_wbs_datrd[19]
port 193 nsew signal tristate
flabel metal2 s 19152 0 19264 800 0 FreeSans 448 90 0 0 io_wbs_datrd[1]
port 194 nsew signal tristate
flabel metal2 s 99792 0 99904 800 0 FreeSans 448 90 0 0 io_wbs_datrd[20]
port 195 nsew signal tristate
flabel metal2 s 103824 0 103936 800 0 FreeSans 448 90 0 0 io_wbs_datrd[21]
port 196 nsew signal tristate
flabel metal2 s 107856 0 107968 800 0 FreeSans 448 90 0 0 io_wbs_datrd[22]
port 197 nsew signal tristate
flabel metal2 s 111888 0 112000 800 0 FreeSans 448 90 0 0 io_wbs_datrd[23]
port 198 nsew signal tristate
flabel metal2 s 115920 0 116032 800 0 FreeSans 448 90 0 0 io_wbs_datrd[24]
port 199 nsew signal tristate
flabel metal2 s 119952 0 120064 800 0 FreeSans 448 90 0 0 io_wbs_datrd[25]
port 200 nsew signal tristate
flabel metal2 s 123984 0 124096 800 0 FreeSans 448 90 0 0 io_wbs_datrd[26]
port 201 nsew signal tristate
flabel metal2 s 128016 0 128128 800 0 FreeSans 448 90 0 0 io_wbs_datrd[27]
port 202 nsew signal tristate
flabel metal2 s 132048 0 132160 800 0 FreeSans 448 90 0 0 io_wbs_datrd[28]
port 203 nsew signal tristate
flabel metal2 s 136080 0 136192 800 0 FreeSans 448 90 0 0 io_wbs_datrd[29]
port 204 nsew signal tristate
flabel metal2 s 24528 0 24640 800 0 FreeSans 448 90 0 0 io_wbs_datrd[2]
port 205 nsew signal tristate
flabel metal2 s 140112 0 140224 800 0 FreeSans 448 90 0 0 io_wbs_datrd[30]
port 206 nsew signal tristate
flabel metal2 s 144144 0 144256 800 0 FreeSans 448 90 0 0 io_wbs_datrd[31]
port 207 nsew signal tristate
flabel metal2 s 29904 0 30016 800 0 FreeSans 448 90 0 0 io_wbs_datrd[3]
port 208 nsew signal tristate
flabel metal2 s 35280 0 35392 800 0 FreeSans 448 90 0 0 io_wbs_datrd[4]
port 209 nsew signal tristate
flabel metal2 s 39312 0 39424 800 0 FreeSans 448 90 0 0 io_wbs_datrd[5]
port 210 nsew signal tristate
flabel metal2 s 43344 0 43456 800 0 FreeSans 448 90 0 0 io_wbs_datrd[6]
port 211 nsew signal tristate
flabel metal2 s 47376 0 47488 800 0 FreeSans 448 90 0 0 io_wbs_datrd[7]
port 212 nsew signal tristate
flabel metal2 s 51408 0 51520 800 0 FreeSans 448 90 0 0 io_wbs_datrd[8]
port 213 nsew signal tristate
flabel metal2 s 55440 0 55552 800 0 FreeSans 448 90 0 0 io_wbs_datrd[9]
port 214 nsew signal tristate
flabel metal2 s 15120 0 15232 800 0 FreeSans 448 90 0 0 io_wbs_datwr[0]
port 215 nsew signal input
flabel metal2 s 60816 0 60928 800 0 FreeSans 448 90 0 0 io_wbs_datwr[10]
port 216 nsew signal input
flabel metal2 s 64848 0 64960 800 0 FreeSans 448 90 0 0 io_wbs_datwr[11]
port 217 nsew signal input
flabel metal2 s 68880 0 68992 800 0 FreeSans 448 90 0 0 io_wbs_datwr[12]
port 218 nsew signal input
flabel metal2 s 72912 0 73024 800 0 FreeSans 448 90 0 0 io_wbs_datwr[13]
port 219 nsew signal input
flabel metal2 s 76944 0 77056 800 0 FreeSans 448 90 0 0 io_wbs_datwr[14]
port 220 nsew signal input
flabel metal2 s 80976 0 81088 800 0 FreeSans 448 90 0 0 io_wbs_datwr[15]
port 221 nsew signal input
flabel metal2 s 85008 0 85120 800 0 FreeSans 448 90 0 0 io_wbs_datwr[16]
port 222 nsew signal input
flabel metal2 s 89040 0 89152 800 0 FreeSans 448 90 0 0 io_wbs_datwr[17]
port 223 nsew signal input
flabel metal2 s 93072 0 93184 800 0 FreeSans 448 90 0 0 io_wbs_datwr[18]
port 224 nsew signal input
flabel metal2 s 97104 0 97216 800 0 FreeSans 448 90 0 0 io_wbs_datwr[19]
port 225 nsew signal input
flabel metal2 s 20496 0 20608 800 0 FreeSans 448 90 0 0 io_wbs_datwr[1]
port 226 nsew signal input
flabel metal2 s 101136 0 101248 800 0 FreeSans 448 90 0 0 io_wbs_datwr[20]
port 227 nsew signal input
flabel metal2 s 105168 0 105280 800 0 FreeSans 448 90 0 0 io_wbs_datwr[21]
port 228 nsew signal input
flabel metal2 s 109200 0 109312 800 0 FreeSans 448 90 0 0 io_wbs_datwr[22]
port 229 nsew signal input
flabel metal2 s 113232 0 113344 800 0 FreeSans 448 90 0 0 io_wbs_datwr[23]
port 230 nsew signal input
flabel metal2 s 117264 0 117376 800 0 FreeSans 448 90 0 0 io_wbs_datwr[24]
port 231 nsew signal input
flabel metal2 s 121296 0 121408 800 0 FreeSans 448 90 0 0 io_wbs_datwr[25]
port 232 nsew signal input
flabel metal2 s 125328 0 125440 800 0 FreeSans 448 90 0 0 io_wbs_datwr[26]
port 233 nsew signal input
flabel metal2 s 129360 0 129472 800 0 FreeSans 448 90 0 0 io_wbs_datwr[27]
port 234 nsew signal input
flabel metal2 s 133392 0 133504 800 0 FreeSans 448 90 0 0 io_wbs_datwr[28]
port 235 nsew signal input
flabel metal2 s 137424 0 137536 800 0 FreeSans 448 90 0 0 io_wbs_datwr[29]
port 236 nsew signal input
flabel metal2 s 25872 0 25984 800 0 FreeSans 448 90 0 0 io_wbs_datwr[2]
port 237 nsew signal input
flabel metal2 s 141456 0 141568 800 0 FreeSans 448 90 0 0 io_wbs_datwr[30]
port 238 nsew signal input
flabel metal2 s 145488 0 145600 800 0 FreeSans 448 90 0 0 io_wbs_datwr[31]
port 239 nsew signal input
flabel metal2 s 31248 0 31360 800 0 FreeSans 448 90 0 0 io_wbs_datwr[3]
port 240 nsew signal input
flabel metal2 s 36624 0 36736 800 0 FreeSans 448 90 0 0 io_wbs_datwr[4]
port 241 nsew signal input
flabel metal2 s 40656 0 40768 800 0 FreeSans 448 90 0 0 io_wbs_datwr[5]
port 242 nsew signal input
flabel metal2 s 44688 0 44800 800 0 FreeSans 448 90 0 0 io_wbs_datwr[6]
port 243 nsew signal input
flabel metal2 s 48720 0 48832 800 0 FreeSans 448 90 0 0 io_wbs_datwr[7]
port 244 nsew signal input
flabel metal2 s 52752 0 52864 800 0 FreeSans 448 90 0 0 io_wbs_datwr[8]
port 245 nsew signal input
flabel metal2 s 56784 0 56896 800 0 FreeSans 448 90 0 0 io_wbs_datwr[9]
port 246 nsew signal input
flabel metal2 s 8400 0 8512 800 0 FreeSans 448 90 0 0 io_wbs_rst
port 247 nsew signal input
flabel metal2 s 16464 0 16576 800 0 FreeSans 448 90 0 0 io_wbs_sel[0]
port 248 nsew signal input
flabel metal2 s 21840 0 21952 800 0 FreeSans 448 90 0 0 io_wbs_sel[1]
port 249 nsew signal input
flabel metal2 s 27216 0 27328 800 0 FreeSans 448 90 0 0 io_wbs_sel[2]
port 250 nsew signal input
flabel metal2 s 32592 0 32704 800 0 FreeSans 448 90 0 0 io_wbs_sel[3]
port 251 nsew signal input
flabel metal2 s 9744 0 9856 800 0 FreeSans 448 90 0 0 io_wbs_stb
port 252 nsew signal input
flabel metal2 s 11088 0 11200 800 0 FreeSans 448 90 0 0 io_wbs_we
port 253 nsew signal input
flabel metal4 s 19594 3076 19914 36908 0 FreeSans 1280 90 0 0 vdd
port 254 nsew power bidirectional
flabel metal4 s 56414 3076 56734 36908 0 FreeSans 1280 90 0 0 vdd
port 254 nsew power bidirectional
flabel metal4 s 93234 3076 93554 36908 0 FreeSans 1280 90 0 0 vdd
port 254 nsew power bidirectional
flabel metal4 s 130054 3076 130374 36908 0 FreeSans 1280 90 0 0 vdd
port 254 nsew power bidirectional
flabel metal4 s 38004 3076 38324 36908 0 FreeSans 1280 90 0 0 vss
port 255 nsew ground bidirectional
flabel metal4 s 74824 3076 75144 36908 0 FreeSans 1280 90 0 0 vss
port 255 nsew ground bidirectional
flabel metal4 s 111644 3076 111964 36908 0 FreeSans 1280 90 0 0 vss
port 255 nsew ground bidirectional
flabel metal4 s 148464 3076 148784 36908 0 FreeSans 1280 90 0 0 vss
port 255 nsew ground bidirectional
flabel metal2 s 5488 39200 5600 40000 0 FreeSans 448 90 0 0 web_mem0
port 256 nsew signal tristate
flabel metal2 s 76272 39200 76384 40000 0 FreeSans 448 90 0 0 web_mem1
port 257 nsew signal tristate
flabel metal2 s 9072 39200 9184 40000 0 FreeSans 448 90 0 0 wmask_mem0[0]
port 258 nsew signal tristate
flabel metal2 s 12656 39200 12768 40000 0 FreeSans 448 90 0 0 wmask_mem0[1]
port 259 nsew signal tristate
flabel metal2 s 16240 39200 16352 40000 0 FreeSans 448 90 0 0 wmask_mem0[2]
port 260 nsew signal tristate
flabel metal2 s 19824 39200 19936 40000 0 FreeSans 448 90 0 0 wmask_mem0[3]
port 261 nsew signal tristate
flabel metal2 s 79856 39200 79968 40000 0 FreeSans 448 90 0 0 wmask_mem1[0]
port 262 nsew signal tristate
flabel metal2 s 83440 39200 83552 40000 0 FreeSans 448 90 0 0 wmask_mem1[1]
port 263 nsew signal tristate
flabel metal2 s 87024 39200 87136 40000 0 FreeSans 448 90 0 0 wmask_mem1[2]
port 264 nsew signal tristate
flabel metal2 s 90608 39200 90720 40000 0 FreeSans 448 90 0 0 wmask_mem1[3]
port 265 nsew signal tristate
rlabel metal1 74984 36848 74984 36848 0 vdd
rlabel via1 75064 36064 75064 36064 0 vss
rlabel metal2 8120 6384 8120 6384 0 _000_
rlabel metal2 7896 4368 7896 4368 0 _001_
rlabel metal3 21000 4872 21000 4872 0 _002_
rlabel metal2 19208 6272 19208 6272 0 _003_
rlabel metal2 28168 4704 28168 4704 0 _004_
rlabel metal2 30968 5712 30968 5712 0 _005_
rlabel metal2 38248 5320 38248 5320 0 _006_
rlabel metal2 38584 4816 38584 4816 0 _007_
rlabel metal2 48328 4704 48328 4704 0 _008_
rlabel metal2 49896 5040 49896 5040 0 _009_
rlabel metal2 64232 5880 64232 5880 0 _010_
rlabel metal3 67368 6440 67368 6440 0 _011_
rlabel metal3 70672 5992 70672 5992 0 _012_
rlabel metal2 68488 4648 68488 4648 0 _013_
rlabel metal2 77112 4872 77112 4872 0 _014_
rlabel metal2 80248 4312 80248 4312 0 _015_
rlabel metal2 92120 4704 92120 4704 0 _016_
rlabel metal2 88424 5040 88424 5040 0 _017_
rlabel metal2 97944 4704 97944 4704 0 _018_
rlabel metal2 102088 4704 102088 4704 0 _019_
rlabel metal2 120064 4312 120064 4312 0 _020_
rlabel metal2 116312 5376 116312 5376 0 _021_
rlabel metal3 133560 8008 133560 8008 0 _022_
rlabel metal2 133672 7112 133672 7112 0 _023_
rlabel metal3 129696 3752 129696 3752 0 _024_
rlabel metal3 132888 3752 132888 3752 0 _025_
rlabel metal2 111664 3752 111664 3752 0 _026_
rlabel metal2 116200 4144 116200 4144 0 _027_
rlabel metal2 119672 3752 119672 3752 0 _028_
rlabel metal2 115472 3752 115472 3752 0 _029_
rlabel metal2 131880 5096 131880 5096 0 _030_
rlabel metal3 132552 6104 132552 6104 0 _031_
rlabel metal2 130984 4984 130984 4984 0 _032_
rlabel metal2 130984 6496 130984 6496 0 _033_
rlabel metal2 16072 4704 16072 4704 0 _034_
rlabel metal3 10976 5096 10976 5096 0 _035_
rlabel metal3 11200 4536 11200 4536 0 _036_
rlabel metal2 16968 5768 16968 5768 0 _037_
rlabel metal3 16408 6104 16408 6104 0 _038_
rlabel metal2 25704 5768 25704 5768 0 _039_
rlabel metal2 28392 6720 28392 6720 0 _040_
rlabel metal3 40096 5992 40096 5992 0 _041_
rlabel metal2 36120 4592 36120 4592 0 _042_
rlabel metal2 45864 5152 45864 5152 0 _043_
rlabel metal2 52248 5768 52248 5768 0 _044_
rlabel metal2 61768 4704 61768 4704 0 _045_
rlabel metal2 62944 6664 62944 6664 0 _046_
rlabel metal2 67704 6720 67704 6720 0 _047_
rlabel metal3 65240 6552 65240 6552 0 _048_
rlabel metal2 79352 6160 79352 6160 0 _049_
rlabel metal2 76104 5768 76104 5768 0 _050_
rlabel metal2 89712 5992 89712 5992 0 _051_
rlabel metal2 85960 5544 85960 5544 0 _052_
rlabel metal3 93744 5992 93744 5992 0 _053_
rlabel metal2 99624 5936 99624 5936 0 _054_
rlabel metal2 117712 5096 117712 5096 0 _055_
rlabel metal3 120736 5880 120736 5880 0 _056_
rlabel metal2 143808 3304 143808 3304 0 _057_
rlabel metal2 143696 4536 143696 4536 0 _058_
rlabel metal2 128576 3640 128576 3640 0 _059_
rlabel metal2 135912 4816 135912 4816 0 _060_
rlabel metal2 108360 4592 108360 4592 0 _061_
rlabel metal3 112504 4872 112504 4872 0 _062_
rlabel metal2 119000 5600 119000 5600 0 _063_
rlabel metal2 112392 5544 112392 5544 0 _064_
rlabel metal2 141512 5992 141512 5992 0 _065_
rlabel metal2 142408 7448 142408 7448 0 _066_
rlabel metal2 127736 7448 127736 7448 0 _067_
rlabel metal2 128408 7532 128408 7532 0 _068_
rlabel metal3 52248 31752 52248 31752 0 _069_
rlabel metal3 127792 9912 127792 9912 0 _070_
rlabel metal3 141120 5880 141120 5880 0 _071_
rlabel metal2 142520 7000 142520 7000 0 _072_
rlabel metal3 128632 9016 128632 9016 0 _073_
rlabel metal2 127400 7056 127400 7056 0 _074_
rlabel metal2 127064 7896 127064 7896 0 _075_
rlabel metal2 22120 33040 22120 33040 0 _076_
rlabel metal2 141848 33208 141848 33208 0 _077_
rlabel metal3 144144 5992 144144 5992 0 _078_
rlabel metal3 143192 6104 143192 6104 0 _079_
rlabel metal2 142240 6888 142240 6888 0 _080_
rlabel metal2 141848 7168 141848 7168 0 _081_
rlabel metal3 115080 6776 115080 6776 0 _082_
rlabel metal3 118888 8120 118888 8120 0 _083_
rlabel metal3 113064 5992 113064 5992 0 _084_
rlabel metal3 119896 8232 119896 8232 0 _085_
rlabel metal2 119336 5264 119336 5264 0 _086_
rlabel metal3 139160 34776 139160 34776 0 _087_
rlabel metal3 115024 5992 115024 5992 0 _088_
rlabel metal2 111048 5320 111048 5320 0 _089_
rlabel metal3 107576 6104 107576 6104 0 _090_
rlabel metal2 108136 5544 108136 5544 0 _091_
rlabel metal3 139272 5208 139272 5208 0 _092_
rlabel metal2 145208 4760 145208 4760 0 _093_
rlabel metal2 136248 4816 136248 4816 0 _094_
rlabel metal3 139832 6104 139832 6104 0 _095_
rlabel metal2 137368 5320 137368 5320 0 _096_
rlabel metal2 75096 33936 75096 33936 0 _097_
rlabel metal2 102760 35840 102760 35840 0 _098_
rlabel metal3 146888 5208 146888 5208 0 _099_
rlabel metal2 144144 4424 144144 4424 0 _100_
rlabel metal3 146664 6104 146664 6104 0 _101_
rlabel metal3 144592 3528 144592 3528 0 _102_
rlabel metal3 122696 7448 122696 7448 0 _103_
rlabel metal2 50344 6272 50344 6272 0 _104_
rlabel metal2 100296 7000 100296 7000 0 _105_
rlabel metal2 122136 6944 122136 6944 0 _106_
rlabel metal2 121464 7728 121464 7728 0 _107_
rlabel metal2 118776 7448 118776 7448 0 _108_
rlabel metal3 99792 35672 99792 35672 0 _109_
rlabel metal2 101080 6776 101080 6776 0 _110_
rlabel metal2 99232 6888 99232 6888 0 _111_
rlabel metal2 90440 7112 90440 7112 0 _112_
rlabel metal2 91560 6048 91560 6048 0 _113_
rlabel metal2 88032 7448 88032 7448 0 _114_
rlabel metal2 77896 7280 77896 7280 0 _115_
rlabel metal2 86520 6216 86520 6216 0 _116_
rlabel metal3 92624 7672 92624 7672 0 _117_
rlabel metal2 89488 5880 89488 5880 0 _118_
rlabel metal2 76216 34720 76216 34720 0 _119_
rlabel metal2 75488 7336 75488 7336 0 _120_
rlabel metal2 75768 6328 75768 6328 0 _121_
rlabel metal3 77672 7448 77672 7448 0 _122_
rlabel metal2 78232 6944 78232 6944 0 _123_
rlabel metal2 67760 5320 67760 5320 0 _124_
rlabel metal2 67928 5768 67928 5768 0 _125_
rlabel metal2 67368 5656 67368 5656 0 _126_
rlabel metal2 69496 7112 69496 7112 0 _127_
rlabel metal2 68488 7168 68488 7168 0 _128_
rlabel metal2 49560 34832 49560 34832 0 _129_
rlabel metal2 65856 7448 65856 7448 0 _130_
rlabel metal3 64736 7448 64736 7448 0 _131_
rlabel metal2 65968 9016 65968 9016 0 _132_
rlabel metal3 64232 8792 64232 8792 0 _133_
rlabel metal2 50176 6888 50176 6888 0 _134_
rlabel metal2 48104 6496 48104 6496 0 _135_
rlabel metal3 51352 6552 51352 6552 0 _136_
rlabel metal3 48328 7448 48328 7448 0 _137_
rlabel metal3 47264 5992 47264 5992 0 _138_
rlabel metal2 30856 33992 30856 33992 0 _139_
rlabel metal3 38584 7336 38584 7336 0 _140_
rlabel metal2 36792 5320 36792 5320 0 _141_
rlabel metal2 40208 6776 40208 6776 0 _142_
rlabel metal2 39480 6160 39480 6160 0 _143_
rlabel metal2 31584 6664 31584 6664 0 _144_
rlabel metal3 29568 6552 29568 6552 0 _145_
rlabel metal2 29736 6944 29736 6944 0 _146_
rlabel metal3 28168 7336 28168 7336 0 _147_
rlabel metal2 26488 6552 26488 6552 0 _148_
rlabel metal2 21056 35448 21056 35448 0 _149_
rlabel metal3 17136 5880 17136 5880 0 _150_
rlabel metal3 19264 7672 19264 7672 0 _151_
rlabel metal2 16632 6608 16632 6608 0 _152_
rlabel metal3 12320 3416 12320 3416 0 _153_
rlabel metal2 9688 4816 9688 4816 0 _154_
rlabel metal2 52752 35112 52752 35112 0 _155_
rlabel metal2 50232 34384 50232 34384 0 _156_
rlabel metal2 59864 4144 59864 4144 0 _157_
rlabel metal2 29512 3640 29512 3640 0 _158_
rlabel metal2 29288 3696 29288 3696 0 _159_
rlabel metal3 71736 4984 71736 4984 0 _160_
rlabel metal3 48384 5096 48384 5096 0 _161_
rlabel metal2 69496 5936 69496 5936 0 _162_
rlabel metal3 92680 5208 92680 5208 0 _163_
rlabel metal2 97832 4816 97832 4816 0 _164_
rlabel metal3 134344 4536 134344 4536 0 _165_
rlabel metal3 117880 3416 117880 3416 0 _166_
rlabel metal2 132160 6552 132160 6552 0 _167_
rlabel metal2 6440 37394 6440 37394 0 addr_mem0[0]
rlabel metal3 10136 35000 10136 35000 0 addr_mem0[1]
rlabel metal2 13888 35000 13888 35000 0 addr_mem0[2]
rlabel metal2 17192 37114 17192 37114 0 addr_mem0[3]
rlabel metal2 21896 35056 21896 35056 0 addr_mem0[4]
rlabel metal2 23632 35000 23632 35000 0 addr_mem0[5]
rlabel metal2 26152 37114 26152 37114 0 addr_mem0[6]
rlabel metal2 28168 35056 28168 35056 0 addr_mem0[7]
rlabel metal2 31752 35056 31752 35056 0 addr_mem0[8]
rlabel metal2 77224 38010 77224 38010 0 addr_mem1[0]
rlabel metal2 82600 35056 82600 35056 0 addr_mem1[1]
rlabel metal2 84392 37170 84392 37170 0 addr_mem1[2]
rlabel metal3 88592 33432 88592 33432 0 addr_mem1[3]
rlabel metal2 93352 35056 93352 35056 0 addr_mem1[4]
rlabel metal2 95816 35056 95816 35056 0 addr_mem1[5]
rlabel metal2 96936 36610 96936 36610 0 addr_mem1[6]
rlabel metal3 100016 33992 100016 33992 0 addr_mem1[7]
rlabel metal2 102312 37002 102312 37002 0 addr_mem1[8]
rlabel metal3 68936 4312 68936 4312 0 clknet_0_io_wbs_clk
rlabel metal3 29960 5880 29960 5880 0 clknet_2_0__leaf_io_wbs_clk
rlabel metal2 7448 6552 7448 6552 0 clknet_2_1__leaf_io_wbs_clk
rlabel metal2 76720 3640 76720 3640 0 clknet_2_2__leaf_io_wbs_clk
rlabel metal3 99288 4312 99288 4312 0 clknet_2_3__leaf_io_wbs_clk
rlabel metal2 7336 37170 7336 37170 0 din_mem0[0]
rlabel metal2 36008 37114 36008 37114 0 din_mem0[10]
rlabel metal2 37968 34216 37968 34216 0 din_mem0[11]
rlabel metal2 39928 36008 39928 36008 0 din_mem0[12]
rlabel metal2 41832 36008 41832 36008 0 din_mem0[13]
rlabel metal2 43512 36008 43512 36008 0 din_mem0[14]
rlabel metal2 45248 34216 45248 34216 0 din_mem0[15]
rlabel metal2 47040 34216 47040 34216 0 din_mem0[16]
rlabel metal3 49112 34216 49112 34216 0 din_mem0[17]
rlabel metal3 50624 35000 50624 35000 0 din_mem0[18]
rlabel metal2 52416 34216 52416 34216 0 din_mem0[19]
rlabel metal2 10976 35560 10976 35560 0 din_mem0[1]
rlabel metal2 54096 35000 54096 35000 0 din_mem0[20]
rlabel metal2 55608 36456 55608 36456 0 din_mem0[21]
rlabel metal2 57736 36008 57736 36008 0 din_mem0[22]
rlabel metal2 59472 35000 59472 35000 0 din_mem0[23]
rlabel metal2 61432 35392 61432 35392 0 din_mem0[24]
rlabel metal2 62944 35000 62944 35000 0 din_mem0[25]
rlabel metal2 65016 35112 65016 35112 0 din_mem0[26]
rlabel metal2 66472 36610 66472 36610 0 din_mem0[27]
rlabel metal2 69944 34272 69944 34272 0 din_mem0[28]
rlabel metal2 70392 36008 70392 36008 0 din_mem0[29]
rlabel metal2 14560 35560 14560 35560 0 din_mem0[2]
rlabel metal2 72240 35000 72240 35000 0 din_mem0[30]
rlabel metal3 74088 35000 74088 35000 0 din_mem0[31]
rlabel metal2 17808 35784 17808 35784 0 din_mem0[3]
rlabel metal2 21840 35784 21840 35784 0 din_mem0[4]
rlabel metal2 24304 35560 24304 35560 0 din_mem0[5]
rlabel metal2 26824 35896 26824 35896 0 din_mem0[6]
rlabel metal2 29960 35392 29960 35392 0 din_mem0[7]
rlabel metal2 32424 37114 32424 37114 0 din_mem0[8]
rlabel metal2 34216 37114 34216 37114 0 din_mem0[9]
rlabel metal2 78456 36176 78456 36176 0 din_mem1[0]
rlabel metal3 107240 33992 107240 33992 0 din_mem1[10]
rlabel metal2 108584 37170 108584 37170 0 din_mem1[11]
rlabel metal2 111608 35056 111608 35056 0 din_mem1[12]
rlabel metal2 113064 33488 113064 33488 0 din_mem1[13]
rlabel metal2 115528 35056 115528 35056 0 din_mem1[14]
rlabel metal3 116200 33992 116200 33992 0 din_mem1[15]
rlabel metal2 118440 35112 118440 35112 0 din_mem1[16]
rlabel metal2 119336 36610 119336 36610 0 din_mem1[17]
rlabel metal2 121464 35112 121464 35112 0 din_mem1[18]
rlabel metal3 123368 33992 123368 33992 0 din_mem1[19]
rlabel metal2 82712 34160 82712 34160 0 din_mem1[1]
rlabel metal2 125160 36064 125160 36064 0 din_mem1[20]
rlabel metal2 127736 35056 127736 35056 0 din_mem1[21]
rlabel metal2 128464 33432 128464 33432 0 din_mem1[22]
rlabel metal2 130536 33656 130536 33656 0 din_mem1[23]
rlabel metal2 133672 35056 133672 35056 0 din_mem1[24]
rlabel metal2 135688 35672 135688 35672 0 din_mem1[25]
rlabel metal2 136360 35056 136360 35056 0 din_mem1[26]
rlabel metal2 137256 36330 137256 36330 0 din_mem1[27]
rlabel metal2 140728 34552 140728 34552 0 din_mem1[28]
rlabel metal3 141288 35000 141288 35000 0 din_mem1[29]
rlabel metal2 85288 37506 85288 37506 0 din_mem1[2]
rlabel metal3 145096 36568 145096 36568 0 din_mem1[30]
rlabel metal3 145040 33992 145040 33992 0 din_mem1[31]
rlabel metal2 90776 33488 90776 33488 0 din_mem1[3]
rlabel metal2 95928 35224 95928 35224 0 din_mem1[4]
rlabel metal2 97608 35112 97608 35112 0 din_mem1[5]
rlabel metal2 99288 35056 99288 35056 0 din_mem1[6]
rlabel metal2 101864 35056 101864 35056 0 din_mem1[7]
rlabel metal2 103880 34216 103880 34216 0 din_mem1[8]
rlabel metal3 105448 33992 105448 33992 0 din_mem1[9]
rlabel metal2 7896 36792 7896 36792 0 dout_mem0[0]
rlabel metal2 37072 35784 37072 35784 0 dout_mem0[10]
rlabel metal2 38920 36848 38920 36848 0 dout_mem0[11]
rlabel metal2 41720 36232 41720 36232 0 dout_mem0[12]
rlabel metal2 42448 36344 42448 36344 0 dout_mem0[13]
rlabel metal2 43848 36064 43848 36064 0 dout_mem0[14]
rlabel metal2 46200 36232 46200 36232 0 dout_mem0[15]
rlabel metal3 47264 36344 47264 36344 0 dout_mem0[16]
rlabel metal2 49784 36344 49784 36344 0 dout_mem0[17]
rlabel metal2 51016 36848 51016 36848 0 dout_mem0[18]
rlabel metal2 53200 35784 53200 35784 0 dout_mem0[19]
rlabel metal2 11760 36344 11760 36344 0 dout_mem0[1]
rlabel metal2 54824 37786 54824 37786 0 dout_mem0[20]
rlabel metal3 57232 35784 57232 35784 0 dout_mem0[21]
rlabel metal2 58464 36344 58464 36344 0 dout_mem0[22]
rlabel metal2 60368 35784 60368 35784 0 dout_mem0[23]
rlabel metal2 62328 35784 62328 35784 0 dout_mem0[24]
rlabel metal3 64120 31864 64120 31864 0 dout_mem0[25]
rlabel metal3 63392 36344 63392 36344 0 dout_mem0[26]
rlabel metal2 67536 36568 67536 36568 0 dout_mem0[27]
rlabel metal2 69328 36344 69328 36344 0 dout_mem0[28]
rlabel metal2 71288 37296 71288 37296 0 dout_mem0[29]
rlabel metal2 15400 37786 15400 37786 0 dout_mem0[2]
rlabel metal2 73472 35784 73472 35784 0 dout_mem0[30]
rlabel metal2 74536 37786 74536 37786 0 dout_mem0[31]
rlabel metal2 19320 36400 19320 36400 0 dout_mem0[3]
rlabel metal3 22736 36344 22736 36344 0 dout_mem0[4]
rlabel metal2 25592 36400 25592 36400 0 dout_mem0[5]
rlabel metal2 28280 36176 28280 36176 0 dout_mem0[6]
rlabel metal2 30968 36848 30968 36848 0 dout_mem0[7]
rlabel metal2 33544 35784 33544 35784 0 dout_mem0[8]
rlabel metal2 35112 37786 35112 37786 0 dout_mem0[9]
rlabel metal3 80192 36344 80192 36344 0 dout_mem1[0]
rlabel metal3 108304 36344 108304 36344 0 dout_mem1[10]
rlabel metal3 110208 35784 110208 35784 0 dout_mem1[11]
rlabel metal3 111944 36344 111944 36344 0 dout_mem1[12]
rlabel metal3 113680 35784 113680 35784 0 dout_mem1[13]
rlabel metal3 115696 36344 115696 36344 0 dout_mem1[14]
rlabel metal2 117880 35448 117880 35448 0 dout_mem1[15]
rlabel metal2 120456 36512 120456 36512 0 dout_mem1[16]
rlabel metal2 120344 35448 120344 35448 0 dout_mem1[17]
rlabel metal3 123200 36344 123200 36344 0 dout_mem1[18]
rlabel metal2 124432 35784 124432 35784 0 dout_mem1[19]
rlabel metal2 83832 36568 83832 36568 0 dout_mem1[1]
rlabel metal2 126112 35784 126112 35784 0 dout_mem1[20]
rlabel metal2 127680 36344 127680 36344 0 dout_mem1[21]
rlabel metal2 129360 35784 129360 35784 0 dout_mem1[22]
rlabel metal2 131152 36344 131152 36344 0 dout_mem1[23]
rlabel metal2 133952 35784 133952 35784 0 dout_mem1[24]
rlabel via2 135352 36344 135352 36344 0 dout_mem1[25]
rlabel metal2 138040 35560 138040 35560 0 dout_mem1[26]
rlabel metal3 139104 36344 139104 36344 0 dout_mem1[27]
rlabel metal2 140280 36344 140280 36344 0 dout_mem1[28]
rlabel metal2 142800 36344 142800 36344 0 dout_mem1[29]
rlabel metal2 86856 36400 86856 36400 0 dout_mem1[2]
rlabel metal2 143416 35000 143416 35000 0 dout_mem1[30]
rlabel metal2 146216 36232 146216 36232 0 dout_mem1[31]
rlabel metal3 90328 36344 90328 36344 0 dout_mem1[3]
rlabel metal2 94584 36624 94584 36624 0 dout_mem1[4]
rlabel metal3 98280 36344 98280 36344 0 dout_mem1[5]
rlabel metal2 100856 36400 100856 36400 0 dout_mem1[6]
rlabel metal2 102424 35336 102424 35336 0 dout_mem1[7]
rlabel metal3 104720 36344 104720 36344 0 dout_mem1[8]
rlabel metal3 106512 35784 106512 35784 0 dout_mem1[9]
rlabel metal2 4424 2478 4424 2478 0 io_wbs_ack
rlabel metal2 58072 3416 58072 3416 0 io_wbs_adr[10]
rlabel metal2 61936 3416 61936 3416 0 io_wbs_adr[11]
rlabel metal3 23688 3416 23688 3416 0 io_wbs_adr[2]
rlabel metal2 28952 3920 28952 3920 0 io_wbs_adr[3]
rlabel metal2 33880 4872 33880 4872 0 io_wbs_adr[4]
rlabel metal2 37800 2856 37800 2856 0 io_wbs_adr[5]
rlabel metal2 41944 3416 41944 3416 0 io_wbs_adr[6]
rlabel metal2 45976 3416 45976 3416 0 io_wbs_adr[7]
rlabel metal2 50008 3416 50008 3416 0 io_wbs_adr[8]
rlabel metal2 54040 3416 54040 3416 0 io_wbs_adr[9]
rlabel metal2 5768 1638 5768 1638 0 io_wbs_clk
rlabel metal2 6832 4200 6832 4200 0 io_wbs_cyc
rlabel metal2 13832 2870 13832 2870 0 io_wbs_datrd[0]
rlabel metal2 59528 2310 59528 2310 0 io_wbs_datrd[10]
rlabel metal2 63560 3262 63560 3262 0 io_wbs_datrd[11]
rlabel metal2 67592 2926 67592 2926 0 io_wbs_datrd[12]
rlabel metal2 71624 2478 71624 2478 0 io_wbs_datrd[13]
rlabel metal2 75656 2086 75656 2086 0 io_wbs_datrd[14]
rlabel metal2 79688 3654 79688 3654 0 io_wbs_datrd[15]
rlabel metal2 83720 2478 83720 2478 0 io_wbs_datrd[16]
rlabel metal2 87752 2478 87752 2478 0 io_wbs_datrd[17]
rlabel metal2 91784 2478 91784 2478 0 io_wbs_datrd[18]
rlabel metal2 95816 2478 95816 2478 0 io_wbs_datrd[19]
rlabel metal2 19208 2478 19208 2478 0 io_wbs_datrd[1]
rlabel metal2 99848 1806 99848 1806 0 io_wbs_datrd[20]
rlabel metal2 103880 2926 103880 2926 0 io_wbs_datrd[21]
rlabel metal2 107912 2926 107912 2926 0 io_wbs_datrd[22]
rlabel metal2 111944 854 111944 854 0 io_wbs_datrd[23]
rlabel metal2 115976 2478 115976 2478 0 io_wbs_datrd[24]
rlabel metal2 120008 1414 120008 1414 0 io_wbs_datrd[25]
rlabel metal2 124040 2086 124040 2086 0 io_wbs_datrd[26]
rlabel metal2 128072 1806 128072 1806 0 io_wbs_datrd[27]
rlabel metal2 132104 2478 132104 2478 0 io_wbs_datrd[28]
rlabel metal2 136136 2086 136136 2086 0 io_wbs_datrd[29]
rlabel metal2 24584 3262 24584 3262 0 io_wbs_datrd[2]
rlabel metal2 140168 2198 140168 2198 0 io_wbs_datrd[30]
rlabel metal2 144200 2198 144200 2198 0 io_wbs_datrd[31]
rlabel metal2 29960 2926 29960 2926 0 io_wbs_datrd[3]
rlabel metal2 35336 854 35336 854 0 io_wbs_datrd[4]
rlabel metal2 39368 2478 39368 2478 0 io_wbs_datrd[5]
rlabel metal2 43400 2870 43400 2870 0 io_wbs_datrd[6]
rlabel metal2 47432 3262 47432 3262 0 io_wbs_datrd[7]
rlabel metal2 51464 854 51464 854 0 io_wbs_datrd[8]
rlabel metal2 55496 2478 55496 2478 0 io_wbs_datrd[9]
rlabel metal3 15736 3416 15736 3416 0 io_wbs_datwr[0]
rlabel metal2 60536 4536 60536 4536 0 io_wbs_datwr[10]
rlabel metal2 65240 3472 65240 3472 0 io_wbs_datwr[11]
rlabel metal2 69832 3416 69832 3416 0 io_wbs_datwr[12]
rlabel metal2 73080 3416 73080 3416 0 io_wbs_datwr[13]
rlabel metal2 77336 3472 77336 3472 0 io_wbs_datwr[14]
rlabel metal3 81984 3416 81984 3416 0 io_wbs_datwr[15]
rlabel metal3 85960 3416 85960 3416 0 io_wbs_datwr[16]
rlabel metal3 91504 3416 91504 3416 0 io_wbs_datwr[17]
rlabel metal3 93912 3416 93912 3416 0 io_wbs_datwr[18]
rlabel metal2 97048 3416 97048 3416 0 io_wbs_datwr[19]
rlabel metal3 20832 4424 20832 4424 0 io_wbs_datwr[1]
rlabel metal2 101080 3416 101080 3416 0 io_wbs_datwr[20]
rlabel metal2 105112 3416 105112 3416 0 io_wbs_datwr[21]
rlabel metal2 109088 3416 109088 3416 0 io_wbs_datwr[22]
rlabel metal2 114632 3528 114632 3528 0 io_wbs_datwr[23]
rlabel metal2 118552 3472 118552 3472 0 io_wbs_datwr[24]
rlabel metal2 122136 2072 122136 2072 0 io_wbs_datwr[25]
rlabel metal2 125384 1246 125384 1246 0 io_wbs_datwr[26]
rlabel metal2 130312 3472 130312 3472 0 io_wbs_datwr[27]
rlabel metal2 133448 2086 133448 2086 0 io_wbs_datwr[28]
rlabel metal2 137480 2590 137480 2590 0 io_wbs_datwr[29]
rlabel metal2 25816 4200 25816 4200 0 io_wbs_datwr[2]
rlabel metal2 141400 4200 141400 4200 0 io_wbs_datwr[30]
rlabel metal2 145600 3416 145600 3416 0 io_wbs_datwr[31]
rlabel metal2 31304 2590 31304 2590 0 io_wbs_datwr[3]
rlabel metal2 36960 3416 36960 3416 0 io_wbs_datwr[4]
rlabel metal3 40992 3416 40992 3416 0 io_wbs_datwr[5]
rlabel metal3 45192 4984 45192 4984 0 io_wbs_datwr[6]
rlabel metal2 49224 2968 49224 2968 0 io_wbs_datwr[7]
rlabel metal2 52696 4200 52696 4200 0 io_wbs_datwr[8]
rlabel metal3 57232 4424 57232 4424 0 io_wbs_datwr[9]
rlabel metal2 8344 3976 8344 3976 0 io_wbs_rst
rlabel metal3 17080 3416 17080 3416 0 io_wbs_sel[0]
rlabel metal2 21896 2086 21896 2086 0 io_wbs_sel[1]
rlabel metal2 27272 2086 27272 2086 0 io_wbs_sel[2]
rlabel metal2 32480 3416 32480 3416 0 io_wbs_sel[3]
rlabel metal3 10416 4424 10416 4424 0 io_wbs_stb
rlabel metal2 12376 3472 12376 3472 0 io_wbs_we
rlabel metal2 17864 34552 17864 34552 0 net1
rlabel metal2 52080 36568 52080 36568 0 net10
rlabel metal2 74200 34608 74200 34608 0 net100
rlabel metal3 28728 4872 28728 4872 0 net101
rlabel metal2 31528 34720 31528 34720 0 net102
rlabel metal3 51016 27720 51016 27720 0 net103
rlabel metal2 47040 5208 47040 5208 0 net104
rlabel metal3 47936 4200 47936 4200 0 net105
rlabel metal2 46872 32760 46872 32760 0 net106
rlabel metal2 48328 32872 48328 32872 0 net107
rlabel metal2 8904 3416 8904 3416 0 net108
rlabel metal3 15176 6776 15176 6776 0 net109
rlabel metal2 54432 35560 54432 35560 0 net11
rlabel metal2 23744 4200 23744 4200 0 net110
rlabel metal2 28560 3640 28560 3640 0 net111
rlabel metal3 32088 3640 32088 3640 0 net112
rlabel metal2 10360 3360 10360 3360 0 net113
rlabel metal2 6440 3584 6440 3584 0 net114
rlabel metal2 7784 34496 7784 34496 0 net115
rlabel metal2 10920 34608 10920 34608 0 net116
rlabel metal3 15512 34328 15512 34328 0 net117
rlabel metal2 21896 36120 21896 36120 0 net118
rlabel metal2 22904 34552 22904 34552 0 net119
rlabel metal2 12824 36176 12824 36176 0 net12
rlabel metal2 25592 35448 25592 35448 0 net120
rlabel metal2 27048 35392 27048 35392 0 net121
rlabel metal2 28840 33656 28840 33656 0 net122
rlabel metal2 46088 34496 46088 34496 0 net123
rlabel metal2 30184 30464 30184 30464 0 net124
rlabel metal2 44632 32648 44632 32648 0 net125
rlabel metal2 51632 33432 51632 33432 0 net126
rlabel metal2 60816 34216 60816 34216 0 net127
rlabel metal3 76104 26264 76104 26264 0 net128
rlabel metal2 77784 34048 77784 34048 0 net129
rlabel metal3 90888 25704 90888 25704 0 net13
rlabel metal2 84504 36176 84504 36176 0 net130
rlabel metal2 100240 35000 100240 35000 0 net131
rlabel metal2 77224 32760 77224 32760 0 net132
rlabel metal2 6888 35616 6888 35616 0 net133
rlabel metal2 51240 33320 51240 33320 0 net134
rlabel metal2 45752 36120 45752 36120 0 net135
rlabel metal2 51464 33992 51464 33992 0 net136
rlabel metal2 53592 35672 53592 35672 0 net137
rlabel metal2 44632 36064 44632 36064 0 net138
rlabel metal2 46312 35112 46312 35112 0 net139
rlabel metal2 59024 35560 59024 35560 0 net14
rlabel metal2 48216 34216 48216 34216 0 net140
rlabel metal2 50792 34160 50792 34160 0 net141
rlabel metal2 52024 34832 52024 34832 0 net142
rlabel metal2 53592 33768 53592 33768 0 net143
rlabel metal2 10472 35952 10472 35952 0 net144
rlabel metal2 61320 35560 61320 35560 0 net145
rlabel metal2 56392 35672 56392 35672 0 net146
rlabel metal3 74032 23128 74032 23128 0 net147
rlabel metal2 99064 31444 99064 31444 0 net148
rlabel metal2 62552 35896 62552 35896 0 net149
rlabel metal3 98392 26824 98392 26824 0 net15
rlabel metal2 64120 36176 64120 36176 0 net150
rlabel metal3 67480 31864 67480 31864 0 net151
rlabel metal2 68208 33432 68208 33432 0 net152
rlabel metal2 71064 34048 71064 34048 0 net153
rlabel metal2 71736 34888 71736 34888 0 net154
rlabel metal2 14280 35672 14280 35672 0 net155
rlabel metal3 75768 34776 75768 34776 0 net156
rlabel metal2 73808 34328 73808 34328 0 net157
rlabel metal2 19208 35000 19208 35000 0 net158
rlabel metal2 23128 35616 23128 35616 0 net159
rlabel metal3 98840 24136 98840 24136 0 net16
rlabel metal2 24472 34384 24472 34384 0 net160
rlabel metal2 27608 35952 27608 35952 0 net161
rlabel metal2 31416 32704 31416 32704 0 net162
rlabel metal2 46424 33824 46424 33824 0 net163
rlabel metal2 47992 33376 47992 33376 0 net164
rlabel metal3 48776 29624 48776 29624 0 net165
rlabel metal2 82600 36736 82600 36736 0 net166
rlabel metal2 98056 34944 98056 34944 0 net167
rlabel metal2 104104 35616 104104 35616 0 net168
rlabel metal2 108248 33992 108248 33992 0 net169
rlabel metal2 63672 37184 63672 37184 0 net17
rlabel metal2 112056 35504 112056 35504 0 net170
rlabel metal2 115640 35728 115640 35728 0 net171
rlabel metal2 117824 36232 117824 36232 0 net172
rlabel metal2 120120 35168 120120 35168 0 net173
rlabel metal2 122584 34944 122584 34944 0 net174
rlabel metal2 108472 35560 108472 35560 0 net175
rlabel metal2 22232 32088 22232 32088 0 net176
rlabel metal2 113960 36064 113960 36064 0 net177
rlabel metal2 126616 33600 126616 33600 0 net178
rlabel metal2 129640 34776 129640 34776 0 net179
rlabel metal2 64680 34384 64680 34384 0 net18
rlabel metal2 131432 34552 131432 34552 0 net180
rlabel metal2 133000 34832 133000 34832 0 net181
rlabel metal2 132664 35000 132664 35000 0 net182
rlabel metal3 134792 34328 134792 34328 0 net183
rlabel metal2 135128 33992 135128 33992 0 net184
rlabel metal2 137480 35168 137480 35168 0 net185
rlabel metal2 139384 35504 139384 35504 0 net186
rlabel metal2 36568 29596 36568 29596 0 net187
rlabel metal3 144536 36344 144536 36344 0 net188
rlabel metal2 145040 36232 145040 36232 0 net189
rlabel metal2 67256 37464 67256 37464 0 net19
rlabel metal2 42504 30688 42504 30688 0 net190
rlabel metal2 58968 32928 58968 32928 0 net191
rlabel metal2 67312 32760 67312 32760 0 net192
rlabel metal2 98616 34832 98616 34832 0 net193
rlabel metal2 98616 36120 98616 36120 0 net194
rlabel metal2 103208 34160 103208 34160 0 net195
rlabel metal2 105224 34328 105224 34328 0 net196
rlabel metal2 6440 4088 6440 4088 0 net197
rlabel metal2 20832 5320 20832 5320 0 net198
rlabel metal2 69160 6608 69160 6608 0 net199
rlabel metal2 68152 34440 68152 34440 0 net2
rlabel metal2 69048 36568 69048 36568 0 net20
rlabel metal2 68264 5824 68264 5824 0 net200
rlabel metal3 73416 5656 73416 5656 0 net201
rlabel metal2 72968 5656 72968 5656 0 net202
rlabel metal2 74648 5824 74648 5824 0 net203
rlabel metal3 88592 6552 88592 6552 0 net204
rlabel metal2 93688 5880 93688 5880 0 net205
rlabel metal2 101640 5432 101640 5432 0 net206
rlabel metal2 95928 3752 95928 3752 0 net207
rlabel metal2 97160 5656 97160 5656 0 net208
rlabel metal2 19712 5992 19712 5992 0 net209
rlabel metal2 70840 37408 70840 37408 0 net21
rlabel metal2 101752 6888 101752 6888 0 net210
rlabel metal2 143528 4984 143528 4984 0 net211
rlabel metal3 138320 5992 138320 5992 0 net212
rlabel metal2 138936 5208 138936 5208 0 net213
rlabel metal2 118216 4200 118216 4200 0 net214
rlabel metal2 116760 4872 116760 4872 0 net215
rlabel metal3 123200 6440 123200 6440 0 net216
rlabel metal2 116312 6384 116312 6384 0 net217
rlabel metal2 141288 6104 141288 6104 0 net218
rlabel metal2 141736 4984 141736 4984 0 net219
rlabel metal2 72408 32032 72408 32032 0 net22
rlabel metal2 27944 5936 27944 5936 0 net220
rlabel metal2 139944 5208 139944 5208 0 net221
rlabel metal2 146552 5768 146552 5768 0 net222
rlabel metal2 31472 6104 31472 6104 0 net223
rlabel metal2 37464 5936 37464 5936 0 net224
rlabel metal3 38808 4536 38808 4536 0 net225
rlabel metal2 48888 4984 48888 4984 0 net226
rlabel via2 49112 5880 49112 5880 0 net227
rlabel metal3 53144 5880 53144 5880 0 net228
rlabel metal2 67256 7280 67256 7280 0 net229
rlabel metal2 30632 34552 30632 34552 0 net23
rlabel metal2 6776 34440 6776 34440 0 net230
rlabel metal3 75040 35672 75040 35672 0 net231
rlabel metal2 9352 35224 9352 35224 0 net232
rlabel metal2 14280 34832 14280 34832 0 net233
rlabel metal3 17640 34328 17640 34328 0 net234
rlabel metal2 20216 35168 20216 35168 0 net235
rlabel metal3 59472 27832 59472 27832 0 net236
rlabel metal2 26152 30184 26152 30184 0 net237
rlabel metal2 28504 31360 28504 31360 0 net238
rlabel metal2 40880 33096 40880 33096 0 net239
rlabel metal3 75992 35560 75992 35560 0 net24
rlabel metal2 4760 36344 4760 36344 0 net240
rlabel metal2 75544 34328 75544 34328 0 net241
rlabel metal2 75600 36568 75600 36568 0 net25
rlabel metal3 28000 36344 28000 36344 0 net26
rlabel metal2 24248 36624 24248 36624 0 net27
rlabel metal2 26936 36512 26936 36512 0 net28
rlabel metal2 29624 35840 29624 35840 0 net29
rlabel metal3 47880 36400 47880 36400 0 net3
rlabel metal2 47488 33432 47488 33432 0 net30
rlabel metal2 34888 33768 34888 33768 0 net31
rlabel metal2 36344 37240 36344 37240 0 net32
rlabel metal3 22512 34664 22512 34664 0 net33
rlabel metal2 69832 35672 69832 35672 0 net34
rlabel metal3 69048 35112 69048 35112 0 net35
rlabel metal2 77280 36568 77280 36568 0 net36
rlabel metal2 78232 33936 78232 33936 0 net37
rlabel metal3 94640 33432 94640 33432 0 net38
rlabel metal2 90048 34888 90048 34888 0 net39
rlabel metal2 76440 37184 76440 37184 0 net4
rlabel metal3 102480 36680 102480 36680 0 net40
rlabel metal2 102088 34888 102088 34888 0 net41
rlabel metal2 120680 35840 120680 35840 0 net42
rlabel metal2 123144 35224 123144 35224 0 net43
rlabel metal2 22792 36624 22792 36624 0 net44
rlabel metal3 129416 34104 129416 34104 0 net45
rlabel metal2 130760 35448 130760 35448 0 net46
rlabel metal2 139048 34272 139048 34272 0 net47
rlabel metal2 138824 35168 138824 35168 0 net48
rlabel metal2 107688 33488 107688 33488 0 net49
rlabel metal2 43960 37632 43960 37632 0 net5
rlabel metal2 135128 36512 135128 36512 0 net50
rlabel metal3 120232 35448 120232 35448 0 net51
rlabel metal2 139048 36344 139048 36344 0 net52
rlabel metal2 141624 35616 141624 35616 0 net53
rlabel metal2 143808 34104 143808 34104 0 net54
rlabel metal2 30072 36960 30072 36960 0 net55
rlabel metal2 143752 36008 143752 36008 0 net56
rlabel metal2 144872 31780 144872 31780 0 net57
rlabel metal2 31304 34160 31304 34160 0 net58
rlabel metal3 67480 24808 67480 24808 0 net59
rlabel metal2 45640 35560 45640 35560 0 net6
rlabel metal3 49560 34608 49560 34608 0 net60
rlabel metal3 46760 34888 46760 34888 0 net61
rlabel metal2 49784 35168 49784 35168 0 net62
rlabel metal2 69496 32032 69496 32032 0 net63
rlabel metal3 66696 35448 66696 35448 0 net64
rlabel metal2 46424 35112 46424 35112 0 net65
rlabel metal2 63952 3752 63952 3752 0 net66
rlabel metal3 24192 3640 24192 3640 0 net67
rlabel metal2 30408 4200 30408 4200 0 net68
rlabel metal3 45696 36344 45696 36344 0 net69
rlabel metal2 47264 35560 47264 35560 0 net7
rlabel metal2 22288 36344 22288 36344 0 net70
rlabel metal2 43848 3640 43848 3640 0 net71
rlabel metal3 47152 3640 47152 3640 0 net72
rlabel metal2 51520 3640 51520 3640 0 net73
rlabel metal3 51072 23464 51072 23464 0 net74
rlabel metal2 6664 3864 6664 3864 0 net75
rlabel metal2 6664 35560 6664 35560 0 net76
rlabel metal2 52024 32984 52024 32984 0 net77
rlabel metal2 67704 3808 67704 3808 0 net78
rlabel metal2 71792 3752 71792 3752 0 net79
rlabel metal3 51772 36568 51772 36568 0 net8
rlabel metal2 75768 3752 75768 3752 0 net80
rlabel metal3 76104 11704 76104 11704 0 net81
rlabel metal3 81984 8344 81984 8344 0 net82
rlabel metal3 101976 22904 101976 22904 0 net83
rlabel metal2 54488 34048 54488 34048 0 net84
rlabel metal3 95424 8344 95424 8344 0 net85
rlabel metal3 100352 3640 100352 3640 0 net86
rlabel metal2 21896 34328 21896 34328 0 net87
rlabel metal3 103936 3640 103936 3640 0 net88
rlabel metal3 112168 26152 112168 26152 0 net89
rlabel metal2 51128 35784 51128 35784 0 net9
rlabel metal3 109704 3640 109704 3640 0 net90
rlabel metal2 100072 33208 100072 33208 0 net91
rlabel metal3 116536 4872 116536 4872 0 net92
rlabel metal2 121128 5992 121128 5992 0 net93
rlabel metal2 125160 14896 125160 14896 0 net94
rlabel metal2 129136 20160 129136 20160 0 net95
rlabel metal3 139496 36232 139496 36232 0 net96
rlabel metal2 138880 4200 138880 4200 0 net97
rlabel metal3 28728 4200 28728 4200 0 net98
rlabel metal2 143248 4200 143248 4200 0 net99
rlabel metal2 20776 7280 20776 7280 0 operation
rlabel metal2 52584 34160 52584 34160 0 web_mem
rlabel metal2 5712 35000 5712 35000 0 web_mem0
rlabel metal2 78120 35672 78120 35672 0 web_mem1
rlabel metal2 8456 36232 8456 36232 0 wmask_mem0[0]
rlabel metal2 12712 37394 12712 37394 0 wmask_mem0[1]
rlabel metal2 16296 37394 16296 37394 0 wmask_mem0[2]
rlabel metal2 20776 34104 20776 34104 0 wmask_mem0[3]
rlabel metal2 80808 35112 80808 35112 0 wmask_mem1[0]
rlabel metal3 84224 35784 84224 35784 0 wmask_mem1[1]
rlabel metal2 87976 35056 87976 35056 0 wmask_mem1[2]
rlabel metal2 92792 34608 92792 34608 0 wmask_mem1[3]
<< properties >>
string FIXED_BBOX 0 0 150000 40000
<< end >>
