VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_memory
  CLASS BLOCK ;
  FOREIGN wb_memory ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 200.000 ;
  PIN addr_mem0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 31.920 196.000 32.480 200.000 ;
    END
  END addr_mem0[0]
  PIN addr_mem0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.840 196.000 50.400 200.000 ;
    END
  END addr_mem0[1]
  PIN addr_mem0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.760 196.000 68.320 200.000 ;
    END
  END addr_mem0[2]
  PIN addr_mem0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 85.680 196.000 86.240 200.000 ;
    END
  END addr_mem0[3]
  PIN addr_mem0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.600 196.000 104.160 200.000 ;
    END
  END addr_mem0[4]
  PIN addr_mem0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.040 196.000 117.600 200.000 ;
    END
  END addr_mem0[5]
  PIN addr_mem0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.480 196.000 131.040 200.000 ;
    END
  END addr_mem0[6]
  PIN addr_mem0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 143.920 196.000 144.480 200.000 ;
    END
  END addr_mem0[7]
  PIN addr_mem0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.360 196.000 157.920 200.000 ;
    END
  END addr_mem0[8]
  PIN addr_mem1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 385.840 196.000 386.400 200.000 ;
    END
  END addr_mem1[0]
  PIN addr_mem1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.760 196.000 404.320 200.000 ;
    END
  END addr_mem1[1]
  PIN addr_mem1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 421.680 196.000 422.240 200.000 ;
    END
  END addr_mem1[2]
  PIN addr_mem1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.600 196.000 440.160 200.000 ;
    END
  END addr_mem1[3]
  PIN addr_mem1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 457.520 196.000 458.080 200.000 ;
    END
  END addr_mem1[4]
  PIN addr_mem1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.960 196.000 471.520 200.000 ;
    END
  END addr_mem1[5]
  PIN addr_mem1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 484.400 196.000 484.960 200.000 ;
    END
  END addr_mem1[6]
  PIN addr_mem1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.840 196.000 498.400 200.000 ;
    END
  END addr_mem1[7]
  PIN addr_mem1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 511.280 196.000 511.840 200.000 ;
    END
  END addr_mem1[8]
  PIN csb_mem0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.960 196.000 23.520 200.000 ;
    END
  END csb_mem0
  PIN csb_mem1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.880 196.000 377.440 200.000 ;
    END
  END csb_mem1
  PIN din_mem0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.400 196.000 36.960 200.000 ;
    END
  END din_mem0[0]
  PIN din_mem0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.760 196.000 180.320 200.000 ;
    END
  END din_mem0[10]
  PIN din_mem0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.720 196.000 189.280 200.000 ;
    END
  END din_mem0[11]
  PIN din_mem0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.680 196.000 198.240 200.000 ;
    END
  END din_mem0[12]
  PIN din_mem0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 206.640 196.000 207.200 200.000 ;
    END
  END din_mem0[13]
  PIN din_mem0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.600 196.000 216.160 200.000 ;
    END
  END din_mem0[14]
  PIN din_mem0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 224.560 196.000 225.120 200.000 ;
    END
  END din_mem0[15]
  PIN din_mem0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 233.520 196.000 234.080 200.000 ;
    END
  END din_mem0[16]
  PIN din_mem0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 242.480 196.000 243.040 200.000 ;
    END
  END din_mem0[17]
  PIN din_mem0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 251.440 196.000 252.000 200.000 ;
    END
  END din_mem0[18]
  PIN din_mem0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 260.400 196.000 260.960 200.000 ;
    END
  END din_mem0[19]
  PIN din_mem0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 54.320 196.000 54.880 200.000 ;
    END
  END din_mem0[1]
  PIN din_mem0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.360 196.000 269.920 200.000 ;
    END
  END din_mem0[20]
  PIN din_mem0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.320 196.000 278.880 200.000 ;
    END
  END din_mem0[21]
  PIN din_mem0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 287.280 196.000 287.840 200.000 ;
    END
  END din_mem0[22]
  PIN din_mem0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.240 196.000 296.800 200.000 ;
    END
  END din_mem0[23]
  PIN din_mem0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.200 196.000 305.760 200.000 ;
    END
  END din_mem0[24]
  PIN din_mem0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 314.160 196.000 314.720 200.000 ;
    END
  END din_mem0[25]
  PIN din_mem0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.120 196.000 323.680 200.000 ;
    END
  END din_mem0[26]
  PIN din_mem0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.080 196.000 332.640 200.000 ;
    END
  END din_mem0[27]
  PIN din_mem0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 341.040 196.000 341.600 200.000 ;
    END
  END din_mem0[28]
  PIN din_mem0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 350.000 196.000 350.560 200.000 ;
    END
  END din_mem0[29]
  PIN din_mem0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.240 196.000 72.800 200.000 ;
    END
  END din_mem0[2]
  PIN din_mem0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 358.960 196.000 359.520 200.000 ;
    END
  END din_mem0[30]
  PIN din_mem0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 367.920 196.000 368.480 200.000 ;
    END
  END din_mem0[31]
  PIN din_mem0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.160 196.000 90.720 200.000 ;
    END
  END din_mem0[3]
  PIN din_mem0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.080 196.000 108.640 200.000 ;
    END
  END din_mem0[4]
  PIN din_mem0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 121.520 196.000 122.080 200.000 ;
    END
  END din_mem0[5]
  PIN din_mem0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.960 196.000 135.520 200.000 ;
    END
  END din_mem0[6]
  PIN din_mem0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.400 196.000 148.960 200.000 ;
    END
  END din_mem0[7]
  PIN din_mem0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.840 196.000 162.400 200.000 ;
    END
  END din_mem0[8]
  PIN din_mem0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.800 196.000 171.360 200.000 ;
    END
  END din_mem0[9]
  PIN din_mem1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.320 196.000 390.880 200.000 ;
    END
  END din_mem1[0]
  PIN din_mem1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 533.680 196.000 534.240 200.000 ;
    END
  END din_mem1[10]
  PIN din_mem1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 542.640 196.000 543.200 200.000 ;
    END
  END din_mem1[11]
  PIN din_mem1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.600 196.000 552.160 200.000 ;
    END
  END din_mem1[12]
  PIN din_mem1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 560.560 196.000 561.120 200.000 ;
    END
  END din_mem1[13]
  PIN din_mem1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 569.520 196.000 570.080 200.000 ;
    END
  END din_mem1[14]
  PIN din_mem1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 578.480 196.000 579.040 200.000 ;
    END
  END din_mem1[15]
  PIN din_mem1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 587.440 196.000 588.000 200.000 ;
    END
  END din_mem1[16]
  PIN din_mem1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 596.400 196.000 596.960 200.000 ;
    END
  END din_mem1[17]
  PIN din_mem1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 605.360 196.000 605.920 200.000 ;
    END
  END din_mem1[18]
  PIN din_mem1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 614.320 196.000 614.880 200.000 ;
    END
  END din_mem1[19]
  PIN din_mem1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 408.240 196.000 408.800 200.000 ;
    END
  END din_mem1[1]
  PIN din_mem1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 623.280 196.000 623.840 200.000 ;
    END
  END din_mem1[20]
  PIN din_mem1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 632.240 196.000 632.800 200.000 ;
    END
  END din_mem1[21]
  PIN din_mem1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 641.200 196.000 641.760 200.000 ;
    END
  END din_mem1[22]
  PIN din_mem1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 650.160 196.000 650.720 200.000 ;
    END
  END din_mem1[23]
  PIN din_mem1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 659.120 196.000 659.680 200.000 ;
    END
  END din_mem1[24]
  PIN din_mem1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 668.080 196.000 668.640 200.000 ;
    END
  END din_mem1[25]
  PIN din_mem1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 677.040 196.000 677.600 200.000 ;
    END
  END din_mem1[26]
  PIN din_mem1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 686.000 196.000 686.560 200.000 ;
    END
  END din_mem1[27]
  PIN din_mem1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 694.960 196.000 695.520 200.000 ;
    END
  END din_mem1[28]
  PIN din_mem1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 703.920 196.000 704.480 200.000 ;
    END
  END din_mem1[29]
  PIN din_mem1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.160 196.000 426.720 200.000 ;
    END
  END din_mem1[2]
  PIN din_mem1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 712.880 196.000 713.440 200.000 ;
    END
  END din_mem1[30]
  PIN din_mem1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 721.840 196.000 722.400 200.000 ;
    END
  END din_mem1[31]
  PIN din_mem1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 444.080 196.000 444.640 200.000 ;
    END
  END din_mem1[3]
  PIN din_mem1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 462.000 196.000 462.560 200.000 ;
    END
  END din_mem1[4]
  PIN din_mem1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 475.440 196.000 476.000 200.000 ;
    END
  END din_mem1[5]
  PIN din_mem1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 488.880 196.000 489.440 200.000 ;
    END
  END din_mem1[6]
  PIN din_mem1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 502.320 196.000 502.880 200.000 ;
    END
  END din_mem1[7]
  PIN din_mem1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 515.760 196.000 516.320 200.000 ;
    END
  END din_mem1[8]
  PIN din_mem1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.720 196.000 525.280 200.000 ;
    END
  END din_mem1[9]
  PIN dout_mem0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.880 196.000 41.440 200.000 ;
    END
  END dout_mem0[0]
  PIN dout_mem0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.240 196.000 184.800 200.000 ;
    END
  END dout_mem0[10]
  PIN dout_mem0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 193.200 196.000 193.760 200.000 ;
    END
  END dout_mem0[11]
  PIN dout_mem0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 202.160 196.000 202.720 200.000 ;
    END
  END dout_mem0[12]
  PIN dout_mem0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.120 196.000 211.680 200.000 ;
    END
  END dout_mem0[13]
  PIN dout_mem0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 220.080 196.000 220.640 200.000 ;
    END
  END dout_mem0[14]
  PIN dout_mem0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.040 196.000 229.600 200.000 ;
    END
  END dout_mem0[15]
  PIN dout_mem0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.000 196.000 238.560 200.000 ;
    END
  END dout_mem0[16]
  PIN dout_mem0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 246.960 196.000 247.520 200.000 ;
    END
  END dout_mem0[17]
  PIN dout_mem0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.920 196.000 256.480 200.000 ;
    END
  END dout_mem0[18]
  PIN dout_mem0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 264.880 196.000 265.440 200.000 ;
    END
  END dout_mem0[19]
  PIN dout_mem0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.800 196.000 59.360 200.000 ;
    END
  END dout_mem0[1]
  PIN dout_mem0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.840 196.000 274.400 200.000 ;
    END
  END dout_mem0[20]
  PIN dout_mem0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.800 196.000 283.360 200.000 ;
    END
  END dout_mem0[21]
  PIN dout_mem0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.760 196.000 292.320 200.000 ;
    END
  END dout_mem0[22]
  PIN dout_mem0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 300.720 196.000 301.280 200.000 ;
    END
  END dout_mem0[23]
  PIN dout_mem0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.680 196.000 310.240 200.000 ;
    END
  END dout_mem0[24]
  PIN dout_mem0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.640 196.000 319.200 200.000 ;
    END
  END dout_mem0[25]
  PIN dout_mem0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 327.600 196.000 328.160 200.000 ;
    END
  END dout_mem0[26]
  PIN dout_mem0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.560 196.000 337.120 200.000 ;
    END
  END dout_mem0[27]
  PIN dout_mem0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 345.520 196.000 346.080 200.000 ;
    END
  END dout_mem0[28]
  PIN dout_mem0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 354.480 196.000 355.040 200.000 ;
    END
  END dout_mem0[29]
  PIN dout_mem0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 76.720 196.000 77.280 200.000 ;
    END
  END dout_mem0[2]
  PIN dout_mem0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 363.440 196.000 364.000 200.000 ;
    END
  END dout_mem0[30]
  PIN dout_mem0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.400 196.000 372.960 200.000 ;
    END
  END dout_mem0[31]
  PIN dout_mem0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.640 196.000 95.200 200.000 ;
    END
  END dout_mem0[3]
  PIN dout_mem0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.560 196.000 113.120 200.000 ;
    END
  END dout_mem0[4]
  PIN dout_mem0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.000 196.000 126.560 200.000 ;
    END
  END dout_mem0[5]
  PIN dout_mem0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 139.440 196.000 140.000 200.000 ;
    END
  END dout_mem0[6]
  PIN dout_mem0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.880 196.000 153.440 200.000 ;
    END
  END dout_mem0[7]
  PIN dout_mem0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.320 196.000 166.880 200.000 ;
    END
  END dout_mem0[8]
  PIN dout_mem0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.280 196.000 175.840 200.000 ;
    END
  END dout_mem0[9]
  PIN dout_mem1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 394.800 196.000 395.360 200.000 ;
    END
  END dout_mem1[0]
  PIN dout_mem1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 538.160 196.000 538.720 200.000 ;
    END
  END dout_mem1[10]
  PIN dout_mem1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.120 196.000 547.680 200.000 ;
    END
  END dout_mem1[11]
  PIN dout_mem1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 556.080 196.000 556.640 200.000 ;
    END
  END dout_mem1[12]
  PIN dout_mem1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 565.040 196.000 565.600 200.000 ;
    END
  END dout_mem1[13]
  PIN dout_mem1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 574.000 196.000 574.560 200.000 ;
    END
  END dout_mem1[14]
  PIN dout_mem1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 582.960 196.000 583.520 200.000 ;
    END
  END dout_mem1[15]
  PIN dout_mem1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.920 196.000 592.480 200.000 ;
    END
  END dout_mem1[16]
  PIN dout_mem1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 600.880 196.000 601.440 200.000 ;
    END
  END dout_mem1[17]
  PIN dout_mem1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 609.840 196.000 610.400 200.000 ;
    END
  END dout_mem1[18]
  PIN dout_mem1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.800 196.000 619.360 200.000 ;
    END
  END dout_mem1[19]
  PIN dout_mem1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 412.720 196.000 413.280 200.000 ;
    END
  END dout_mem1[1]
  PIN dout_mem1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 627.760 196.000 628.320 200.000 ;
    END
  END dout_mem1[20]
  PIN dout_mem1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 636.720 196.000 637.280 200.000 ;
    END
  END dout_mem1[21]
  PIN dout_mem1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.680 196.000 646.240 200.000 ;
    END
  END dout_mem1[22]
  PIN dout_mem1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 654.640 196.000 655.200 200.000 ;
    END
  END dout_mem1[23]
  PIN dout_mem1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 663.600 196.000 664.160 200.000 ;
    END
  END dout_mem1[24]
  PIN dout_mem1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.560 196.000 673.120 200.000 ;
    END
  END dout_mem1[25]
  PIN dout_mem1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 681.520 196.000 682.080 200.000 ;
    END
  END dout_mem1[26]
  PIN dout_mem1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 690.480 196.000 691.040 200.000 ;
    END
  END dout_mem1[27]
  PIN dout_mem1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 699.440 196.000 700.000 200.000 ;
    END
  END dout_mem1[28]
  PIN dout_mem1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 708.400 196.000 708.960 200.000 ;
    END
  END dout_mem1[29]
  PIN dout_mem1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.640 196.000 431.200 200.000 ;
    END
  END dout_mem1[2]
  PIN dout_mem1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 717.360 196.000 717.920 200.000 ;
    END
  END dout_mem1[30]
  PIN dout_mem1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 726.320 196.000 726.880 200.000 ;
    END
  END dout_mem1[31]
  PIN dout_mem1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 448.560 196.000 449.120 200.000 ;
    END
  END dout_mem1[3]
  PIN dout_mem1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 466.480 196.000 467.040 200.000 ;
    END
  END dout_mem1[4]
  PIN dout_mem1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 479.920 196.000 480.480 200.000 ;
    END
  END dout_mem1[5]
  PIN dout_mem1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 493.360 196.000 493.920 200.000 ;
    END
  END dout_mem1[6]
  PIN dout_mem1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 506.800 196.000 507.360 200.000 ;
    END
  END dout_mem1[7]
  PIN dout_mem1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.240 196.000 520.800 200.000 ;
    END
  END dout_mem1[8]
  PIN dout_mem1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 529.200 196.000 529.760 200.000 ;
    END
  END dout_mem1[9]
  PIN io_wbs_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.840 0.000 22.400 4.000 ;
    END
  END io_wbs_ack
  PIN io_wbs_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 62.160 0.000 62.720 4.000 ;
    END
  END io_wbs_adr[0]
  PIN io_wbs_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 290.640 0.000 291.200 4.000 ;
    END
  END io_wbs_adr[10]
  PIN io_wbs_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 310.800 0.000 311.360 4.000 ;
    END
  END io_wbs_adr[11]
  PIN io_wbs_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 330.960 0.000 331.520 4.000 ;
    END
  END io_wbs_adr[12]
  PIN io_wbs_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.120 0.000 351.680 4.000 ;
    END
  END io_wbs_adr[13]
  PIN io_wbs_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.280 0.000 371.840 4.000 ;
    END
  END io_wbs_adr[14]
  PIN io_wbs_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 391.440 0.000 392.000 4.000 ;
    END
  END io_wbs_adr[15]
  PIN io_wbs_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 411.600 0.000 412.160 4.000 ;
    END
  END io_wbs_adr[16]
  PIN io_wbs_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 431.760 0.000 432.320 4.000 ;
    END
  END io_wbs_adr[17]
  PIN io_wbs_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 451.920 0.000 452.480 4.000 ;
    END
  END io_wbs_adr[18]
  PIN io_wbs_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 472.080 0.000 472.640 4.000 ;
    END
  END io_wbs_adr[19]
  PIN io_wbs_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.040 0.000 89.600 4.000 ;
    END
  END io_wbs_adr[1]
  PIN io_wbs_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 492.240 0.000 492.800 4.000 ;
    END
  END io_wbs_adr[20]
  PIN io_wbs_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 512.400 0.000 512.960 4.000 ;
    END
  END io_wbs_adr[21]
  PIN io_wbs_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.560 0.000 533.120 4.000 ;
    END
  END io_wbs_adr[22]
  PIN io_wbs_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 552.720 0.000 553.280 4.000 ;
    END
  END io_wbs_adr[23]
  PIN io_wbs_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 572.880 0.000 573.440 4.000 ;
    END
  END io_wbs_adr[24]
  PIN io_wbs_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 593.040 0.000 593.600 4.000 ;
    END
  END io_wbs_adr[25]
  PIN io_wbs_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 613.200 0.000 613.760 4.000 ;
    END
  END io_wbs_adr[26]
  PIN io_wbs_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 633.360 0.000 633.920 4.000 ;
    END
  END io_wbs_adr[27]
  PIN io_wbs_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 653.520 0.000 654.080 4.000 ;
    END
  END io_wbs_adr[28]
  PIN io_wbs_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 673.680 0.000 674.240 4.000 ;
    END
  END io_wbs_adr[29]
  PIN io_wbs_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 115.920 0.000 116.480 4.000 ;
    END
  END io_wbs_adr[2]
  PIN io_wbs_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 693.840 0.000 694.400 4.000 ;
    END
  END io_wbs_adr[30]
  PIN io_wbs_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 714.000 0.000 714.560 4.000 ;
    END
  END io_wbs_adr[31]
  PIN io_wbs_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.800 0.000 143.360 4.000 ;
    END
  END io_wbs_adr[3]
  PIN io_wbs_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.680 0.000 170.240 4.000 ;
    END
  END io_wbs_adr[4]
  PIN io_wbs_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 189.840 0.000 190.400 4.000 ;
    END
  END io_wbs_adr[5]
  PIN io_wbs_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 210.000 0.000 210.560 4.000 ;
    END
  END io_wbs_adr[6]
  PIN io_wbs_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 230.160 0.000 230.720 4.000 ;
    END
  END io_wbs_adr[7]
  PIN io_wbs_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 250.320 0.000 250.880 4.000 ;
    END
  END io_wbs_adr[8]
  PIN io_wbs_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 270.480 0.000 271.040 4.000 ;
    END
  END io_wbs_adr[9]
  PIN io_wbs_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 28.560 0.000 29.120 4.000 ;
    END
  END io_wbs_clk
  PIN io_wbs_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 35.280 0.000 35.840 4.000 ;
    END
  END io_wbs_cyc
  PIN io_wbs_datrd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.880 0.000 69.440 4.000 ;
    END
  END io_wbs_datrd[0]
  PIN io_wbs_datrd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 297.360 0.000 297.920 4.000 ;
    END
  END io_wbs_datrd[10]
  PIN io_wbs_datrd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 317.520 0.000 318.080 4.000 ;
    END
  END io_wbs_datrd[11]
  PIN io_wbs_datrd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 337.680 0.000 338.240 4.000 ;
    END
  END io_wbs_datrd[12]
  PIN io_wbs_datrd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 357.840 0.000 358.400 4.000 ;
    END
  END io_wbs_datrd[13]
  PIN io_wbs_datrd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.000 0.000 378.560 4.000 ;
    END
  END io_wbs_datrd[14]
  PIN io_wbs_datrd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 398.160 0.000 398.720 4.000 ;
    END
  END io_wbs_datrd[15]
  PIN io_wbs_datrd[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.320 0.000 418.880 4.000 ;
    END
  END io_wbs_datrd[16]
  PIN io_wbs_datrd[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 438.480 0.000 439.040 4.000 ;
    END
  END io_wbs_datrd[17]
  PIN io_wbs_datrd[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 458.640 0.000 459.200 4.000 ;
    END
  END io_wbs_datrd[18]
  PIN io_wbs_datrd[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 478.800 0.000 479.360 4.000 ;
    END
  END io_wbs_datrd[19]
  PIN io_wbs_datrd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.760 0.000 96.320 4.000 ;
    END
  END io_wbs_datrd[1]
  PIN io_wbs_datrd[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 498.960 0.000 499.520 4.000 ;
    END
  END io_wbs_datrd[20]
  PIN io_wbs_datrd[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 519.120 0.000 519.680 4.000 ;
    END
  END io_wbs_datrd[21]
  PIN io_wbs_datrd[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 539.280 0.000 539.840 4.000 ;
    END
  END io_wbs_datrd[22]
  PIN io_wbs_datrd[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 559.440 0.000 560.000 4.000 ;
    END
  END io_wbs_datrd[23]
  PIN io_wbs_datrd[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 579.600 0.000 580.160 4.000 ;
    END
  END io_wbs_datrd[24]
  PIN io_wbs_datrd[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.760 0.000 600.320 4.000 ;
    END
  END io_wbs_datrd[25]
  PIN io_wbs_datrd[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 619.920 0.000 620.480 4.000 ;
    END
  END io_wbs_datrd[26]
  PIN io_wbs_datrd[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 640.080 0.000 640.640 4.000 ;
    END
  END io_wbs_datrd[27]
  PIN io_wbs_datrd[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 660.240 0.000 660.800 4.000 ;
    END
  END io_wbs_datrd[28]
  PIN io_wbs_datrd[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 680.400 0.000 680.960 4.000 ;
    END
  END io_wbs_datrd[29]
  PIN io_wbs_datrd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 122.640 0.000 123.200 4.000 ;
    END
  END io_wbs_datrd[2]
  PIN io_wbs_datrd[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 700.560 0.000 701.120 4.000 ;
    END
  END io_wbs_datrd[30]
  PIN io_wbs_datrd[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.720 0.000 721.280 4.000 ;
    END
  END io_wbs_datrd[31]
  PIN io_wbs_datrd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 149.520 0.000 150.080 4.000 ;
    END
  END io_wbs_datrd[3]
  PIN io_wbs_datrd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.400 0.000 176.960 4.000 ;
    END
  END io_wbs_datrd[4]
  PIN io_wbs_datrd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 196.560 0.000 197.120 4.000 ;
    END
  END io_wbs_datrd[5]
  PIN io_wbs_datrd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 216.720 0.000 217.280 4.000 ;
    END
  END io_wbs_datrd[6]
  PIN io_wbs_datrd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 236.880 0.000 237.440 4.000 ;
    END
  END io_wbs_datrd[7]
  PIN io_wbs_datrd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 257.040 0.000 257.600 4.000 ;
    END
  END io_wbs_datrd[8]
  PIN io_wbs_datrd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 277.200 0.000 277.760 4.000 ;
    END
  END io_wbs_datrd[9]
  PIN io_wbs_datwr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.600 0.000 76.160 4.000 ;
    END
  END io_wbs_datwr[0]
  PIN io_wbs_datwr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.080 0.000 304.640 4.000 ;
    END
  END io_wbs_datwr[10]
  PIN io_wbs_datwr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 324.240 0.000 324.800 4.000 ;
    END
  END io_wbs_datwr[11]
  PIN io_wbs_datwr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 344.400 0.000 344.960 4.000 ;
    END
  END io_wbs_datwr[12]
  PIN io_wbs_datwr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.560 0.000 365.120 4.000 ;
    END
  END io_wbs_datwr[13]
  PIN io_wbs_datwr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 384.720 0.000 385.280 4.000 ;
    END
  END io_wbs_datwr[14]
  PIN io_wbs_datwr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 404.880 0.000 405.440 4.000 ;
    END
  END io_wbs_datwr[15]
  PIN io_wbs_datwr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 425.040 0.000 425.600 4.000 ;
    END
  END io_wbs_datwr[16]
  PIN io_wbs_datwr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.200 0.000 445.760 4.000 ;
    END
  END io_wbs_datwr[17]
  PIN io_wbs_datwr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 465.360 0.000 465.920 4.000 ;
    END
  END io_wbs_datwr[18]
  PIN io_wbs_datwr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 485.520 0.000 486.080 4.000 ;
    END
  END io_wbs_datwr[19]
  PIN io_wbs_datwr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 102.480 0.000 103.040 4.000 ;
    END
  END io_wbs_datwr[1]
  PIN io_wbs_datwr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 505.680 0.000 506.240 4.000 ;
    END
  END io_wbs_datwr[20]
  PIN io_wbs_datwr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 525.840 0.000 526.400 4.000 ;
    END
  END io_wbs_datwr[21]
  PIN io_wbs_datwr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 546.000 0.000 546.560 4.000 ;
    END
  END io_wbs_datwr[22]
  PIN io_wbs_datwr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 566.160 0.000 566.720 4.000 ;
    END
  END io_wbs_datwr[23]
  PIN io_wbs_datwr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 586.320 0.000 586.880 4.000 ;
    END
  END io_wbs_datwr[24]
  PIN io_wbs_datwr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 606.480 0.000 607.040 4.000 ;
    END
  END io_wbs_datwr[25]
  PIN io_wbs_datwr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 626.640 0.000 627.200 4.000 ;
    END
  END io_wbs_datwr[26]
  PIN io_wbs_datwr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 646.800 0.000 647.360 4.000 ;
    END
  END io_wbs_datwr[27]
  PIN io_wbs_datwr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 666.960 0.000 667.520 4.000 ;
    END
  END io_wbs_datwr[28]
  PIN io_wbs_datwr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 687.120 0.000 687.680 4.000 ;
    END
  END io_wbs_datwr[29]
  PIN io_wbs_datwr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 129.360 0.000 129.920 4.000 ;
    END
  END io_wbs_datwr[2]
  PIN io_wbs_datwr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 707.280 0.000 707.840 4.000 ;
    END
  END io_wbs_datwr[30]
  PIN io_wbs_datwr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 727.440 0.000 728.000 4.000 ;
    END
  END io_wbs_datwr[31]
  PIN io_wbs_datwr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 156.240 0.000 156.800 4.000 ;
    END
  END io_wbs_datwr[3]
  PIN io_wbs_datwr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.120 0.000 183.680 4.000 ;
    END
  END io_wbs_datwr[4]
  PIN io_wbs_datwr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 203.280 0.000 203.840 4.000 ;
    END
  END io_wbs_datwr[5]
  PIN io_wbs_datwr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 223.440 0.000 224.000 4.000 ;
    END
  END io_wbs_datwr[6]
  PIN io_wbs_datwr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 243.600 0.000 244.160 4.000 ;
    END
  END io_wbs_datwr[7]
  PIN io_wbs_datwr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 263.760 0.000 264.320 4.000 ;
    END
  END io_wbs_datwr[8]
  PIN io_wbs_datwr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 283.920 0.000 284.480 4.000 ;
    END
  END io_wbs_datwr[9]
  PIN io_wbs_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 42.000 0.000 42.560 4.000 ;
    END
  END io_wbs_rst
  PIN io_wbs_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 82.320 0.000 82.880 4.000 ;
    END
  END io_wbs_sel[0]
  PIN io_wbs_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 109.200 0.000 109.760 4.000 ;
    END
  END io_wbs_sel[1]
  PIN io_wbs_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.080 0.000 136.640 4.000 ;
    END
  END io_wbs_sel[2]
  PIN io_wbs_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.960 0.000 163.520 4.000 ;
    END
  END io_wbs_sel[3]
  PIN io_wbs_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 48.720 0.000 49.280 4.000 ;
    END
  END io_wbs_stb
  PIN io_wbs_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 55.440 0.000 56.000 4.000 ;
    END
  END io_wbs_we
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 97.970 15.380 99.570 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 282.070 15.380 283.670 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 466.170 15.380 467.770 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 650.270 15.380 651.870 184.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 190.020 15.380 191.620 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.120 15.380 375.720 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 558.220 15.380 559.820 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 742.320 15.380 743.920 184.540 ;
    END
  END vss
  PIN web_mem0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 27.440 196.000 28.000 200.000 ;
    END
  END web_mem0
  PIN web_mem1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 381.360 196.000 381.920 200.000 ;
    END
  END web_mem1
  PIN wmask_mem0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.360 196.000 45.920 200.000 ;
    END
  END wmask_mem0[0]
  PIN wmask_mem0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.280 196.000 63.840 200.000 ;
    END
  END wmask_mem0[1]
  PIN wmask_mem0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.200 196.000 81.760 200.000 ;
    END
  END wmask_mem0[2]
  PIN wmask_mem0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 99.120 196.000 99.680 200.000 ;
    END
  END wmask_mem0[3]
  PIN wmask_mem1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.280 196.000 399.840 200.000 ;
    END
  END wmask_mem1[0]
  PIN wmask_mem1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 417.200 196.000 417.760 200.000 ;
    END
  END wmask_mem1[1]
  PIN wmask_mem1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 435.120 196.000 435.680 200.000 ;
    END
  END wmask_mem1[2]
  PIN wmask_mem1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.040 196.000 453.600 200.000 ;
    END
  END wmask_mem1[3]
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 743.920 186.890 ;
      LAYER Metal2 ;
        RECT 21.980 195.700 22.660 196.420 ;
        RECT 23.820 195.700 27.140 196.420 ;
        RECT 28.300 195.700 31.620 196.420 ;
        RECT 32.780 195.700 36.100 196.420 ;
        RECT 37.260 195.700 40.580 196.420 ;
        RECT 41.740 195.700 45.060 196.420 ;
        RECT 46.220 195.700 49.540 196.420 ;
        RECT 50.700 195.700 54.020 196.420 ;
        RECT 55.180 195.700 58.500 196.420 ;
        RECT 59.660 195.700 62.980 196.420 ;
        RECT 64.140 195.700 67.460 196.420 ;
        RECT 68.620 195.700 71.940 196.420 ;
        RECT 73.100 195.700 76.420 196.420 ;
        RECT 77.580 195.700 80.900 196.420 ;
        RECT 82.060 195.700 85.380 196.420 ;
        RECT 86.540 195.700 89.860 196.420 ;
        RECT 91.020 195.700 94.340 196.420 ;
        RECT 95.500 195.700 98.820 196.420 ;
        RECT 99.980 195.700 103.300 196.420 ;
        RECT 104.460 195.700 107.780 196.420 ;
        RECT 108.940 195.700 112.260 196.420 ;
        RECT 113.420 195.700 116.740 196.420 ;
        RECT 117.900 195.700 121.220 196.420 ;
        RECT 122.380 195.700 125.700 196.420 ;
        RECT 126.860 195.700 130.180 196.420 ;
        RECT 131.340 195.700 134.660 196.420 ;
        RECT 135.820 195.700 139.140 196.420 ;
        RECT 140.300 195.700 143.620 196.420 ;
        RECT 144.780 195.700 148.100 196.420 ;
        RECT 149.260 195.700 152.580 196.420 ;
        RECT 153.740 195.700 157.060 196.420 ;
        RECT 158.220 195.700 161.540 196.420 ;
        RECT 162.700 195.700 166.020 196.420 ;
        RECT 167.180 195.700 170.500 196.420 ;
        RECT 171.660 195.700 174.980 196.420 ;
        RECT 176.140 195.700 179.460 196.420 ;
        RECT 180.620 195.700 183.940 196.420 ;
        RECT 185.100 195.700 188.420 196.420 ;
        RECT 189.580 195.700 192.900 196.420 ;
        RECT 194.060 195.700 197.380 196.420 ;
        RECT 198.540 195.700 201.860 196.420 ;
        RECT 203.020 195.700 206.340 196.420 ;
        RECT 207.500 195.700 210.820 196.420 ;
        RECT 211.980 195.700 215.300 196.420 ;
        RECT 216.460 195.700 219.780 196.420 ;
        RECT 220.940 195.700 224.260 196.420 ;
        RECT 225.420 195.700 228.740 196.420 ;
        RECT 229.900 195.700 233.220 196.420 ;
        RECT 234.380 195.700 237.700 196.420 ;
        RECT 238.860 195.700 242.180 196.420 ;
        RECT 243.340 195.700 246.660 196.420 ;
        RECT 247.820 195.700 251.140 196.420 ;
        RECT 252.300 195.700 255.620 196.420 ;
        RECT 256.780 195.700 260.100 196.420 ;
        RECT 261.260 195.700 264.580 196.420 ;
        RECT 265.740 195.700 269.060 196.420 ;
        RECT 270.220 195.700 273.540 196.420 ;
        RECT 274.700 195.700 278.020 196.420 ;
        RECT 279.180 195.700 282.500 196.420 ;
        RECT 283.660 195.700 286.980 196.420 ;
        RECT 288.140 195.700 291.460 196.420 ;
        RECT 292.620 195.700 295.940 196.420 ;
        RECT 297.100 195.700 300.420 196.420 ;
        RECT 301.580 195.700 304.900 196.420 ;
        RECT 306.060 195.700 309.380 196.420 ;
        RECT 310.540 195.700 313.860 196.420 ;
        RECT 315.020 195.700 318.340 196.420 ;
        RECT 319.500 195.700 322.820 196.420 ;
        RECT 323.980 195.700 327.300 196.420 ;
        RECT 328.460 195.700 331.780 196.420 ;
        RECT 332.940 195.700 336.260 196.420 ;
        RECT 337.420 195.700 340.740 196.420 ;
        RECT 341.900 195.700 345.220 196.420 ;
        RECT 346.380 195.700 349.700 196.420 ;
        RECT 350.860 195.700 354.180 196.420 ;
        RECT 355.340 195.700 358.660 196.420 ;
        RECT 359.820 195.700 363.140 196.420 ;
        RECT 364.300 195.700 367.620 196.420 ;
        RECT 368.780 195.700 372.100 196.420 ;
        RECT 373.260 195.700 376.580 196.420 ;
        RECT 377.740 195.700 381.060 196.420 ;
        RECT 382.220 195.700 385.540 196.420 ;
        RECT 386.700 195.700 390.020 196.420 ;
        RECT 391.180 195.700 394.500 196.420 ;
        RECT 395.660 195.700 398.980 196.420 ;
        RECT 400.140 195.700 403.460 196.420 ;
        RECT 404.620 195.700 407.940 196.420 ;
        RECT 409.100 195.700 412.420 196.420 ;
        RECT 413.580 195.700 416.900 196.420 ;
        RECT 418.060 195.700 421.380 196.420 ;
        RECT 422.540 195.700 425.860 196.420 ;
        RECT 427.020 195.700 430.340 196.420 ;
        RECT 431.500 195.700 434.820 196.420 ;
        RECT 435.980 195.700 439.300 196.420 ;
        RECT 440.460 195.700 443.780 196.420 ;
        RECT 444.940 195.700 448.260 196.420 ;
        RECT 449.420 195.700 452.740 196.420 ;
        RECT 453.900 195.700 457.220 196.420 ;
        RECT 458.380 195.700 461.700 196.420 ;
        RECT 462.860 195.700 466.180 196.420 ;
        RECT 467.340 195.700 470.660 196.420 ;
        RECT 471.820 195.700 475.140 196.420 ;
        RECT 476.300 195.700 479.620 196.420 ;
        RECT 480.780 195.700 484.100 196.420 ;
        RECT 485.260 195.700 488.580 196.420 ;
        RECT 489.740 195.700 493.060 196.420 ;
        RECT 494.220 195.700 497.540 196.420 ;
        RECT 498.700 195.700 502.020 196.420 ;
        RECT 503.180 195.700 506.500 196.420 ;
        RECT 507.660 195.700 510.980 196.420 ;
        RECT 512.140 195.700 515.460 196.420 ;
        RECT 516.620 195.700 519.940 196.420 ;
        RECT 521.100 195.700 524.420 196.420 ;
        RECT 525.580 195.700 528.900 196.420 ;
        RECT 530.060 195.700 533.380 196.420 ;
        RECT 534.540 195.700 537.860 196.420 ;
        RECT 539.020 195.700 542.340 196.420 ;
        RECT 543.500 195.700 546.820 196.420 ;
        RECT 547.980 195.700 551.300 196.420 ;
        RECT 552.460 195.700 555.780 196.420 ;
        RECT 556.940 195.700 560.260 196.420 ;
        RECT 561.420 195.700 564.740 196.420 ;
        RECT 565.900 195.700 569.220 196.420 ;
        RECT 570.380 195.700 573.700 196.420 ;
        RECT 574.860 195.700 578.180 196.420 ;
        RECT 579.340 195.700 582.660 196.420 ;
        RECT 583.820 195.700 587.140 196.420 ;
        RECT 588.300 195.700 591.620 196.420 ;
        RECT 592.780 195.700 596.100 196.420 ;
        RECT 597.260 195.700 600.580 196.420 ;
        RECT 601.740 195.700 605.060 196.420 ;
        RECT 606.220 195.700 609.540 196.420 ;
        RECT 610.700 195.700 614.020 196.420 ;
        RECT 615.180 195.700 618.500 196.420 ;
        RECT 619.660 195.700 622.980 196.420 ;
        RECT 624.140 195.700 627.460 196.420 ;
        RECT 628.620 195.700 631.940 196.420 ;
        RECT 633.100 195.700 636.420 196.420 ;
        RECT 637.580 195.700 640.900 196.420 ;
        RECT 642.060 195.700 645.380 196.420 ;
        RECT 646.540 195.700 649.860 196.420 ;
        RECT 651.020 195.700 654.340 196.420 ;
        RECT 655.500 195.700 658.820 196.420 ;
        RECT 659.980 195.700 663.300 196.420 ;
        RECT 664.460 195.700 667.780 196.420 ;
        RECT 668.940 195.700 672.260 196.420 ;
        RECT 673.420 195.700 676.740 196.420 ;
        RECT 677.900 195.700 681.220 196.420 ;
        RECT 682.380 195.700 685.700 196.420 ;
        RECT 686.860 195.700 690.180 196.420 ;
        RECT 691.340 195.700 694.660 196.420 ;
        RECT 695.820 195.700 699.140 196.420 ;
        RECT 700.300 195.700 703.620 196.420 ;
        RECT 704.780 195.700 708.100 196.420 ;
        RECT 709.260 195.700 712.580 196.420 ;
        RECT 713.740 195.700 717.060 196.420 ;
        RECT 718.220 195.700 721.540 196.420 ;
        RECT 722.700 195.700 726.020 196.420 ;
        RECT 727.180 195.700 743.780 196.420 ;
        RECT 21.980 4.300 743.780 195.700 ;
        RECT 22.700 3.500 28.260 4.300 ;
        RECT 29.420 3.500 34.980 4.300 ;
        RECT 36.140 3.500 41.700 4.300 ;
        RECT 42.860 3.500 48.420 4.300 ;
        RECT 49.580 3.500 55.140 4.300 ;
        RECT 56.300 3.500 61.860 4.300 ;
        RECT 63.020 3.500 68.580 4.300 ;
        RECT 69.740 3.500 75.300 4.300 ;
        RECT 76.460 3.500 82.020 4.300 ;
        RECT 83.180 3.500 88.740 4.300 ;
        RECT 89.900 3.500 95.460 4.300 ;
        RECT 96.620 3.500 102.180 4.300 ;
        RECT 103.340 3.500 108.900 4.300 ;
        RECT 110.060 3.500 115.620 4.300 ;
        RECT 116.780 3.500 122.340 4.300 ;
        RECT 123.500 3.500 129.060 4.300 ;
        RECT 130.220 3.500 135.780 4.300 ;
        RECT 136.940 3.500 142.500 4.300 ;
        RECT 143.660 3.500 149.220 4.300 ;
        RECT 150.380 3.500 155.940 4.300 ;
        RECT 157.100 3.500 162.660 4.300 ;
        RECT 163.820 3.500 169.380 4.300 ;
        RECT 170.540 3.500 176.100 4.300 ;
        RECT 177.260 3.500 182.820 4.300 ;
        RECT 183.980 3.500 189.540 4.300 ;
        RECT 190.700 3.500 196.260 4.300 ;
        RECT 197.420 3.500 202.980 4.300 ;
        RECT 204.140 3.500 209.700 4.300 ;
        RECT 210.860 3.500 216.420 4.300 ;
        RECT 217.580 3.500 223.140 4.300 ;
        RECT 224.300 3.500 229.860 4.300 ;
        RECT 231.020 3.500 236.580 4.300 ;
        RECT 237.740 3.500 243.300 4.300 ;
        RECT 244.460 3.500 250.020 4.300 ;
        RECT 251.180 3.500 256.740 4.300 ;
        RECT 257.900 3.500 263.460 4.300 ;
        RECT 264.620 3.500 270.180 4.300 ;
        RECT 271.340 3.500 276.900 4.300 ;
        RECT 278.060 3.500 283.620 4.300 ;
        RECT 284.780 3.500 290.340 4.300 ;
        RECT 291.500 3.500 297.060 4.300 ;
        RECT 298.220 3.500 303.780 4.300 ;
        RECT 304.940 3.500 310.500 4.300 ;
        RECT 311.660 3.500 317.220 4.300 ;
        RECT 318.380 3.500 323.940 4.300 ;
        RECT 325.100 3.500 330.660 4.300 ;
        RECT 331.820 3.500 337.380 4.300 ;
        RECT 338.540 3.500 344.100 4.300 ;
        RECT 345.260 3.500 350.820 4.300 ;
        RECT 351.980 3.500 357.540 4.300 ;
        RECT 358.700 3.500 364.260 4.300 ;
        RECT 365.420 3.500 370.980 4.300 ;
        RECT 372.140 3.500 377.700 4.300 ;
        RECT 378.860 3.500 384.420 4.300 ;
        RECT 385.580 3.500 391.140 4.300 ;
        RECT 392.300 3.500 397.860 4.300 ;
        RECT 399.020 3.500 404.580 4.300 ;
        RECT 405.740 3.500 411.300 4.300 ;
        RECT 412.460 3.500 418.020 4.300 ;
        RECT 419.180 3.500 424.740 4.300 ;
        RECT 425.900 3.500 431.460 4.300 ;
        RECT 432.620 3.500 438.180 4.300 ;
        RECT 439.340 3.500 444.900 4.300 ;
        RECT 446.060 3.500 451.620 4.300 ;
        RECT 452.780 3.500 458.340 4.300 ;
        RECT 459.500 3.500 465.060 4.300 ;
        RECT 466.220 3.500 471.780 4.300 ;
        RECT 472.940 3.500 478.500 4.300 ;
        RECT 479.660 3.500 485.220 4.300 ;
        RECT 486.380 3.500 491.940 4.300 ;
        RECT 493.100 3.500 498.660 4.300 ;
        RECT 499.820 3.500 505.380 4.300 ;
        RECT 506.540 3.500 512.100 4.300 ;
        RECT 513.260 3.500 518.820 4.300 ;
        RECT 519.980 3.500 525.540 4.300 ;
        RECT 526.700 3.500 532.260 4.300 ;
        RECT 533.420 3.500 538.980 4.300 ;
        RECT 540.140 3.500 545.700 4.300 ;
        RECT 546.860 3.500 552.420 4.300 ;
        RECT 553.580 3.500 559.140 4.300 ;
        RECT 560.300 3.500 565.860 4.300 ;
        RECT 567.020 3.500 572.580 4.300 ;
        RECT 573.740 3.500 579.300 4.300 ;
        RECT 580.460 3.500 586.020 4.300 ;
        RECT 587.180 3.500 592.740 4.300 ;
        RECT 593.900 3.500 599.460 4.300 ;
        RECT 600.620 3.500 606.180 4.300 ;
        RECT 607.340 3.500 612.900 4.300 ;
        RECT 614.060 3.500 619.620 4.300 ;
        RECT 620.780 3.500 626.340 4.300 ;
        RECT 627.500 3.500 633.060 4.300 ;
        RECT 634.220 3.500 639.780 4.300 ;
        RECT 640.940 3.500 646.500 4.300 ;
        RECT 647.660 3.500 653.220 4.300 ;
        RECT 654.380 3.500 659.940 4.300 ;
        RECT 661.100 3.500 666.660 4.300 ;
        RECT 667.820 3.500 673.380 4.300 ;
        RECT 674.540 3.500 680.100 4.300 ;
        RECT 681.260 3.500 686.820 4.300 ;
        RECT 687.980 3.500 693.540 4.300 ;
        RECT 694.700 3.500 700.260 4.300 ;
        RECT 701.420 3.500 706.980 4.300 ;
        RECT 708.140 3.500 713.700 4.300 ;
        RECT 714.860 3.500 720.420 4.300 ;
        RECT 721.580 3.500 727.140 4.300 ;
        RECT 728.300 3.500 743.780 4.300 ;
      LAYER Metal3 ;
        RECT 28.650 12.460 743.830 194.740 ;
      LAYER Metal4 ;
        RECT 217.980 125.530 281.770 181.910 ;
        RECT 283.970 125.530 373.820 181.910 ;
        RECT 376.020 125.530 465.870 181.910 ;
        RECT 468.070 125.530 557.920 181.910 ;
        RECT 560.120 125.530 575.540 181.910 ;
  END
END wb_memory
END LIBRARY

